magic
tech sky130A
magscale 1 2
timestamp 1724369829
<< pwell >>
rect 5780 1530 5860 1570
rect 5980 1540 6080 1590
rect 1360 -1610 1420 -1550
rect 1220 -1990 1310 -1900
rect 1230 -2560 1300 -2400
rect 1600 -2690 1690 -2620
rect 1600 -2920 1690 -2850
rect 1230 -3010 1300 -2940
rect 1230 -3240 1300 -3170
rect 1970 -3450 2050 -3370
rect 1230 -3730 1300 -3580
rect 1230 -4170 1300 -4100
rect 1230 -4400 1300 -4330
rect 1230 -4830 1300 -4760
rect 3270 -9200 3490 -7712
<< locali >>
rect 880 4410 930 4420
<< viali >>
rect 540 4700 720 4750
rect 980 4690 1230 4740
rect 450 4360 500 4650
rect 880 4600 930 4650
rect 880 4370 930 4410
rect 1280 4370 1320 4640
rect 540 4270 720 4320
rect 1120 4280 1230 4320
rect 1720 3170 2030 3220
rect 1470 2880 1520 3130
rect 1570 2690 1770 2830
rect 5290 2500 5470 2550
rect 5900 2510 6160 2550
rect 5290 2090 5470 2140
rect 5300 1830 5460 1880
rect 1570 1680 1730 1810
rect 5800 1510 5840 1560
rect 6210 1510 6260 2460
rect 5300 1420 5460 1470
rect 5900 1420 6160 1460
rect 5340 970 5500 1020
rect 6160 980 6280 1030
rect 1570 660 1740 800
rect 5340 560 5500 610
rect 5340 170 5500 220
rect 2220 100 2460 150
rect 1570 -50 1740 -10
rect 1570 -280 1740 -240
rect 2500 -340 2560 60
rect 5340 -240 5500 -190
rect 2220 -430 2460 -380
rect 5910 -810 5960 -140
rect 6320 -810 6380 920
rect 6010 -910 6270 -860
rect 1570 -1010 1740 -950
rect 1480 -1180 1650 -1130
rect 5340 -1390 5500 -1340
rect 6030 -1380 6270 -1340
rect 2050 -1470 2660 -1420
rect 1480 -1700 1650 -1650
rect 1480 -1960 1650 -1910
rect 2690 -2080 2750 -1500
rect 5340 -1800 5500 -1750
rect 2050 -2160 2660 -2110
rect 5340 -2190 5500 -2140
rect 1480 -2470 1650 -2420
rect 1750 -2580 1910 -2540
rect 5340 -2600 5500 -2550
rect 2480 -2910 2660 -2860
rect 1750 -3000 1910 -2960
rect 1750 -3220 1910 -3180
rect 2700 -3230 2760 -2950
rect 2480 -3320 2660 -3270
rect 1750 -3640 1910 -3600
rect 1550 -3730 1710 -3690
rect 2140 -4070 2700 -4010
rect 1550 -4150 1710 -4110
rect 1550 -4390 1710 -4350
rect 2740 -4390 2800 -4110
rect 2140 -4490 2700 -4430
rect 1550 -4810 1710 -4770
rect 5900 -4780 5960 -2500
rect 6320 -4780 6380 -1430
rect 890 -5990 6200 -5920
rect 6820 -7260 6870 -6040
rect 890 -7370 6200 -7300
rect 890 -7790 6200 -7720
rect 3420 -9070 3610 -7840
rect 6820 -9060 6870 -7840
rect 1000 -9250 6710 -9120
rect 6820 -10520 6870 -9300
rect 890 -10640 6200 -10570
<< metal1 >>
rect 1350 4920 1442 5196
rect 1718 4920 1810 5196
rect 2086 4920 2178 5196
rect 2454 4920 2546 5196
rect 2822 4920 2914 5196
rect 3190 4920 3282 5196
rect 3558 4920 3650 5196
rect 3926 4920 4018 5196
rect 4294 4920 4386 5196
rect 4662 4920 4754 5196
rect 5030 4920 5122 5196
rect 5398 4920 5490 5196
rect 5766 4920 5858 5196
rect 6134 4920 6226 5196
rect 6502 4920 6594 5196
rect 6870 4920 6962 5196
rect 1360 4860 1620 4920
rect 420 4750 740 4780
rect 420 4700 540 4750
rect 720 4700 740 4750
rect 420 4690 740 4700
rect 870 4740 1470 4750
rect 870 4690 980 4740
rect 1230 4690 1470 4740
rect 420 4650 530 4690
rect 870 4680 1470 4690
rect 870 4660 950 4680
rect 420 4360 450 4650
rect 500 4570 530 4650
rect 590 4600 880 4660
rect 940 4600 950 4660
rect 1190 4640 1470 4680
rect 710 4590 950 4600
rect 980 4590 1160 4640
rect 500 4450 610 4570
rect 980 4560 1070 4590
rect 1190 4560 1280 4640
rect 650 4460 1070 4560
rect 1160 4460 1280 4560
rect 500 4360 530 4450
rect 710 4420 940 4430
rect 590 4360 850 4420
rect 420 4330 530 4360
rect 840 4350 850 4360
rect 930 4350 940 4420
rect 840 4340 940 4350
rect 970 4420 1070 4460
rect 1170 4450 1280 4460
rect 970 4370 1160 4420
rect 1190 4370 1280 4450
rect 1320 4370 1470 4640
rect 420 4320 740 4330
rect 420 4270 540 4320
rect 720 4270 740 4320
rect 420 4180 740 4270
rect 970 4210 1070 4370
rect 1190 4340 1470 4370
rect 420 4020 440 4180
rect 720 4020 740 4180
rect 420 4000 740 4020
rect 890 3970 1070 4210
rect 1100 4320 1470 4340
rect 1100 4280 1120 4320
rect 1230 4280 1470 4320
rect 1100 4150 1470 4280
rect 1560 4320 1620 4860
rect 1730 4440 1790 4920
rect 2105 4545 2155 4920
rect 2475 4645 2525 4920
rect 2845 4735 2895 4920
rect 3215 4865 3265 4920
rect 3215 4815 3355 4865
rect 2845 4685 3185 4735
rect 2475 4595 2995 4645
rect 2105 4495 2695 4545
rect 1730 4380 2540 4440
rect 1560 4260 2390 4320
rect 1100 4100 1530 4150
rect 890 3950 1100 3970
rect 890 3850 910 3950
rect 1080 3850 1100 3950
rect 890 3830 1100 3850
rect 1160 3800 1530 4100
rect 1160 3600 1180 3800
rect 1470 3600 1530 3800
rect 1160 3490 1530 3600
rect 1220 3130 1530 3490
rect 1710 3780 2040 3800
rect 1710 3620 1730 3780
rect 2020 3620 2040 3780
rect 1560 3460 1660 3470
rect 1560 3350 1570 3460
rect 1650 3350 1660 3460
rect 1560 3340 1660 3350
rect 1220 2880 1470 3130
rect 1520 2880 1530 3130
rect 1570 2950 1620 3340
rect 1710 3220 2040 3620
rect 2090 3460 2190 3470
rect 2090 3350 2100 3460
rect 2180 3350 2190 3460
rect 2090 3340 2190 3350
rect 1710 3170 1720 3220
rect 2030 3170 2040 3220
rect 1710 3120 2040 3170
rect 1650 3060 2070 3120
rect 2100 2950 2150 3340
rect 2330 3250 2390 4260
rect 2480 3250 2540 4380
rect 2645 3250 2695 4495
rect 2945 3250 2995 4595
rect 2324 3190 2330 3250
rect 2390 3190 2396 3250
rect 2474 3190 2480 3250
rect 2540 3190 2546 3250
rect 2630 3246 2710 3250
rect 2630 3194 2644 3246
rect 2696 3194 2710 3246
rect 2630 3190 2710 3194
rect 2930 3246 3010 3250
rect 3135 3246 3185 4685
rect 3305 3246 3355 4815
rect 3585 4645 3635 4920
rect 3465 4595 3635 4645
rect 3465 3246 3515 4595
rect 3945 4545 3995 4920
rect 3625 4495 3995 4545
rect 3625 3246 3675 4495
rect 4325 4435 4375 4920
rect 3765 4385 4375 4435
rect 3765 3246 3815 4385
rect 4685 4315 4735 4920
rect 3915 4265 4735 4315
rect 5045 4265 5095 4920
rect 3915 3246 3965 4265
rect 5045 4215 5260 4265
rect 2930 3194 2944 3246
rect 2996 3194 3010 3246
rect 3128 3194 3134 3246
rect 3186 3194 3192 3246
rect 3298 3194 3304 3246
rect 3356 3194 3362 3246
rect 3458 3194 3464 3246
rect 3516 3194 3522 3246
rect 3618 3194 3624 3246
rect 3676 3194 3682 3246
rect 3758 3194 3764 3246
rect 3816 3194 3822 3246
rect 3908 3194 3914 3246
rect 3966 3194 3972 3246
rect 2930 3190 3010 3194
rect 1650 2890 2070 2950
rect 1220 2850 1530 2880
rect 1220 2830 1790 2850
rect 1220 2810 1570 2830
rect 1220 2700 1240 2810
rect 1350 2700 1570 2810
rect 1220 2690 1570 2700
rect 1770 2690 1790 2830
rect 1220 2680 1790 2690
rect 1610 2580 1710 2640
rect 1770 2580 1780 2640
rect 1850 2540 2060 2890
rect 5210 2845 5260 4215
rect 5415 2966 5465 4920
rect 5780 3520 5840 4920
rect 6150 3660 6210 4920
rect 6520 4200 6580 4920
rect 6890 4390 6950 4920
rect 6890 4330 6986 4390
rect 6520 4140 6868 4200
rect 6150 3600 6480 3660
rect 5780 3460 6340 3520
rect 6280 3250 6340 3460
rect 6420 3250 6480 3600
rect 6274 3190 6280 3250
rect 6340 3190 6346 3250
rect 6414 3190 6420 3250
rect 6480 3190 6486 3250
rect 6808 3248 6868 4140
rect 6926 3248 6986 4330
rect 6802 3188 6808 3248
rect 6868 3188 6874 3248
rect 6920 3188 6926 3248
rect 6986 3188 6992 3248
rect 5408 2914 5414 2966
rect 5466 2914 5472 2966
rect 5210 2795 5680 2845
rect 610 2520 1630 2540
rect 610 1980 630 2520
rect 790 1980 1630 2520
rect 610 1960 1630 1980
rect 1670 1960 2060 2540
rect 4900 2560 5490 2570
rect 4900 2490 4910 2560
rect 5030 2550 5490 2560
rect 5030 2500 5290 2550
rect 5470 2500 5490 2550
rect 5030 2490 5490 2500
rect 4900 2480 5490 2490
rect 5630 2450 5680 2795
rect 5880 2550 6750 2570
rect 5270 2400 5680 2450
rect 5730 2510 5830 2520
rect 5730 2430 5740 2510
rect 5820 2470 5830 2510
rect 5880 2510 5900 2550
rect 6160 2510 6570 2550
rect 5880 2500 6570 2510
rect 5820 2430 6080 2470
rect 5730 2420 6080 2430
rect 4050 2360 5360 2370
rect 4050 2280 4060 2360
rect 4240 2280 5360 2360
rect 4050 2270 5360 2280
rect 5400 2360 5590 2370
rect 5400 2280 5510 2360
rect 5580 2280 5590 2360
rect 5400 2270 5590 2280
rect 5630 2240 5680 2400
rect 5980 2390 6080 2420
rect 6200 2460 6570 2500
rect 5340 2190 5680 2240
rect 4900 2150 5490 2160
rect 4900 2080 4910 2150
rect 5030 2140 5490 2150
rect 5030 2090 5290 2140
rect 5470 2090 5490 2140
rect 5030 2080 5490 2090
rect 4900 2070 5490 2080
rect 1610 1860 1710 1920
rect 1770 1860 1780 1920
rect 1220 1810 1790 1820
rect 1220 1800 1570 1810
rect 1220 1690 1240 1800
rect 1350 1690 1570 1800
rect 1220 1680 1570 1690
rect 1730 1680 1790 1810
rect 1220 1670 1790 1680
rect 1610 1570 1710 1630
rect 1770 1570 1780 1630
rect 1850 1530 2060 1960
rect 4620 2020 6165 2030
rect 4620 1950 4630 2020
rect 4810 1950 6165 2020
rect 4620 1940 6165 1950
rect 4900 1890 5490 1900
rect 4900 1820 4910 1890
rect 5030 1880 5490 1890
rect 5030 1830 5300 1880
rect 5460 1830 5490 1880
rect 5030 1820 5490 1830
rect 4900 1810 5490 1820
rect 5629 1876 5681 1882
rect 5629 1818 5681 1824
rect 5630 1780 5680 1818
rect 5280 1730 5680 1780
rect 4330 1630 5360 1700
rect 4330 1550 4350 1630
rect 4510 1600 5360 1630
rect 5400 1690 5590 1700
rect 5400 1610 5510 1690
rect 5580 1610 5590 1690
rect 5400 1600 5590 1610
rect 4510 1550 4600 1600
rect 5630 1570 5680 1730
rect 4330 1530 4600 1550
rect 290 1510 1630 1530
rect 290 970 310 1510
rect 470 970 1630 1510
rect 290 950 1630 970
rect 1670 950 2060 1530
rect 5340 1520 5680 1570
rect 5780 1560 5860 1570
rect 5780 1510 5800 1560
rect 5840 1550 5860 1560
rect 5980 1550 6080 1590
rect 6200 1550 6210 2460
rect 5840 1510 6210 1550
rect 6260 1510 6570 2460
rect 4900 1480 5490 1490
rect 4900 1410 4910 1480
rect 5030 1470 5490 1480
rect 5030 1420 5300 1470
rect 5460 1420 5490 1470
rect 5030 1410 5490 1420
rect 4900 1400 5490 1410
rect 5780 1460 6570 1510
rect 5780 1420 5900 1460
rect 6160 1420 6570 1460
rect 6730 1420 6750 2550
rect 5780 1400 6750 1420
rect 4900 1030 5520 1040
rect 4900 970 4910 1030
rect 5030 1020 5520 1030
rect 5030 970 5340 1020
rect 5500 970 5520 1020
rect 6140 1030 6750 1050
rect 4900 960 5520 970
rect 5990 980 6110 990
rect 5620 930 5700 940
rect 5620 920 5630 930
rect 1220 870 1370 890
rect 1220 760 1240 870
rect 1350 810 1370 870
rect 1610 850 1710 910
rect 1770 850 1780 910
rect 5390 870 5630 920
rect 5690 870 5700 930
rect 5990 900 6000 980
rect 6080 940 6110 980
rect 6140 980 6160 1030
rect 6280 980 6570 1030
rect 6140 970 6570 980
rect 6080 900 6190 940
rect 5990 890 6190 900
rect 5620 860 5700 870
rect 6090 860 6190 890
rect 6310 920 6570 970
rect 4050 830 4250 850
rect 1350 800 1790 810
rect 1350 760 1570 800
rect 1220 730 1570 760
rect 1220 660 1230 730
rect 1300 670 1570 730
rect 1300 660 1310 670
rect 1220 650 1310 660
rect 1550 660 1570 670
rect 1740 740 1790 800
rect 4050 750 4070 830
rect 4220 750 5400 830
rect 5440 820 5980 830
rect 5440 760 5890 820
rect 5970 760 5980 820
rect 5440 750 5980 760
rect 1740 710 2830 740
rect 4050 730 4250 750
rect 5620 710 5700 720
rect 1740 660 2650 710
rect 1550 650 2650 660
rect 2630 640 2650 650
rect 2810 640 2830 710
rect 5390 660 5630 710
rect 5620 650 5630 660
rect 5690 650 5700 710
rect 5620 640 5700 650
rect 1350 630 1430 640
rect 1350 570 1360 630
rect 1420 610 1430 630
rect 2630 620 2830 640
rect 2273 610 2279 611
rect 1420 570 2279 610
rect 1350 560 2279 570
rect 2273 559 2279 560
rect 2331 559 2337 611
rect 4900 610 5520 620
rect 4900 550 4910 610
rect 5030 560 5340 610
rect 5500 560 5520 610
rect 5030 550 5520 560
rect 4900 540 5520 550
rect 610 510 1620 530
rect 610 160 630 510
rect 790 160 1620 510
rect 610 140 1620 160
rect 1670 510 1870 520
rect 1670 150 1780 510
rect 1860 150 1870 510
rect 4620 440 6280 450
rect 4620 350 4630 440
rect 4810 350 6280 440
rect 4620 340 6280 350
rect 4900 230 5520 240
rect 1670 140 1870 150
rect 2200 160 2830 180
rect 4900 170 4910 230
rect 5030 220 5520 230
rect 5030 170 5340 220
rect 5500 170 5520 220
rect 4900 160 5520 170
rect 2200 150 2650 160
rect 2200 100 2220 150
rect 2460 100 2650 150
rect 1350 90 1680 100
rect 2200 90 2650 100
rect 1350 30 1360 90
rect 1420 50 1680 90
rect 2480 60 2650 90
rect 1420 30 1430 50
rect 1350 20 1430 30
rect 1220 10 1300 20
rect 1220 -50 1230 10
rect 1290 -20 1300 10
rect 1910 0 2380 50
rect 1550 -10 1760 0
rect 1550 -20 1570 -10
rect 1290 -50 1570 -20
rect 1740 -50 1760 -10
rect 1220 -60 1760 -50
rect 890 -100 1090 -80
rect 1910 -100 1960 0
rect 2480 -30 2500 60
rect 890 -190 910 -100
rect 1070 -190 1960 -100
rect 890 -210 1090 -190
rect 1220 -240 1760 -230
rect 1220 -300 1230 -240
rect 1290 -270 1570 -240
rect 1290 -300 1300 -270
rect 1550 -280 1570 -270
rect 1740 -280 1760 -240
rect 1550 -290 1760 -280
rect 1910 -280 1960 -190
rect 2000 -50 2280 -40
rect 2000 -230 2010 -50
rect 2140 -230 2280 -50
rect 2000 -240 2280 -230
rect 2390 -250 2500 -30
rect 1220 -310 1300 -300
rect 1350 -320 1430 -310
rect 1350 -380 1360 -320
rect 1420 -340 1430 -320
rect 1910 -330 2380 -280
rect 2480 -340 2500 -250
rect 2560 -340 2650 60
rect 1420 -380 1680 -340
rect 2480 -370 2650 -340
rect 1350 -390 1680 -380
rect 2200 -380 2650 -370
rect 290 -440 1620 -420
rect 2200 -430 2220 -380
rect 2460 -430 2650 -380
rect 290 -790 310 -440
rect 470 -790 1620 -440
rect 290 -810 1620 -790
rect 1670 -440 1870 -430
rect 1670 -800 1780 -440
rect 1860 -800 1870 -440
rect 2200 -440 2650 -430
rect 2810 -440 2830 160
rect 5620 130 5700 140
rect 5620 120 5630 130
rect 5390 70 5630 120
rect 5690 70 5700 130
rect 5620 60 5700 70
rect 4330 30 4530 50
rect 4330 -50 4350 30
rect 4510 -50 5400 30
rect 5440 20 5980 30
rect 5440 -40 5890 20
rect 5970 -40 5980 20
rect 5440 -50 5980 -40
rect 4330 -70 4530 -50
rect 5620 -90 5700 -80
rect 5390 -140 5630 -90
rect 5620 -150 5630 -140
rect 5690 -150 5700 -90
rect 5620 -160 5700 -150
rect 5890 -140 5980 -110
rect 4900 -190 5520 -180
rect 4900 -250 4910 -190
rect 5030 -240 5340 -190
rect 5500 -240 5520 -190
rect 5030 -250 5520 -240
rect 4900 -260 5520 -250
rect 2200 -460 2830 -440
rect 1670 -810 1870 -800
rect 5890 -810 5910 -140
rect 5960 -780 5980 -140
rect 6090 -780 6190 -750
rect 6310 -780 6320 920
rect 5960 -810 6320 -780
rect 6380 -810 6570 920
rect 2273 -850 2279 -849
rect 1350 -860 2279 -850
rect 1350 -920 1360 -860
rect 1420 -900 2279 -860
rect 1420 -920 1430 -900
rect 2273 -901 2279 -900
rect 2331 -901 2337 -849
rect 5890 -860 6570 -810
rect 5890 -910 6010 -860
rect 6270 -910 6570 -860
rect 6730 -910 6750 1030
rect 1350 -930 1430 -920
rect 2630 -930 2830 -910
rect 5890 -930 6750 -910
rect 2630 -940 2650 -930
rect 1220 -950 1310 -940
rect 1220 -1020 1230 -950
rect 1300 -960 1310 -950
rect 1550 -950 2650 -940
rect 1550 -960 1570 -950
rect 1300 -1010 1570 -960
rect 1740 -1010 2650 -950
rect 1300 -1020 2650 -1010
rect 1220 -1030 2650 -1020
rect 1460 -1130 2650 -1030
rect 1460 -1180 1480 -1130
rect 1650 -1170 2650 -1130
rect 2810 -1170 2830 -930
rect 1650 -1180 2830 -1170
rect 1460 -1190 2830 -1180
rect 1350 -1210 1430 -1200
rect 1350 -1270 1360 -1210
rect 1420 -1230 1430 -1210
rect 2273 -1230 2279 -1229
rect 1420 -1270 2279 -1230
rect 1350 -1280 2279 -1270
rect 2273 -1281 2279 -1280
rect 2331 -1281 2337 -1229
rect 610 -1330 1540 -1310
rect 610 -1490 630 -1330
rect 790 -1490 1540 -1330
rect 610 -1510 1540 -1490
rect 1580 -1320 1770 -1310
rect 1580 -1500 1690 -1320
rect 1760 -1500 1770 -1320
rect 4900 -1330 5520 -1320
rect 4900 -1390 4910 -1330
rect 5030 -1340 5520 -1330
rect 5030 -1390 5340 -1340
rect 5500 -1390 5520 -1340
rect 6010 -1340 6750 -1320
rect 4900 -1400 5520 -1390
rect 5880 -1380 5980 -1370
rect 2030 -1420 3030 -1410
rect 2030 -1470 2050 -1420
rect 2660 -1430 3030 -1420
rect 2660 -1470 2850 -1430
rect 2030 -1480 2850 -1470
rect 1580 -1510 1770 -1500
rect 2680 -1500 2850 -1480
rect 1350 -1550 1600 -1540
rect 1350 -1610 1360 -1550
rect 1420 -1590 1600 -1550
rect 1800 -1570 2570 -1520
rect 1420 -1610 1430 -1590
rect 1350 -1620 1430 -1610
rect 1220 -1630 1310 -1620
rect 1220 -1700 1230 -1630
rect 1300 -1650 1310 -1630
rect 1460 -1650 1670 -1640
rect 1300 -1700 1480 -1650
rect 1650 -1700 1670 -1650
rect 1220 -1710 1670 -1700
rect 890 -1720 1090 -1710
rect 890 -1870 910 -1720
rect 1070 -1740 1090 -1720
rect 1800 -1740 1850 -1570
rect 2680 -1600 2690 -1500
rect 1070 -1860 1850 -1740
rect 1070 -1870 1090 -1860
rect 890 -1890 1090 -1870
rect 1220 -1910 1670 -1890
rect 1220 -1980 1230 -1910
rect 1300 -1950 1480 -1910
rect 1300 -1980 1310 -1950
rect 1460 -1960 1480 -1950
rect 1650 -1960 1670 -1910
rect 1460 -1970 1670 -1960
rect 1220 -1990 1310 -1980
rect 1350 -1990 1430 -1980
rect 1350 -2050 1360 -1990
rect 1420 -2010 1430 -1990
rect 1800 -2010 1850 -1860
rect 1890 -1620 2110 -1610
rect 1890 -1960 1900 -1620
rect 1990 -1960 2110 -1620
rect 1890 -1970 2110 -1960
rect 2580 -1980 2690 -1600
rect 1420 -2050 1600 -2010
rect 1350 -2060 1600 -2050
rect 1800 -2060 2570 -2010
rect 2680 -2080 2690 -1980
rect 2750 -2080 2850 -1500
rect 290 -2110 1540 -2090
rect 290 -2270 310 -2110
rect 470 -2270 1540 -2110
rect 290 -2290 1540 -2270
rect 1580 -2100 1770 -2090
rect 2680 -2100 2850 -2080
rect 1580 -2280 1690 -2100
rect 1760 -2280 1770 -2100
rect 2030 -2110 2850 -2100
rect 2030 -2160 2050 -2110
rect 2660 -2150 2850 -2110
rect 3010 -2150 3030 -1430
rect 5620 -1430 5700 -1420
rect 5620 -1440 5630 -1430
rect 5390 -1490 5630 -1440
rect 5690 -1490 5700 -1430
rect 5880 -1440 5890 -1380
rect 5970 -1420 5980 -1380
rect 6010 -1380 6030 -1340
rect 6270 -1380 6570 -1340
rect 6010 -1390 6570 -1380
rect 5970 -1440 6190 -1420
rect 5880 -1480 6190 -1440
rect 6310 -1430 6570 -1390
rect 5620 -1500 5700 -1490
rect 4050 -1530 4250 -1510
rect 4050 -1610 4070 -1530
rect 4220 -1610 5400 -1530
rect 5440 -1540 5980 -1530
rect 5440 -1600 5890 -1540
rect 5970 -1600 5980 -1540
rect 5440 -1610 5980 -1600
rect 4050 -1630 4250 -1610
rect 5620 -1650 5700 -1640
rect 5390 -1700 5630 -1650
rect 5620 -1710 5630 -1700
rect 5690 -1710 5700 -1650
rect 5620 -1720 5700 -1710
rect 4900 -1750 5520 -1740
rect 4900 -1810 4910 -1750
rect 5030 -1800 5340 -1750
rect 5500 -1800 5520 -1750
rect 5030 -1810 5520 -1800
rect 4900 -1820 5520 -1810
rect 4620 -1920 6280 -1910
rect 4620 -2020 4630 -1920
rect 4810 -2020 6280 -1920
rect 4620 -2030 6280 -2020
rect 2660 -2160 3030 -2150
rect 2030 -2170 3030 -2160
rect 4900 -2130 5520 -2120
rect 4900 -2190 4910 -2130
rect 5030 -2140 5520 -2130
rect 5030 -2190 5340 -2140
rect 5500 -2190 5520 -2140
rect 4900 -2200 5520 -2190
rect 5620 -2230 5700 -2220
rect 5620 -2240 5630 -2230
rect 1580 -2290 1770 -2280
rect 5390 -2290 5630 -2240
rect 5690 -2290 5700 -2230
rect 5620 -2300 5700 -2290
rect 2273 -2320 2279 -2319
rect 1350 -2330 2279 -2320
rect 1350 -2390 1360 -2330
rect 1420 -2370 2279 -2330
rect 1420 -2390 1430 -2370
rect 2273 -2371 2279 -2370
rect 2331 -2371 2337 -2319
rect 4330 -2330 4530 -2310
rect 1220 -2400 1310 -2390
rect 1350 -2400 1430 -2390
rect 1220 -2560 1230 -2400
rect 1300 -2430 1310 -2400
rect 4330 -2410 4350 -2330
rect 4510 -2410 5400 -2330
rect 5440 -2340 5980 -2330
rect 5440 -2400 5890 -2340
rect 5970 -2400 5980 -2340
rect 5440 -2410 5980 -2400
rect 1460 -2420 3030 -2410
rect 1460 -2430 1480 -2420
rect 1300 -2470 1480 -2430
rect 1650 -2430 3030 -2420
rect 4330 -2430 4530 -2410
rect 1650 -2470 2850 -2430
rect 1300 -2540 2850 -2470
rect 1300 -2560 1750 -2540
rect 1220 -2570 1750 -2560
rect 1730 -2580 1750 -2570
rect 1910 -2550 2850 -2540
rect 3010 -2550 3030 -2430
rect 5620 -2450 5700 -2440
rect 5390 -2500 5630 -2450
rect 5620 -2510 5630 -2500
rect 5690 -2510 5700 -2450
rect 5620 -2520 5700 -2510
rect 5890 -2500 5970 -2480
rect 1910 -2570 3030 -2550
rect 4900 -2550 5520 -2540
rect 1910 -2580 1930 -2570
rect 1730 -2600 1930 -2580
rect 4900 -2610 4910 -2550
rect 5030 -2600 5340 -2550
rect 5500 -2600 5520 -2550
rect 5030 -2610 5520 -2600
rect 4900 -2620 5520 -2610
rect 1600 -2680 1610 -2620
rect 1680 -2640 1690 -2620
rect 2303 -2640 2309 -2639
rect 1680 -2680 2309 -2640
rect 610 -2700 810 -2680
rect 1600 -2690 2309 -2680
rect 2303 -2691 2309 -2690
rect 2361 -2691 2367 -2639
rect 610 -2840 630 -2700
rect 790 -2720 810 -2700
rect 790 -2820 1810 -2720
rect 1860 -2730 2060 -2720
rect 1860 -2810 1970 -2730
rect 2050 -2810 2060 -2730
rect 1860 -2820 2060 -2810
rect 790 -2840 810 -2820
rect 610 -2860 810 -2840
rect 1600 -2860 1880 -2850
rect 1600 -2920 1610 -2860
rect 1680 -2900 1880 -2860
rect 2460 -2860 3030 -2850
rect 1680 -2920 1690 -2900
rect 2460 -2910 2480 -2860
rect 2660 -2870 3030 -2860
rect 2660 -2910 2850 -2870
rect 2460 -2920 2850 -2910
rect 1220 -2940 1310 -2930
rect 1220 -3010 1230 -2940
rect 1300 -2950 1310 -2940
rect 1730 -2950 1940 -2940
rect 1300 -2960 1940 -2950
rect 1300 -3000 1750 -2960
rect 1910 -3000 1940 -2960
rect 1300 -3010 1940 -3000
rect 1220 -3020 1940 -3010
rect 2060 -2960 2430 -2930
rect 2620 -2950 2850 -2920
rect 2060 -2970 2580 -2960
rect 890 -3040 1090 -3020
rect 890 -3140 910 -3040
rect 1070 -3050 1090 -3040
rect 2060 -3050 2100 -2970
rect 1070 -3130 2100 -3050
rect 1070 -3140 1090 -3130
rect 890 -3160 1090 -3140
rect 1220 -3170 1940 -3160
rect 1220 -3240 1230 -3170
rect 1300 -3180 1940 -3170
rect 1300 -3220 1750 -3180
rect 1910 -3220 1940 -3180
rect 1300 -3230 1940 -3220
rect 1300 -3240 1310 -3230
rect 1730 -3240 1940 -3230
rect 2060 -3210 2100 -3130
rect 2130 -3010 2360 -3000
rect 2390 -3010 2580 -2970
rect 2130 -3170 2140 -3010
rect 2270 -3030 2360 -3010
rect 2620 -3030 2700 -2950
rect 2270 -3050 2370 -3030
rect 2600 -3050 2700 -3030
rect 2270 -3130 2380 -3050
rect 2590 -3130 2700 -3050
rect 2270 -3150 2370 -3130
rect 2600 -3150 2700 -3130
rect 2270 -3170 2360 -3150
rect 2130 -3180 2360 -3170
rect 2390 -3210 2580 -3170
rect 2060 -3220 2580 -3210
rect 1220 -3250 1310 -3240
rect 2060 -3250 2430 -3220
rect 2620 -3230 2700 -3150
rect 2760 -3230 2850 -2950
rect 2620 -3260 2850 -3230
rect 1600 -3320 1610 -3260
rect 1680 -3280 1690 -3260
rect 2460 -3270 2850 -3260
rect 1680 -3320 1880 -3280
rect 1600 -3330 1880 -3320
rect 2460 -3320 2480 -3270
rect 2660 -3310 2850 -3270
rect 3010 -3310 3030 -2870
rect 2660 -3320 3030 -3310
rect 2460 -3330 3030 -3320
rect 290 -3360 490 -3340
rect 290 -3460 310 -3360
rect 470 -3460 1810 -3360
rect 1860 -3370 2060 -3360
rect 1860 -3450 1970 -3370
rect 2050 -3450 2060 -3370
rect 1860 -3460 2060 -3450
rect 290 -3480 490 -3460
rect 2298 -3490 2304 -3489
rect 1600 -3500 2304 -3490
rect 1600 -3560 1610 -3500
rect 1680 -3540 2304 -3500
rect 1680 -3560 1690 -3540
rect 2298 -3541 2304 -3540
rect 2356 -3541 2362 -3489
rect 1220 -3580 1310 -3570
rect 1220 -3730 1230 -3580
rect 1300 -3590 1310 -3580
rect 1730 -3590 1940 -3580
rect 1300 -3600 3030 -3590
rect 1300 -3640 1750 -3600
rect 1910 -3610 3030 -3600
rect 1910 -3640 2850 -3610
rect 1300 -3690 2850 -3640
rect 1300 -3720 1550 -3690
rect 1220 -3740 1300 -3730
rect 1530 -3730 1550 -3720
rect 1710 -3730 2850 -3690
rect 3010 -3730 3030 -3610
rect 1530 -3750 3030 -3730
rect 1420 -3770 1500 -3760
rect 1420 -3830 1430 -3770
rect 1490 -3790 1500 -3770
rect 2303 -3790 2309 -3789
rect 1490 -3830 2309 -3790
rect 1420 -3840 2309 -3830
rect 2303 -3841 2309 -3840
rect 2361 -3841 2367 -3789
rect 610 -3870 810 -3850
rect 610 -3970 630 -3870
rect 790 -3970 1610 -3870
rect 1650 -3880 1870 -3870
rect 1650 -3960 1790 -3880
rect 1650 -3970 1870 -3960
rect 610 -3990 810 -3970
rect 1420 -4010 1670 -4000
rect 1420 -4070 1430 -4010
rect 1490 -4050 1670 -4010
rect 2120 -4010 3030 -4000
rect 1490 -4070 1500 -4050
rect 1420 -4080 1500 -4070
rect 2120 -4070 2140 -4010
rect 2700 -4020 3030 -4010
rect 2700 -4070 2850 -4020
rect 2120 -4080 2850 -4070
rect 1220 -4100 1300 -4090
rect 1220 -4170 1230 -4100
rect 1530 -4110 1740 -4090
rect 1530 -4120 1550 -4110
rect 1300 -4150 1550 -4120
rect 1710 -4150 1740 -4110
rect 2730 -4110 2850 -4080
rect 1300 -4170 1740 -4150
rect 1860 -4170 2620 -4120
rect 890 -4200 1090 -4180
rect 1860 -4200 1900 -4170
rect 2730 -4200 2740 -4110
rect 890 -4300 910 -4200
rect 1070 -4300 1900 -4200
rect 1930 -4210 2210 -4200
rect 1930 -4290 1940 -4210
rect 2020 -4290 2210 -4210
rect 1930 -4300 2210 -4290
rect 2630 -4300 2740 -4200
rect 890 -4320 1090 -4300
rect 1860 -4330 1900 -4300
rect 1220 -4400 1230 -4330
rect 1300 -4350 1740 -4330
rect 1300 -4390 1550 -4350
rect 1710 -4390 1740 -4350
rect 1860 -4380 2620 -4330
rect 1220 -4410 1300 -4400
rect 1530 -4410 1740 -4390
rect 2730 -4390 2740 -4300
rect 2800 -4390 2850 -4110
rect 2730 -4420 2850 -4390
rect 1420 -4430 1500 -4420
rect 1420 -4490 1430 -4430
rect 1490 -4450 1500 -4430
rect 2120 -4430 2850 -4420
rect 1490 -4490 1670 -4450
rect 1420 -4500 1670 -4490
rect 2120 -4490 2140 -4430
rect 2700 -4480 2850 -4430
rect 3010 -4480 3030 -4020
rect 2700 -4490 3030 -4480
rect 2120 -4500 3030 -4490
rect 290 -4530 490 -4510
rect 290 -4630 310 -4530
rect 470 -4630 1610 -4530
rect 1650 -4540 1870 -4530
rect 1650 -4620 1790 -4540
rect 1650 -4630 1870 -4620
rect 290 -4650 490 -4630
rect 2303 -4660 2309 -4659
rect 1420 -4670 2309 -4660
rect 1420 -4730 1430 -4670
rect 1490 -4710 2309 -4670
rect 1490 -4730 1500 -4710
rect 2303 -4711 2309 -4710
rect 2361 -4711 2367 -4659
rect 1420 -4740 1500 -4730
rect 1220 -4760 1300 -4750
rect 1220 -4830 1230 -4760
rect 1530 -4770 3030 -4750
rect 1530 -4780 1550 -4770
rect 1300 -4810 1550 -4780
rect 1710 -4810 2850 -4770
rect 1300 -4830 2850 -4810
rect 2830 -4890 2850 -4830
rect 3010 -4890 3030 -4770
rect 5890 -4780 5900 -2500
rect 5960 -4740 5970 -2500
rect 6090 -4740 6190 -4710
rect 6310 -4740 6320 -1430
rect 5960 -4780 6320 -4740
rect 6380 -4780 6570 -1430
rect 5890 -4870 6570 -4780
rect 6730 -4870 6750 -1340
rect 5890 -4890 6750 -4870
rect 2830 -4910 3030 -4890
rect 870 -5920 6220 -5900
rect 870 -5990 890 -5920
rect 6200 -5990 6220 -5920
rect 870 -6010 6220 -5990
rect 6800 -6040 6890 -6020
rect 270 -6070 750 -6050
rect 270 -7240 290 -6070
rect 730 -7240 750 -6070
rect 270 -7260 750 -7240
rect 870 -7300 6220 -7280
rect 870 -7370 890 -7300
rect 6200 -7370 6220 -7300
rect 870 -7390 6220 -7370
rect 870 -7720 6220 -7700
rect 870 -7790 890 -7720
rect 6200 -7790 6220 -7720
rect 870 -7810 6220 -7790
rect 3390 -7840 3630 -7810
rect 280 -10500 750 -7860
rect 2880 -7880 3350 -7860
rect 2880 -9020 2900 -7880
rect 3330 -9020 3350 -7880
rect 2880 -9040 3350 -9020
rect 3390 -9070 3420 -7840
rect 3610 -9070 3630 -7840
rect 3680 -7880 4150 -7860
rect 3680 -9020 3700 -7880
rect 4130 -9020 4150 -7880
rect 3680 -9040 4150 -9020
rect 6280 -9040 6750 -6060
rect 6800 -7260 6810 -6040
rect 6870 -7260 6890 -6040
rect 6800 -7280 6890 -7260
rect 6800 -7840 6890 -7820
rect 3390 -9100 3630 -9070
rect 6800 -9060 6810 -7840
rect 6870 -9060 6890 -7840
rect 6800 -9080 6890 -9060
rect 980 -9120 6730 -9100
rect 980 -9250 1000 -9120
rect 6710 -9250 6730 -9120
rect 980 -9270 6730 -9250
rect 6800 -9300 6890 -9280
rect 6280 -9330 6750 -9320
rect 6280 -10490 6290 -9330
rect 6740 -10490 6750 -9330
rect 6280 -10500 6750 -10490
rect 6800 -10520 6810 -9300
rect 6870 -10520 6890 -9300
rect 6800 -10540 6890 -10520
rect 870 -10570 6220 -10550
rect 870 -10640 890 -10570
rect 6200 -10640 6220 -10570
rect 870 -10660 6220 -10640
<< via1 >>
rect 880 4650 940 4660
rect 880 4600 930 4650
rect 930 4600 940 4650
rect 850 4410 930 4420
rect 850 4370 880 4410
rect 880 4370 930 4410
rect 850 4350 930 4370
rect 440 4020 720 4180
rect 910 3850 1080 3950
rect 1180 3600 1470 3800
rect 1730 3620 2020 3780
rect 1570 3350 1650 3460
rect 2100 3350 2180 3460
rect 2330 3190 2390 3250
rect 2480 3190 2540 3250
rect 2644 3194 2696 3246
rect 2944 3194 2996 3246
rect 3134 3194 3186 3246
rect 3304 3194 3356 3246
rect 3464 3194 3516 3246
rect 3624 3194 3676 3246
rect 3764 3194 3816 3246
rect 3914 3194 3966 3246
rect 1240 2700 1350 2810
rect 1710 2580 1770 2640
rect 6280 3190 6340 3250
rect 6420 3190 6480 3250
rect 6808 3188 6868 3248
rect 6926 3188 6986 3248
rect 5414 2914 5466 2966
rect 630 1980 790 2520
rect 4910 2490 5030 2560
rect 5740 2430 5820 2510
rect 4060 2280 4240 2360
rect 5510 2280 5580 2360
rect 4910 2080 5030 2150
rect 1710 1860 1770 1920
rect 1240 1690 1350 1800
rect 1710 1570 1770 1630
rect 4630 1950 4810 2020
rect 4910 1820 5030 1890
rect 5629 1824 5681 1876
rect 4350 1550 4510 1630
rect 5510 1610 5580 1690
rect 310 970 470 1510
rect 4910 1410 5030 1480
rect 6570 1420 6730 2550
rect 4910 970 5030 1030
rect 1240 760 1350 870
rect 1710 850 1770 910
rect 5630 870 5690 930
rect 6000 900 6080 980
rect 1230 660 1300 730
rect 4070 750 4220 830
rect 5890 760 5970 820
rect 2650 640 2810 710
rect 5630 650 5690 710
rect 1360 570 1420 630
rect 2279 559 2331 611
rect 4910 550 5030 610
rect 630 160 790 510
rect 1780 150 1860 510
rect 4630 350 4810 440
rect 4910 170 5030 230
rect 1360 30 1420 90
rect 1230 -50 1290 10
rect 910 -190 1070 -100
rect 1230 -300 1290 -240
rect 2010 -230 2140 -50
rect 1360 -380 1420 -320
rect 310 -790 470 -440
rect 1780 -800 1860 -440
rect 2650 -440 2810 160
rect 5630 70 5690 130
rect 4350 -50 4510 30
rect 5890 -40 5970 20
rect 5630 -150 5690 -90
rect 4910 -250 5030 -190
rect 1360 -920 1420 -860
rect 2279 -901 2331 -849
rect 6570 -910 6730 1030
rect 1230 -1020 1300 -950
rect 2650 -1170 2810 -930
rect 1360 -1270 1420 -1210
rect 2279 -1281 2331 -1229
rect 630 -1490 790 -1330
rect 1690 -1500 1760 -1320
rect 4910 -1390 5030 -1330
rect 1360 -1610 1420 -1550
rect 1230 -1700 1300 -1630
rect 910 -1870 1070 -1720
rect 1230 -1980 1300 -1910
rect 1360 -2050 1420 -1990
rect 1900 -1960 1990 -1620
rect 310 -2270 470 -2110
rect 1690 -2280 1760 -2100
rect 2850 -2150 3010 -1430
rect 5630 -1490 5690 -1430
rect 5890 -1440 5970 -1380
rect 4070 -1610 4220 -1530
rect 5890 -1600 5970 -1540
rect 5630 -1710 5690 -1650
rect 4910 -1810 5030 -1750
rect 4630 -2020 4810 -1920
rect 4910 -2190 5030 -2130
rect 5630 -2290 5690 -2230
rect 1360 -2390 1420 -2330
rect 2279 -2371 2331 -2319
rect 1230 -2560 1300 -2400
rect 4350 -2410 4510 -2330
rect 5890 -2400 5970 -2340
rect 2850 -2550 3010 -2430
rect 5630 -2510 5690 -2450
rect 4910 -2610 5030 -2550
rect 1610 -2680 1680 -2620
rect 2309 -2691 2361 -2639
rect 630 -2840 790 -2700
rect 1970 -2810 2050 -2730
rect 1610 -2920 1680 -2860
rect 1230 -3010 1300 -2940
rect 910 -3140 1070 -3040
rect 1230 -3240 1300 -3170
rect 2140 -3170 2270 -3010
rect 1610 -3320 1680 -3260
rect 2850 -3310 3010 -2870
rect 310 -3460 470 -3360
rect 1970 -3450 2050 -3370
rect 1610 -3560 1680 -3500
rect 2304 -3541 2356 -3489
rect 1230 -3730 1300 -3580
rect 2850 -3730 3010 -3610
rect 1430 -3830 1490 -3770
rect 2309 -3841 2361 -3789
rect 630 -3970 790 -3870
rect 1790 -3960 1870 -3880
rect 1430 -4070 1490 -4010
rect 1230 -4170 1300 -4100
rect 910 -4300 1070 -4200
rect 1940 -4290 2020 -4210
rect 1230 -4400 1300 -4330
rect 1430 -4490 1490 -4430
rect 2850 -4480 3010 -4020
rect 310 -4630 470 -4530
rect 1790 -4620 1870 -4540
rect 1430 -4730 1490 -4670
rect 2309 -4711 2361 -4659
rect 1230 -4830 1300 -4760
rect 2850 -4890 3010 -4770
rect 6570 -4870 6730 -1340
rect 890 -5990 6200 -5920
rect 290 -7240 730 -6070
rect 890 -7370 6200 -7300
rect 890 -7790 6200 -7720
rect 2900 -9020 3330 -7880
rect 3420 -9070 3610 -7840
rect 3700 -9020 4130 -7880
rect 6810 -7260 6820 -6040
rect 6820 -7260 6870 -6040
rect 6810 -9060 6820 -7840
rect 6820 -9060 6870 -7840
rect 1000 -9250 6710 -9120
rect 6290 -10490 6740 -9330
rect 6810 -10520 6820 -9300
rect 6820 -10520 6870 -9300
rect 890 -10640 6200 -10570
<< metal2 >>
rect 870 4660 950 4670
rect 870 4600 880 4660
rect 940 4600 950 4660
rect 870 4440 950 4600
rect 840 4420 950 4440
rect 840 4350 850 4420
rect 930 4350 950 4420
rect 840 4340 950 4350
rect 420 4180 740 4200
rect 420 4020 440 4180
rect 720 4020 740 4180
rect 420 4000 740 4020
rect 890 3950 1100 3970
rect 890 3850 910 3950
rect 1080 3850 1100 3950
rect 890 3470 1100 3850
rect 1160 3800 1490 3820
rect 1160 3600 1180 3800
rect 1470 3600 1490 3800
rect 1710 3780 2040 3800
rect 1710 3620 1730 3780
rect 2020 3620 2040 3780
rect 1710 3600 2040 3620
rect 1160 3580 1490 3600
rect 890 3460 4820 3470
rect 890 3350 1570 3460
rect 1650 3350 2100 3460
rect 2180 3350 4820 3460
rect 890 3340 4820 3350
rect 610 2520 810 2540
rect 610 1980 630 2520
rect 790 1980 810 2520
rect 610 1960 810 1980
rect 290 1510 490 1530
rect 290 970 310 1510
rect 470 970 490 1510
rect 290 950 490 970
rect 610 510 810 530
rect 610 160 630 510
rect 790 160 810 510
rect 610 140 810 160
rect 890 -100 1090 3340
rect 2330 3250 2390 3256
rect 890 -190 910 -100
rect 1070 -190 1090 -100
rect 290 -440 490 -420
rect 290 -790 310 -440
rect 470 -790 490 -440
rect 290 -810 490 -790
rect 610 -1330 810 -1310
rect 610 -1490 630 -1330
rect 790 -1490 810 -1330
rect 610 -1510 810 -1490
rect 890 -1720 1090 -190
rect 890 -1870 910 -1720
rect 1070 -1870 1090 -1720
rect 290 -2110 490 -2090
rect 290 -2270 310 -2110
rect 470 -2270 490 -2110
rect 290 -2290 490 -2270
rect 610 -2700 810 -2680
rect 610 -2840 630 -2700
rect 790 -2840 810 -2700
rect 610 -2860 810 -2840
rect 890 -3040 1090 -1870
rect 890 -3140 910 -3040
rect 1070 -3140 1090 -3040
rect 290 -3360 490 -3340
rect 290 -3460 310 -3360
rect 470 -3460 490 -3360
rect 290 -3480 490 -3460
rect 610 -3870 810 -3850
rect 610 -3970 630 -3870
rect 790 -3970 810 -3870
rect 610 -3990 810 -3970
rect 890 -4200 1090 -3140
rect 890 -4300 910 -4200
rect 1070 -4300 1090 -4200
rect 290 -4530 490 -4510
rect 290 -4630 310 -4530
rect 470 -4630 490 -4530
rect 290 -4650 490 -4630
rect 890 -5000 1090 -4300
rect 1220 2810 1370 2830
rect 1220 2700 1240 2810
rect 1350 2700 1370 2810
rect 1220 1800 1370 2700
rect 2330 2640 2390 3190
rect 1700 2580 1710 2640
rect 1770 2580 2390 2640
rect 2480 3250 2540 3256
rect 2120 1920 2180 2580
rect 2480 2490 2540 3190
rect 2644 3246 2696 3252
rect 2644 3188 2696 3194
rect 2944 3246 2996 3252
rect 2944 3188 2996 3194
rect 3134 3246 3186 3252
rect 3134 3188 3186 3194
rect 3304 3246 3356 3252
rect 3304 3188 3356 3194
rect 3464 3246 3516 3252
rect 3464 3188 3516 3194
rect 3624 3246 3676 3252
rect 3624 3188 3676 3194
rect 3764 3246 3816 3252
rect 3764 3188 3816 3194
rect 3914 3246 3966 3252
rect 3914 3188 3966 3194
rect 1700 1860 1710 1920
rect 1770 1860 2180 1920
rect 2260 2430 2540 2490
rect 1220 1690 1240 1800
rect 1350 1690 1370 1800
rect 1220 870 1370 1690
rect 2260 1630 2320 2430
rect 2645 2275 2695 3188
rect 1700 1570 1710 1630
rect 1770 1570 2320 1630
rect 2455 2225 2695 2275
rect 2120 910 2180 1570
rect 1220 760 1240 870
rect 1350 760 1370 870
rect 1700 850 1710 910
rect 1770 850 2180 910
rect 1220 740 1370 760
rect 1220 730 1300 740
rect 1220 660 1230 730
rect 1220 10 1300 660
rect 1350 630 1430 640
rect 1350 570 1360 630
rect 1420 570 1430 630
rect 1350 90 1430 570
rect 2279 611 2331 617
rect 2455 610 2505 2225
rect 2630 710 2830 730
rect 2630 640 2650 710
rect 2810 640 2830 710
rect 2630 620 2830 640
rect 2331 560 2505 610
rect 2279 553 2331 559
rect 1770 510 2150 520
rect 1770 150 1780 510
rect 1860 150 2150 510
rect 1770 140 2150 150
rect 1350 30 1360 90
rect 1420 30 1430 90
rect 1350 20 1430 30
rect 1220 -50 1230 10
rect 1290 -50 1300 10
rect 1220 -240 1300 -50
rect 1220 -300 1230 -240
rect 1290 -300 1300 -240
rect 1220 -950 1300 -300
rect 2000 -50 2150 140
rect 2000 -230 2010 -50
rect 2140 -230 2150 -50
rect 1350 -320 1430 -310
rect 1350 -380 1360 -320
rect 1420 -380 1430 -320
rect 1350 -860 1430 -380
rect 2000 -430 2150 -230
rect 1770 -440 2150 -430
rect 1770 -800 1780 -440
rect 1860 -800 2150 -440
rect 2630 160 2830 180
rect 2630 -440 2650 160
rect 2810 -440 2830 160
rect 2630 -460 2830 -440
rect 1770 -810 2150 -800
rect 2945 -820 2995 3188
rect 1350 -920 1360 -860
rect 1420 -920 1430 -860
rect 2279 -849 2331 -843
rect 2520 -850 2995 -820
rect 2331 -870 2995 -850
rect 2331 -900 2570 -870
rect 2279 -907 2331 -901
rect 1350 -930 1430 -920
rect 2630 -930 2830 -910
rect 1220 -1020 1230 -950
rect 1220 -1630 1300 -1020
rect 2630 -1170 2650 -930
rect 2810 -1170 2830 -930
rect 2630 -1190 2830 -1170
rect 1350 -1210 1430 -1200
rect 1350 -1270 1360 -1210
rect 1420 -1270 1430 -1210
rect 1350 -1550 1430 -1270
rect 2279 -1229 2331 -1223
rect 3135 -1230 3185 3188
rect 2331 -1280 3185 -1230
rect 2279 -1287 2331 -1281
rect 1680 -1320 2000 -1310
rect 1680 -1500 1690 -1320
rect 1760 -1500 2000 -1320
rect 1680 -1510 2000 -1500
rect 1350 -1610 1360 -1550
rect 1420 -1610 1430 -1550
rect 1350 -1620 1430 -1610
rect 1890 -1620 2000 -1510
rect 1220 -1700 1230 -1630
rect 1220 -1910 1300 -1700
rect 1220 -1980 1230 -1910
rect 1890 -1960 1900 -1620
rect 1990 -1960 2000 -1620
rect 1220 -2400 1300 -1980
rect 1350 -1990 1430 -1980
rect 1350 -2050 1360 -1990
rect 1420 -2050 1430 -1990
rect 1350 -2330 1430 -2050
rect 1890 -2090 2000 -1960
rect 1680 -2100 2000 -2090
rect 1680 -2280 1690 -2100
rect 1760 -2280 2000 -2100
rect 2830 -1430 3030 -1410
rect 2830 -2150 2850 -1430
rect 3010 -2150 3030 -1430
rect 2830 -2170 3030 -2150
rect 1680 -2290 2000 -2280
rect 1350 -2390 1360 -2330
rect 1420 -2390 1430 -2330
rect 2279 -2319 2331 -2313
rect 3305 -2320 3355 3188
rect 2331 -2370 3355 -2320
rect 2279 -2377 2331 -2371
rect 1350 -2400 1430 -2390
rect 1220 -2560 1230 -2400
rect 1220 -2940 1300 -2560
rect 2830 -2430 3030 -2410
rect 2830 -2550 2850 -2430
rect 3010 -2550 3030 -2430
rect 2830 -2570 3030 -2550
rect 1600 -2680 1610 -2620
rect 1680 -2680 1690 -2620
rect 1600 -2860 1690 -2680
rect 2309 -2639 2361 -2633
rect 3465 -2640 3515 3188
rect 2361 -2690 3515 -2640
rect 2309 -2697 2361 -2691
rect 1960 -2730 2280 -2720
rect 1960 -2810 1970 -2730
rect 2050 -2810 2280 -2730
rect 1960 -2820 2280 -2810
rect 1600 -2920 1610 -2860
rect 1680 -2920 1690 -2860
rect 1220 -3010 1230 -2940
rect 1220 -3170 1300 -3010
rect 1220 -3240 1230 -3170
rect 1220 -3580 1300 -3240
rect 2130 -3010 2280 -2820
rect 2130 -3170 2140 -3010
rect 2270 -3170 2280 -3010
rect 1600 -3320 1610 -3260
rect 1680 -3320 1690 -3260
rect 1600 -3500 1690 -3320
rect 2130 -3360 2280 -3170
rect 2830 -2870 3030 -2850
rect 2830 -3310 2850 -2870
rect 3010 -3310 3030 -2870
rect 2830 -3330 3030 -3310
rect 1960 -3370 2280 -3360
rect 1960 -3450 1970 -3370
rect 2050 -3450 2280 -3370
rect 1960 -3460 2280 -3450
rect 1600 -3560 1610 -3500
rect 1680 -3560 1690 -3500
rect 2304 -3489 2356 -3483
rect 3625 -3490 3675 3188
rect 2356 -3540 3675 -3490
rect 2304 -3547 2356 -3541
rect 1220 -3730 1230 -3580
rect 1220 -4100 1300 -3730
rect 2830 -3610 3030 -3590
rect 2830 -3730 2850 -3610
rect 3010 -3730 3030 -3610
rect 2830 -3750 3030 -3730
rect 1420 -3770 1500 -3760
rect 1420 -3830 1430 -3770
rect 1490 -3830 1500 -3770
rect 1420 -4010 1500 -3830
rect 2309 -3789 2361 -3783
rect 3765 -3790 3815 3188
rect 2361 -3840 3815 -3790
rect 2309 -3847 2361 -3841
rect 1780 -3880 2030 -3870
rect 1780 -3960 1790 -3880
rect 1870 -3960 2030 -3880
rect 1780 -3970 2030 -3960
rect 1420 -4070 1430 -4010
rect 1490 -4070 1500 -4010
rect 1420 -4080 1500 -4070
rect 1220 -4170 1230 -4100
rect 1220 -4330 1300 -4170
rect 1220 -4400 1230 -4330
rect 1220 -4760 1300 -4400
rect 1930 -4210 2030 -3970
rect 1930 -4290 1940 -4210
rect 2020 -4290 2030 -4210
rect 1420 -4430 1500 -4420
rect 1420 -4490 1430 -4430
rect 1490 -4490 1500 -4430
rect 1420 -4670 1500 -4490
rect 1930 -4530 2030 -4290
rect 2830 -4020 3030 -4000
rect 2830 -4480 2850 -4020
rect 3010 -4480 3030 -4020
rect 2830 -4500 3030 -4480
rect 1780 -4540 2030 -4530
rect 1780 -4620 1790 -4540
rect 1870 -4620 2030 -4540
rect 1780 -4630 2030 -4620
rect 1420 -4730 1430 -4670
rect 1490 -4730 1500 -4670
rect 2309 -4659 2361 -4653
rect 3915 -4660 3965 3188
rect 4050 2360 4250 2370
rect 4050 2280 4060 2360
rect 4240 2280 4250 2360
rect 4050 2270 4250 2280
rect 4620 2020 4820 3340
rect 6280 3250 6340 3256
rect 4620 1950 4630 2020
rect 4810 1950 4820 2020
rect 4330 1630 4530 1650
rect 4330 1550 4350 1630
rect 4510 1550 4530 1630
rect 4330 1530 4530 1550
rect 4050 830 4250 850
rect 4050 750 4070 830
rect 4230 750 4250 830
rect 4050 730 4250 750
rect 4620 440 4820 1950
rect 4620 350 4630 440
rect 4810 350 4820 440
rect 4330 30 4530 50
rect 4330 -50 4350 30
rect 4510 -50 4530 30
rect 4330 -70 4530 -50
rect 4050 -1530 4250 -1510
rect 4050 -1610 4070 -1530
rect 4230 -1610 4250 -1530
rect 4050 -1630 4250 -1610
rect 4620 -1920 4820 350
rect 4620 -2020 4630 -1920
rect 4810 -2020 4820 -1920
rect 4330 -2330 4530 -2310
rect 4330 -2410 4350 -2330
rect 4510 -2410 4530 -2330
rect 4330 -2430 4530 -2410
rect 2361 -4710 3965 -4660
rect 2309 -4717 2361 -4711
rect 1420 -4740 1500 -4730
rect 1220 -4830 1230 -4760
rect 1220 -4840 1300 -4830
rect 2830 -4770 3030 -4750
rect 2830 -4890 2850 -4770
rect 3010 -4890 3030 -4770
rect 2830 -4910 3030 -4890
rect 4620 -5000 4820 -2020
rect 4900 3149 5040 3160
rect 4900 3031 4911 3149
rect 5029 3031 5040 3149
rect 4900 2560 5040 3031
rect 5414 2966 5466 2972
rect 5414 2908 5466 2914
rect 5415 2715 5465 2908
rect 4900 2490 4910 2560
rect 5030 2490 5040 2560
rect 4900 2150 5040 2490
rect 4900 2080 4910 2150
rect 5030 2080 5040 2150
rect 4900 1890 5040 2080
rect 5075 2665 5465 2715
rect 5075 1965 5125 2665
rect 5730 2510 5830 2520
rect 5730 2430 5740 2510
rect 5820 2430 5830 2510
rect 5730 2370 5830 2430
rect 5500 2360 5830 2370
rect 5500 2280 5510 2360
rect 5580 2280 5830 2360
rect 5500 2270 5830 2280
rect 5075 1915 5680 1965
rect 4900 1820 4910 1890
rect 5030 1820 5040 1890
rect 5630 1876 5680 1915
rect 5623 1824 5629 1876
rect 5681 1824 5687 1876
rect 4900 1480 5040 1820
rect 5730 1700 5830 2270
rect 5500 1690 5830 1700
rect 5500 1610 5510 1690
rect 5580 1610 5830 1690
rect 5500 1600 5830 1610
rect 4900 1410 4910 1480
rect 5030 1410 5040 1480
rect 4900 1030 5040 1410
rect 6280 1300 6340 3190
rect 4900 970 4910 1030
rect 5030 970 5040 1030
rect 4900 610 5040 970
rect 5630 1240 6340 1300
rect 6420 3250 6480 3256
rect 5630 940 5690 1240
rect 6420 1170 6480 3190
rect 6808 3248 6868 3254
rect 6550 2550 6750 2570
rect 6550 1420 6570 2550
rect 6730 1420 6750 2550
rect 6550 1400 6750 1420
rect 5760 1110 6480 1170
rect 5620 930 5700 940
rect 5620 870 5630 930
rect 5690 870 5700 930
rect 5620 860 5700 870
rect 5630 720 5690 860
rect 5620 710 5700 720
rect 5620 650 5630 710
rect 5690 650 5700 710
rect 5620 640 5700 650
rect 4900 550 4910 610
rect 5030 550 5040 610
rect 4900 230 5040 550
rect 5760 270 5820 1110
rect 6550 1030 6750 1050
rect 4900 170 4910 230
rect 5030 170 5040 230
rect 4900 -190 5040 170
rect 5630 210 5820 270
rect 5880 980 6090 990
rect 5880 900 6000 980
rect 6080 900 6090 980
rect 5880 890 6090 900
rect 5880 820 5980 890
rect 5880 760 5890 820
rect 5970 760 5980 820
rect 5630 140 5690 210
rect 5620 130 5700 140
rect 5620 70 5630 130
rect 5690 70 5700 130
rect 5620 60 5700 70
rect 5630 -80 5690 60
rect 5880 20 5980 760
rect 5880 -40 5890 20
rect 5970 -40 5980 20
rect 5880 -50 5980 -40
rect 5620 -90 5700 -80
rect 5620 -150 5630 -90
rect 5690 -150 5700 -90
rect 5620 -160 5700 -150
rect 4900 -250 4910 -190
rect 5030 -250 5040 -190
rect 4900 -1330 5040 -250
rect 6550 -910 6570 1030
rect 6730 -910 6750 1030
rect 6550 -930 6750 -910
rect 6808 -1060 6868 3188
rect 4900 -1390 4910 -1330
rect 5030 -1390 5040 -1330
rect 4900 -1750 5040 -1390
rect 5630 -1120 6868 -1060
rect 6926 3248 6986 3254
rect 5630 -1420 5690 -1120
rect 6926 -1190 6986 3188
rect 5760 -1250 6986 -1190
rect 5620 -1430 5700 -1420
rect 5620 -1490 5630 -1430
rect 5690 -1490 5700 -1430
rect 5620 -1500 5700 -1490
rect 5630 -1640 5690 -1500
rect 5620 -1650 5700 -1640
rect 5620 -1710 5630 -1650
rect 5690 -1710 5700 -1650
rect 5620 -1720 5700 -1710
rect 4900 -1810 4910 -1750
rect 5030 -1810 5040 -1750
rect 4900 -2130 5040 -1810
rect 5760 -2090 5820 -1250
rect 6550 -1340 6750 -1320
rect 4900 -2190 4910 -2130
rect 5030 -2190 5040 -2130
rect 4900 -2550 5040 -2190
rect 5630 -2150 5820 -2090
rect 5880 -1380 5980 -1370
rect 5880 -1440 5890 -1380
rect 5970 -1440 5980 -1380
rect 5880 -1540 5980 -1440
rect 5880 -1600 5890 -1540
rect 5970 -1600 5980 -1540
rect 5630 -2220 5690 -2150
rect 5620 -2230 5700 -2220
rect 5620 -2290 5630 -2230
rect 5690 -2290 5700 -2230
rect 5620 -2300 5700 -2290
rect 5630 -2440 5690 -2300
rect 5880 -2340 5980 -1600
rect 5880 -2400 5890 -2340
rect 5970 -2400 5980 -2340
rect 5880 -2410 5980 -2400
rect 5620 -2450 5700 -2440
rect 5620 -2510 5630 -2450
rect 5690 -2510 5700 -2450
rect 5620 -2520 5700 -2510
rect 4900 -2610 4910 -2550
rect 5030 -2610 5040 -2550
rect 4900 -2620 5040 -2610
rect 6550 -4870 6570 -1340
rect 6730 -4870 6750 -1340
rect 5210 -5000 5430 -4990
rect 890 -5200 5216 -5000
rect 5416 -5200 5430 -5000
rect 5210 -5210 5430 -5200
rect 6550 -5820 6750 -4870
rect 860 -5920 6970 -5820
rect 860 -5990 890 -5920
rect 6200 -5990 6970 -5920
rect 860 -6020 6970 -5990
rect 6770 -6040 6970 -6020
rect 270 -6070 750 -6050
rect 270 -7240 290 -6070
rect 730 -7240 750 -6070
rect 270 -7260 750 -7240
rect 6770 -7260 6810 -6040
rect 6870 -7260 6970 -6040
rect 860 -7300 6970 -7260
rect 860 -7370 890 -7300
rect 6200 -7370 6970 -7300
rect 860 -7460 6970 -7370
rect 6783 -7643 6957 -7460
rect 853 -7720 6957 -7643
rect 853 -7790 890 -7720
rect 6200 -7790 6957 -7720
rect 853 -7817 6957 -7790
rect 3383 -7840 3640 -7817
rect 2880 -7880 3350 -7860
rect 2880 -9020 2900 -7880
rect 3330 -9020 3350 -7880
rect 2880 -9040 3350 -9020
rect 3383 -9070 3420 -7840
rect 3610 -9070 3640 -7840
rect 6783 -7840 6957 -7817
rect 3680 -7880 4150 -7860
rect 3680 -9020 3700 -7880
rect 4130 -9020 4150 -7880
rect 3680 -9040 4150 -9020
rect 3383 -9103 3640 -9070
rect 6783 -9060 6810 -7840
rect 6870 -9060 6957 -7840
rect 6783 -9103 6957 -9060
rect 963 -9120 6957 -9103
rect 963 -9250 1000 -9120
rect 6710 -9250 6957 -9120
rect 963 -9277 6957 -9250
rect 6783 -9300 6957 -9277
rect 6280 -9330 6750 -9320
rect 6280 -10490 6290 -9330
rect 6740 -10490 6750 -9330
rect 6280 -10500 6750 -10490
rect 6783 -10520 6810 -9300
rect 6870 -10520 6957 -9300
rect 6783 -10533 6957 -10520
rect 843 -10570 6957 -10533
rect 843 -10640 890 -10570
rect 6200 -10640 6957 -10570
rect 843 -10707 6957 -10640
<< via2 >>
rect 440 4020 720 4180
rect 1180 3600 1470 3800
rect 1730 3620 2020 3780
rect 630 1980 790 2520
rect 310 970 470 1510
rect 630 160 790 510
rect 310 -790 470 -440
rect 630 -1490 790 -1330
rect 310 -2270 470 -2110
rect 630 -2840 790 -2700
rect 310 -3460 470 -3360
rect 630 -3970 790 -3870
rect 310 -4630 470 -4530
rect 2650 640 2810 710
rect 2650 -440 2810 160
rect 2650 -1170 2810 -930
rect 2850 -2150 3010 -1430
rect 2850 -2550 3010 -2430
rect 2850 -3310 3010 -2870
rect 2850 -3730 3010 -3610
rect 2850 -4480 3010 -4020
rect 4060 2280 4240 2360
rect 4350 1550 4510 1630
rect 4070 750 4220 830
rect 4220 750 4230 830
rect 4350 -50 4510 30
rect 4070 -1610 4220 -1530
rect 4220 -1610 4230 -1530
rect 4350 -2410 4510 -2330
rect 2850 -4890 3010 -4770
rect 4911 3031 5029 3149
rect 6570 1420 6730 2550
rect 6570 -910 6730 1030
rect 6570 -4870 6730 -1340
rect 5216 -5200 5416 -5000
rect 290 -7240 730 -6070
rect 2900 -9020 3330 -7880
rect 3700 -9020 4130 -7880
rect 6290 -10490 6740 -9330
<< metal3 >>
rect 420 4180 740 4200
rect 420 4020 440 4180
rect 720 4020 740 4180
rect 420 3400 740 4020
rect 1160 3800 1490 3820
rect 1160 3600 1180 3800
rect 1470 3780 6750 3800
rect 1470 3620 1730 3780
rect 2020 3620 6750 3780
rect 1470 3600 6750 3620
rect 1160 3580 1490 3600
rect 420 3240 440 3400
rect 720 3240 740 3400
rect 420 3220 740 3240
rect 610 2520 810 2540
rect 610 1980 630 2520
rect 790 1980 810 2520
rect 290 1510 490 1530
rect 290 970 310 1510
rect 470 970 490 1510
rect 290 950 490 970
rect 610 510 810 1980
rect 610 160 630 510
rect 790 160 810 510
rect 290 -440 490 -420
rect 290 -790 310 -440
rect 470 -790 490 -440
rect 290 -810 490 -790
rect 610 -1330 810 160
rect 2630 710 2830 3600
rect 4906 3149 5034 3600
rect 4906 3031 4911 3149
rect 5029 3031 5034 3149
rect 4906 3026 5034 3031
rect 6550 2550 6750 3600
rect 2630 640 2650 710
rect 2810 640 2830 710
rect 2630 160 2830 640
rect 2630 -440 2650 160
rect 2810 -440 2830 160
rect 2630 -930 2830 -440
rect 2630 -1170 2650 -930
rect 2810 -1130 2830 -930
rect 4050 2360 4250 2370
rect 4050 2280 4060 2360
rect 4240 2280 4250 2360
rect 4050 830 4250 2280
rect 4330 1630 4530 1650
rect 4330 1550 4350 1630
rect 4510 1550 4530 1630
rect 4330 1530 4530 1550
rect 4050 750 4070 830
rect 4230 750 4250 830
rect 2810 -1170 3030 -1130
rect 2630 -1330 3030 -1170
rect 610 -1490 630 -1330
rect 790 -1490 810 -1330
rect 290 -2110 490 -2090
rect 290 -2270 310 -2110
rect 470 -2270 490 -2110
rect 290 -2290 490 -2270
rect 610 -2700 810 -1490
rect 610 -2840 630 -2700
rect 790 -2840 810 -2700
rect 290 -3360 490 -3340
rect 290 -3460 310 -3360
rect 470 -3460 490 -3360
rect 290 -3480 490 -3460
rect 610 -3870 810 -2840
rect 610 -3970 630 -3870
rect 790 -3970 810 -3870
rect 290 -4530 490 -4510
rect 290 -4630 310 -4530
rect 470 -4630 490 -4530
rect 290 -4650 490 -4630
rect 610 -5280 810 -3970
rect 2830 -1430 3030 -1330
rect 2830 -2150 2850 -1430
rect 3010 -2150 3030 -1430
rect 2830 -2430 3030 -2150
rect 2830 -2550 2850 -2430
rect 3010 -2550 3030 -2430
rect 2830 -2870 3030 -2550
rect 2830 -3310 2850 -2870
rect 3010 -3310 3030 -2870
rect 2830 -3610 3030 -3310
rect 2830 -3730 2850 -3610
rect 3010 -3730 3030 -3610
rect 2830 -4020 3030 -3730
rect 2830 -4480 2850 -4020
rect 3010 -4480 3030 -4020
rect 2830 -4770 3030 -4480
rect 2830 -4890 2850 -4770
rect 3010 -4890 3030 -4770
rect 2830 -4910 3030 -4890
rect 4050 -1530 4250 750
rect 6550 1420 6570 2550
rect 6730 1420 6750 2550
rect 6550 1030 6750 1420
rect 4330 30 4530 50
rect 4330 -50 4350 30
rect 4510 -50 4530 30
rect 4330 -70 4530 -50
rect 4050 -1610 4070 -1530
rect 4230 -1610 4250 -1530
rect 4050 -5280 4250 -1610
rect 6550 -910 6570 1030
rect 6730 -910 6750 1030
rect 6550 -1340 6750 -910
rect 4330 -2330 4530 -2310
rect 4330 -2410 4350 -2330
rect 4510 -2410 4530 -2330
rect 4330 -2430 4530 -2410
rect 6550 -4870 6570 -1340
rect 6730 -4870 6750 -1340
rect 6550 -4890 6750 -4870
rect 5210 -4995 5430 -4990
rect 5210 -5000 5221 -4995
rect 5210 -5200 5216 -5000
rect 5210 -5205 5221 -5200
rect 5421 -5205 5430 -4995
rect 5210 -5210 5430 -5205
rect 610 -5480 6970 -5280
rect 270 -6070 750 -6050
rect 270 -7240 290 -6070
rect 730 -7240 750 -6070
rect 270 -7260 750 -7240
rect 270 -7710 470 -7260
rect 0 -7730 470 -7710
rect 0 -7910 10 -7730
rect 190 -7910 470 -7730
rect 0 -7920 470 -7910
rect 2880 -7880 3350 -7860
rect 2880 -9020 2900 -7880
rect 3330 -9020 3350 -7880
rect 2880 -9040 3350 -9020
rect 3680 -7880 4150 -7860
rect 3680 -9020 3700 -7880
rect 4130 -9020 4150 -7880
rect 3680 -9040 4150 -9020
rect 6770 -9320 6970 -5480
rect 6280 -9330 6970 -9320
rect 6280 -10490 6290 -9330
rect 6740 -10490 6970 -9330
rect 6280 -10500 6770 -10490
rect 6770 -10696 6970 -10690
<< via3 >>
rect 440 4020 720 4180
rect 1180 3600 1470 3800
rect 440 3240 720 3400
rect 310 970 470 1510
rect 310 -790 470 -440
rect 4350 1550 4510 1630
rect 310 -2270 470 -2110
rect 310 -3460 470 -3360
rect 310 -4630 470 -4530
rect 4350 -50 4510 30
rect 4350 -2410 4510 -2330
rect 5221 -5000 5421 -4995
rect 5221 -5200 5416 -5000
rect 5416 -5200 5421 -5000
rect 5221 -5205 5421 -5200
rect 290 -7240 730 -6070
rect 10 -7910 190 -7730
rect 2900 -9020 3330 -7880
rect 3700 -9020 4130 -7880
rect 6770 -10690 6970 -10490
<< metal4 >>
rect 0 4180 740 4200
rect 0 4020 440 4180
rect 720 4020 740 4180
rect 0 4000 740 4020
rect 1160 3800 1490 3820
rect 0 3600 1180 3800
rect 1470 3600 1490 3800
rect 1160 3580 1490 3600
rect 0 3400 740 3420
rect 0 3240 440 3400
rect 720 3240 740 3400
rect 0 3220 740 3240
rect 0 -7450 200 3220
rect 4330 1630 4530 1650
rect 4330 1550 4350 1630
rect 4510 1550 4530 1630
rect 290 1510 490 1530
rect 290 970 310 1510
rect 470 970 490 1510
rect 290 -440 490 970
rect 290 -790 310 -440
rect 470 -790 490 -440
rect 290 -2110 490 -790
rect 290 -2270 310 -2110
rect 470 -2270 490 -2110
rect 290 -3360 490 -2270
rect 290 -3460 310 -3360
rect 470 -3460 490 -3360
rect 290 -4530 490 -3460
rect 290 -4630 310 -4530
rect 470 -4630 490 -4530
rect 290 -5560 490 -4630
rect 4330 30 4530 1550
rect 4330 -50 4350 30
rect 4510 -50 4530 30
rect 4330 -2330 4530 -50
rect 4330 -2410 4350 -2330
rect 4510 -2410 4530 -2330
rect 4330 -5560 4530 -2410
rect 5210 -4995 5430 -4990
rect 5210 -5205 5221 -4995
rect 5421 -5000 5430 -4995
rect 5421 -5200 6970 -5000
rect 5421 -5205 5430 -5200
rect 5210 -5210 5430 -5205
rect 290 -5760 4530 -5560
rect 290 -6050 490 -5760
rect 270 -6070 750 -6050
rect 270 -7240 290 -6070
rect 730 -7240 750 -6070
rect 270 -7260 750 -7240
rect 0 -7650 4010 -7450
rect 0 -7730 200 -7720
rect 0 -7910 10 -7730
rect 190 -7910 200 -7730
rect 3010 -7860 3210 -7650
rect 3810 -7860 4010 -7650
rect 0 -10950 200 -7910
rect 2880 -7880 3350 -7860
rect 2880 -9020 2900 -7880
rect 3330 -9020 3350 -7880
rect 2880 -9040 3350 -9020
rect 3680 -7880 4150 -7860
rect 3680 -9020 3700 -7880
rect 4130 -9020 4150 -7880
rect 3680 -9040 4150 -9020
rect 6769 -10490 6971 -10489
rect 6769 -10690 6770 -10490
rect 6970 -10690 6971 -10490
rect 6769 -10691 6971 -10690
rect 6770 -10950 6970 -10691
use sky130_fd_pr__nfet_01v8_ATLS57  sky130_fd_pr__nfet_01v8_ATLS57_0 csdac_nom__devices
timestamp 1723780759
transform -1 0 1651 0 -1 -620
box -211 -410 211 410
use sky130_fd_pr__nfet_01v8_HZS9GD  XMB0 csdac_nom__devices
timestamp 1723780759
transform 0 1 6140 -1 0 -3104
box -1796 -260 1796 260
use sky130_fd_pr__nfet_01v8_FMHZDY  XMB1 csdac_nom__devices
timestamp 1723780759
transform 0 1 6140 -1 0 56
box -996 -260 996 260
use sky130_fd_pr__nfet_01v8_AHZR5K  XMB2 csdac_nom__devices
timestamp 1723780759
transform 0 1 6030 -1 0 1986
box -596 -260 596 260
use sky130_fd_pr__nfet_01v8_BHEWB6  XMB3 csdac_nom__devices
timestamp 1723780759
transform 1 0 2416 0 1 -4250
box -406 -260 406 260
use sky130_fd_pr__nfet_01v8_FMMQLY  XMB4 csdac_nom__devices
timestamp 1723780759
transform 1 0 2486 0 1 -3090
box -296 -260 296 260
use sky130_fd_pr__nfet_01v8_C4RU6Y  XMB5 csdac_nom__devices
timestamp 1723780759
transform 1 0 2346 0 1 -1790
box -426 -400 426 400
use sky130_fd_pr__nfet_01v8_N5FCK4  XMB6 csdac_nom__devices
timestamp 1723780759
transform 1 0 2336 0 1 -140
box -246 -320 246 320
use sky130_fd_pr__nfet_01v8_8TEC39  XMB7 csdac_nom__devices
timestamp 1723780759
transform 0 -1 1860 1 0 3006
box -246 -420 246 420
use sky130_fd_pr__nfet_01v8_SMGLWN  XMmirror csdac_nom__devices
timestamp 1723780759
transform 1 0 1105 0 1 4507
box -246 -260 246 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMN0 csdac_nom__devices
timestamp 1723780759
transform 1 0 5421 0 1 -1570
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMN1
timestamp 1723780759
transform 1 0 5421 0 1 790
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMN2
timestamp 1723780759
transform 1 0 5381 0 1 2320
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMN3
timestamp 1723780759
transform 1 0 1631 0 1 -3920
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMN4
timestamp 1723780759
transform 1 0 1831 0 1 -2770
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_648S5X  XMN5 csdac_nom__devices
timestamp 1723780759
transform 1 0 1561 0 1 -1410
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_ATLS57  XMN6
timestamp 1723780759
transform -1 0 1651 0 -1 330
box -211 -410 211 410
use sky130_fd_pr__nfet_01v8_J2SMEF  XMN7 csdac_nom__devices
timestamp 1723780759
transform 1 0 1651 0 1 2250
box -211 -510 211 510
use sky130_fd_pr__nfet_01v8_L9ESAD  XMP0
timestamp 1723780759
transform 1 0 5421 0 1 -2370
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMP1
timestamp 1723780759
transform 1 0 5421 0 1 -10
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMP2
timestamp 1723780759
transform 1 0 5381 0 1 1650
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMP3
timestamp 1723780759
transform 1 0 1631 0 1 -4580
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMP4
timestamp 1723780759
transform 1 0 1831 0 1 -3410
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_648S5X  XMP5
timestamp 1723780759
transform 1 0 1561 0 1 -2190
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_J2SMEF  XMP7
timestamp 1723780759
transform 1 0 1651 0 1 1240
box -211 -510 211 510
use sky130_fd_pr__pfet_01v8_XJ7GBL  XMprog csdac_nom__devices
timestamp 1723780759
transform 1 0 631 0 1 4509
box -211 -269 211 269
use sky130_fd_pr__res_high_po_5p73_CS2QPW  XRLN csdac_nom__devices
timestamp 1724367708
transform 0 1 3512 -1 0 -9911
box -739 -3382 739 3382
use sky130_fd_pr__res_high_po_5p73_CS2QPW  XRLP
timestamp 1724367708
transform 0 1 3512 -1 0 -6651
box -739 -3382 739 3382
use sky130_fd_pr__res_high_po_5p73_69LTDJ  XRSN csdac_nom__devices
timestamp 1724367708
transform 0 1 1812 -1 0 -8451
box -739 -1682 739 1682
use sky130_fd_pr__res_high_po_5p73_69LTDJ  XRSP
timestamp 1724367708
transform 0 1 5212 -1 0 -8451
box -739 -1682 739 1682
<< labels >>
flabel metal4 0 4000 300 4200 0 FreeSans 1120 0 0 0 vcc
port 21 nsew
flabel metal4 0 3600 300 3800 0 FreeSans 1120 0 0 0 vss
port 22 nsew
flabel metal1 1850 950 2060 2950 0 FreeSans 800 0 0 0 IS7
flabel metal2 5880 -2340 5980 -1600 0 FreeSans 800 0 0 0 IS0
flabel metal2 5880 20 5980 760 0 FreeSans 800 0 0 0 IS1
flabel metal2 5580 2270 5830 2370 0 FreeSans 800 0 0 0 IS2
flabel metal1 1350 4920 1442 5196 0 FreeSans 640 0 0 0 n7
port 26 nsew
flabel metal1 3926 4920 4018 5196 0 FreeSans 640 0 0 0 p4
port 33 nsew
flabel metal1 4294 4920 4386 5196 0 FreeSans 640 0 0 0 n3
port 34 nsew
flabel metal1 4662 4920 4754 5196 0 FreeSans 640 0 0 0 p3
port 35 nsew
flabel metal1 5030 4920 5122 5196 0 FreeSans 640 0 0 0 n2
port 36 nsew
flabel metal1 5398 4920 5490 5196 0 FreeSans 640 0 0 0 p2
port 37 nsew
flabel metal1 6502 4920 6594 5196 0 FreeSans 640 0 0 0 n0
port 40 nsew
flabel metal1 6870 4920 6962 5196 0 FreeSans 640 0 0 0 p0
port 41 nsew
flabel metal1 6134 4920 6226 5196 0 FreeSans 640 0 0 0 p1
port 39 nsew
flabel metal1 5766 4920 5858 5196 0 FreeSans 640 0 0 0 n1
port 38 nsew
flabel metal1 3558 4920 3650 5196 0 FreeSans 640 0 0 0 n4
port 32 nsew
flabel metal1 3190 4920 3282 5196 0 FreeSans 640 0 0 0 p5
port 31 nsew
flabel metal1 2822 4920 2914 5196 0 FreeSans 640 0 0 0 n5
port 30 nsew
flabel metal1 2454 4920 2546 5196 0 FreeSans 640 0 0 0 p6
port 29 nsew
flabel metal1 2086 4920 2178 5196 0 FreeSans 640 0 0 0 n6
port 28 nsew
flabel metal1 1718 4920 1810 5196 0 FreeSans 640 0 0 0 p7
port 27 nsew
flabel metal2 2000 -50 2150 520 0 FreeSans 800 0 0 0 IS6
flabel metal2 1760 -1510 2000 -1310 0 FreeSans 800 0 0 0 IS5
flabel metal2 2130 -3010 2280 -2720 0 FreeSans 800 0 0 0 IS4
flabel metal2 1930 -4210 2030 -3870 0 FreeSans 800 0 0 0 IS3
flabel metal4 6770 -5200 6970 -5000 0 FreeSans 640 0 0 0 Vbias
port 42 nsew
flabel metal4 0 -10950 200 -10750 0 FreeSans 640 0 0 0 Vpos
port 44 nsew
flabel metal4 6770 -10950 6970 -10750 0 FreeSans 640 0 0 0 Vneg
port 43 nsew
<< end >>

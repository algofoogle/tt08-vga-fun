magic
tech sky130A
magscale 1 2
timestamp 1724131680
<< metal1 >>
rect 11648 18162 11654 18218
rect 11710 18162 11716 18218
rect 12016 18162 12022 18218
rect 12078 18162 12084 18218
rect 12384 18162 12390 18218
rect 12446 18162 12452 18218
rect 12752 18162 12758 18218
rect 12814 18162 12820 18218
rect 13120 18162 13126 18218
rect 13182 18162 13188 18218
rect 13488 18162 13494 18218
rect 13550 18162 13556 18218
rect 13856 18162 13862 18218
rect 13918 18162 13924 18218
rect 14224 18162 14230 18218
rect 14286 18162 14292 18218
rect 14592 18162 14598 18218
rect 14654 18162 14660 18218
rect 14960 18162 14966 18218
rect 15022 18162 15028 18218
rect 15328 18162 15334 18218
rect 15390 18162 15396 18218
rect 15696 18162 15702 18218
rect 15758 18162 15764 18218
rect 16064 18162 16070 18218
rect 16126 18162 16132 18218
rect 16432 18162 16438 18218
rect 16494 18162 16500 18218
rect 16800 18162 16806 18218
rect 16862 18162 16868 18218
rect 17168 18162 17174 18218
rect 17230 18162 17236 18218
<< via1 >>
rect 11654 18162 11710 18218
rect 12022 18162 12078 18218
rect 12390 18162 12446 18218
rect 12758 18162 12814 18218
rect 13126 18162 13182 18218
rect 13494 18162 13550 18218
rect 13862 18162 13918 18218
rect 14230 18162 14286 18218
rect 14598 18162 14654 18218
rect 14966 18162 15022 18218
rect 15334 18162 15390 18218
rect 15702 18162 15758 18218
rect 16070 18162 16126 18218
rect 16438 18162 16494 18218
rect 16806 18162 16862 18218
rect 17174 18162 17230 18218
<< metal2 >>
rect 10704 44870 10824 44900
rect 10704 44810 10732 44870
rect 10792 44810 10824 44870
rect 10704 44780 10824 44810
rect 11256 44870 11376 44900
rect 11256 44810 11284 44870
rect 11344 44810 11376 44870
rect 11256 44780 11376 44810
rect 11808 44870 11928 44900
rect 11808 44810 11836 44870
rect 11896 44810 11928 44870
rect 11808 44780 11928 44810
rect 12360 44870 12480 44900
rect 12360 44810 12388 44870
rect 12448 44810 12480 44870
rect 12360 44780 12480 44810
rect 12912 44870 13032 44900
rect 12912 44810 12940 44870
rect 13000 44810 13032 44870
rect 12912 44780 13032 44810
rect 13464 44870 13584 44900
rect 13464 44810 13492 44870
rect 13552 44810 13584 44870
rect 13464 44780 13584 44810
rect 14016 44870 14136 44900
rect 14016 44810 14044 44870
rect 14104 44810 14136 44870
rect 14016 44780 14136 44810
rect 14568 44870 14688 44900
rect 14568 44810 14596 44870
rect 14656 44810 14688 44870
rect 14568 44780 14688 44810
rect 15120 44870 15240 44900
rect 15120 44810 15148 44870
rect 15208 44810 15240 44870
rect 15120 44780 15240 44810
rect 15672 44870 15792 44900
rect 15672 44810 15700 44870
rect 15760 44810 15792 44870
rect 15672 44780 15792 44810
rect 20640 44870 20760 44900
rect 20640 44810 20668 44870
rect 20728 44810 20760 44870
rect 20640 44780 20760 44810
rect 21192 44870 21312 44900
rect 21192 44810 21220 44870
rect 21280 44810 21312 44870
rect 21192 44780 21312 44810
rect 21744 44870 21864 44900
rect 21744 44810 21772 44870
rect 21832 44810 21864 44870
rect 21744 44780 21864 44810
rect 22296 44870 22416 44900
rect 22296 44810 22324 44870
rect 22384 44810 22416 44870
rect 22296 44780 22416 44810
rect 22848 44870 22968 44900
rect 22848 44810 22876 44870
rect 22936 44810 22968 44870
rect 22848 44780 22968 44810
rect 23400 44870 23520 44900
rect 23400 44810 23428 44870
rect 23488 44810 23520 44870
rect 23400 44780 23520 44810
rect 23952 44870 24072 44900
rect 23952 44810 23980 44870
rect 24040 44810 24072 44870
rect 23952 44780 24072 44810
rect 24504 44870 24624 44900
rect 24504 44810 24532 44870
rect 24592 44810 24624 44870
rect 24504 44780 24624 44810
rect 25056 44870 25176 44900
rect 25056 44810 25084 44870
rect 25144 44810 25176 44870
rect 25056 44780 25176 44810
rect 25608 44870 25728 44900
rect 25608 44810 25636 44870
rect 25696 44810 25728 44870
rect 25608 44780 25728 44810
rect 10734 43862 10790 44780
rect 11286 43862 11342 44780
rect 11838 43862 11894 44780
rect 12390 43862 12446 44780
rect 12942 43862 12998 44780
rect 13494 43862 13550 44780
rect 14046 43862 14102 44780
rect 14598 43862 14654 44780
rect 15150 43862 15206 44780
rect 15702 43862 15758 44780
rect 20670 43862 20726 44780
rect 21222 43862 21278 44780
rect 21774 43862 21830 44780
rect 22326 43862 22382 44780
rect 22878 43862 22934 44780
rect 23430 43862 23486 44780
rect 23982 43862 24038 44780
rect 24534 43862 24590 44780
rect 25086 43862 25142 44780
rect 25638 43862 25694 44780
rect 11654 18218 11710 20148
rect 11654 18156 11710 18162
rect 12022 18218 12078 20148
rect 12022 18156 12078 18162
rect 12390 18218 12446 20148
rect 12390 18156 12446 18162
rect 12758 18218 12814 20148
rect 12758 18156 12814 18162
rect 13126 18218 13182 20148
rect 13126 18156 13182 18162
rect 13494 18218 13550 20148
rect 13494 18156 13550 18162
rect 13862 18218 13918 20148
rect 13862 18156 13918 18162
rect 14230 18218 14286 20148
rect 14230 18156 14286 18162
rect 14598 18218 14654 20148
rect 14598 18156 14654 18162
rect 14966 18218 15022 20148
rect 14966 18156 15022 18162
rect 15334 18218 15390 20148
rect 15334 18156 15390 18162
rect 15702 18218 15758 20148
rect 15702 18156 15758 18162
rect 16070 18218 16126 20148
rect 16070 18156 16126 18162
rect 16438 18218 16494 20148
rect 16438 18156 16494 18162
rect 16806 18218 16862 20148
rect 16806 18156 16862 18162
rect 17174 18218 17230 20148
rect 17174 18156 17230 18162
<< via2 >>
rect 10732 44810 10792 44870
rect 11284 44810 11344 44870
rect 11836 44810 11896 44870
rect 12388 44810 12448 44870
rect 12940 44810 13000 44870
rect 13492 44810 13552 44870
rect 14044 44810 14104 44870
rect 14596 44810 14656 44870
rect 15148 44810 15208 44870
rect 15700 44810 15760 44870
rect 20668 44810 20728 44870
rect 21220 44810 21280 44870
rect 21772 44810 21832 44870
rect 22324 44810 22384 44870
rect 22876 44810 22936 44870
rect 23428 44810 23488 44870
rect 23980 44810 24040 44870
rect 24532 44810 24592 44870
rect 25084 44810 25144 44870
rect 25636 44810 25696 44870
<< metal3 >>
rect 10704 44875 10824 44900
rect 6310 44798 6316 44862
rect 6380 44798 6386 44862
rect 6862 44798 6868 44862
rect 6932 44798 6938 44862
rect 10704 44805 10727 44875
rect 10797 44805 10824 44875
rect 926 44703 1074 44704
rect 921 44557 927 44703
rect 1073 44557 1079 44703
rect 926 44064 1074 44557
rect 6318 44408 6378 44798
rect 6870 44408 6930 44798
rect 10704 44780 10824 44805
rect 11256 44875 11376 44900
rect 11256 44805 11279 44875
rect 11349 44805 11376 44875
rect 11256 44780 11376 44805
rect 11808 44875 11928 44900
rect 11808 44805 11831 44875
rect 11901 44805 11928 44875
rect 11808 44780 11928 44805
rect 12360 44875 12480 44900
rect 12360 44805 12383 44875
rect 12453 44805 12480 44875
rect 12360 44780 12480 44805
rect 12912 44875 13032 44900
rect 12912 44805 12935 44875
rect 13005 44805 13032 44875
rect 12912 44780 13032 44805
rect 13464 44875 13584 44900
rect 13464 44805 13487 44875
rect 13557 44805 13584 44875
rect 13464 44780 13584 44805
rect 14016 44875 14136 44900
rect 14016 44805 14039 44875
rect 14109 44805 14136 44875
rect 14016 44780 14136 44805
rect 14568 44875 14688 44900
rect 14568 44805 14591 44875
rect 14661 44805 14688 44875
rect 14568 44780 14688 44805
rect 15120 44875 15240 44900
rect 15120 44805 15143 44875
rect 15213 44805 15240 44875
rect 15120 44780 15240 44805
rect 15672 44875 15792 44900
rect 15672 44805 15695 44875
rect 15765 44805 15792 44875
rect 15672 44780 15792 44805
rect 20640 44875 20760 44900
rect 20640 44805 20663 44875
rect 20733 44805 20760 44875
rect 20640 44780 20760 44805
rect 21192 44875 21312 44900
rect 21192 44805 21215 44875
rect 21285 44805 21312 44875
rect 21192 44780 21312 44805
rect 21744 44875 21864 44900
rect 21744 44805 21767 44875
rect 21837 44805 21864 44875
rect 21744 44780 21864 44805
rect 22296 44875 22416 44900
rect 22296 44805 22319 44875
rect 22389 44805 22416 44875
rect 22296 44780 22416 44805
rect 22848 44875 22968 44900
rect 22848 44805 22871 44875
rect 22941 44805 22968 44875
rect 22848 44780 22968 44805
rect 23400 44875 23520 44900
rect 23400 44805 23423 44875
rect 23493 44805 23520 44875
rect 23400 44780 23520 44805
rect 23952 44875 24072 44900
rect 23952 44805 23975 44875
rect 24045 44805 24072 44875
rect 23952 44780 24072 44805
rect 24504 44875 24624 44900
rect 24504 44805 24527 44875
rect 24597 44805 24624 44875
rect 24504 44780 24624 44805
rect 25056 44875 25176 44900
rect 25056 44805 25079 44875
rect 25149 44805 25176 44875
rect 25056 44780 25176 44805
rect 25608 44875 25728 44900
rect 25608 44805 25631 44875
rect 25701 44805 25728 44875
rect 25608 44780 25728 44805
rect 6316 44402 6380 44408
rect 6316 44332 6380 44338
rect 6868 44402 6932 44408
rect 6868 44332 6932 44338
rect 926 43910 1074 43916
rect 3789 19770 4187 19775
rect 200 19769 22190 19770
rect 200 19750 3789 19769
rect 200 19390 220 19750
rect 580 19390 3789 19750
rect 200 19371 3789 19390
rect 4187 19750 22190 19769
rect 4187 19390 9810 19750
rect 10170 19390 15810 19750
rect 16170 19390 21810 19750
rect 22170 19390 22190 19750
rect 4187 19371 22190 19390
rect 200 19370 22190 19371
rect 3789 19365 4187 19370
rect 801 19190 1199 19195
rect 800 19189 1980 19190
rect 800 18791 801 19189
rect 1199 18791 1980 19189
rect 800 18790 1980 18791
rect 2380 18790 2386 19190
rect 6783 18791 6789 19189
rect 7187 18791 7193 19189
rect 801 18785 1199 18790
rect 9120 17199 9320 19370
rect 12783 18791 12789 19189
rect 13187 18791 13193 19189
rect 18783 18791 18789 19189
rect 19187 18791 19193 19189
rect 24783 18791 24789 19189
rect 25187 18791 25193 19189
rect 9120 17001 9121 17199
rect 9319 17001 9320 17199
rect 9120 17000 9320 17001
rect 9121 16995 9319 17000
<< via3 >>
rect 6316 44798 6380 44862
rect 6868 44798 6932 44862
rect 10727 44870 10797 44875
rect 10727 44810 10732 44870
rect 10732 44810 10792 44870
rect 10792 44810 10797 44870
rect 10727 44805 10797 44810
rect 927 44557 1073 44703
rect 11279 44870 11349 44875
rect 11279 44810 11284 44870
rect 11284 44810 11344 44870
rect 11344 44810 11349 44870
rect 11279 44805 11349 44810
rect 11831 44870 11901 44875
rect 11831 44810 11836 44870
rect 11836 44810 11896 44870
rect 11896 44810 11901 44870
rect 11831 44805 11901 44810
rect 12383 44870 12453 44875
rect 12383 44810 12388 44870
rect 12388 44810 12448 44870
rect 12448 44810 12453 44870
rect 12383 44805 12453 44810
rect 12935 44870 13005 44875
rect 12935 44810 12940 44870
rect 12940 44810 13000 44870
rect 13000 44810 13005 44870
rect 12935 44805 13005 44810
rect 13487 44870 13557 44875
rect 13487 44810 13492 44870
rect 13492 44810 13552 44870
rect 13552 44810 13557 44870
rect 13487 44805 13557 44810
rect 14039 44870 14109 44875
rect 14039 44810 14044 44870
rect 14044 44810 14104 44870
rect 14104 44810 14109 44870
rect 14039 44805 14109 44810
rect 14591 44870 14661 44875
rect 14591 44810 14596 44870
rect 14596 44810 14656 44870
rect 14656 44810 14661 44870
rect 14591 44805 14661 44810
rect 15143 44870 15213 44875
rect 15143 44810 15148 44870
rect 15148 44810 15208 44870
rect 15208 44810 15213 44870
rect 15143 44805 15213 44810
rect 15695 44870 15765 44875
rect 15695 44810 15700 44870
rect 15700 44810 15760 44870
rect 15760 44810 15765 44870
rect 15695 44805 15765 44810
rect 20663 44870 20733 44875
rect 20663 44810 20668 44870
rect 20668 44810 20728 44870
rect 20728 44810 20733 44870
rect 20663 44805 20733 44810
rect 21215 44870 21285 44875
rect 21215 44810 21220 44870
rect 21220 44810 21280 44870
rect 21280 44810 21285 44870
rect 21215 44805 21285 44810
rect 21767 44870 21837 44875
rect 21767 44810 21772 44870
rect 21772 44810 21832 44870
rect 21832 44810 21837 44870
rect 21767 44805 21837 44810
rect 22319 44870 22389 44875
rect 22319 44810 22324 44870
rect 22324 44810 22384 44870
rect 22384 44810 22389 44870
rect 22319 44805 22389 44810
rect 22871 44870 22941 44875
rect 22871 44810 22876 44870
rect 22876 44810 22936 44870
rect 22936 44810 22941 44870
rect 22871 44805 22941 44810
rect 23423 44870 23493 44875
rect 23423 44810 23428 44870
rect 23428 44810 23488 44870
rect 23488 44810 23493 44870
rect 23423 44805 23493 44810
rect 23975 44870 24045 44875
rect 23975 44810 23980 44870
rect 23980 44810 24040 44870
rect 24040 44810 24045 44870
rect 23975 44805 24045 44810
rect 24527 44870 24597 44875
rect 24527 44810 24532 44870
rect 24532 44810 24592 44870
rect 24592 44810 24597 44870
rect 24527 44805 24597 44810
rect 25079 44870 25149 44875
rect 25079 44810 25084 44870
rect 25084 44810 25144 44870
rect 25144 44810 25149 44870
rect 25079 44805 25149 44810
rect 25631 44870 25701 44875
rect 25631 44810 25636 44870
rect 25636 44810 25696 44870
rect 25696 44810 25701 44870
rect 25631 44805 25701 44810
rect 6316 44338 6380 44402
rect 6868 44338 6932 44402
rect 926 43916 1074 44064
rect 220 19390 580 19750
rect 3789 19371 4187 19769
rect 9810 19390 10170 19750
rect 15810 19390 16170 19750
rect 21810 19390 22170 19750
rect 801 18791 1199 19189
rect 1980 18790 2380 19190
rect 6789 18791 7187 19189
rect 12789 18791 13187 19189
rect 18789 18791 19187 19189
rect 24789 18791 25187 19189
rect 9121 17001 9319 17199
<< metal4 >>
rect 926 44703 1074 44704
rect 926 44557 927 44703
rect 1073 44696 1074 44703
rect 3006 44696 3066 45152
rect 3558 44696 3618 45152
rect 4110 44696 4170 45152
rect 4662 44696 4722 45152
rect 5214 44696 5274 45152
rect 5766 44696 5826 45152
rect 6318 44863 6378 45152
rect 6870 44863 6930 45152
rect 6315 44862 6381 44863
rect 6315 44798 6316 44862
rect 6380 44798 6381 44862
rect 6315 44797 6381 44798
rect 6867 44862 6933 44863
rect 6867 44798 6868 44862
rect 6932 44798 6933 44862
rect 6867 44797 6933 44798
rect 7422 44696 7482 45152
rect 7974 44696 8034 45152
rect 8526 44696 8586 45152
rect 9078 44696 9138 45152
rect 9630 44696 9690 45152
rect 10182 44696 10242 45152
rect 10734 45010 10794 45152
rect 11286 45010 11346 45152
rect 11838 45010 11898 45152
rect 12390 45010 12450 45152
rect 12942 45010 13002 45152
rect 13494 45010 13554 45152
rect 14046 45010 14106 45152
rect 14598 45010 14658 45152
rect 15150 45010 15210 45152
rect 15702 45010 15762 45152
rect 10724 44900 10804 45010
rect 11276 44900 11356 45010
rect 11828 44900 11908 45010
rect 12380 44900 12460 45010
rect 12932 44900 13012 45010
rect 13484 44900 13564 45010
rect 14036 44900 14116 45010
rect 14588 44900 14668 45010
rect 15140 44900 15220 45010
rect 15692 44900 15772 45010
rect 16254 44952 16314 45152
rect 16806 44952 16866 45152
rect 17358 44952 17418 45152
rect 17910 44952 17970 45152
rect 18462 44952 18522 45152
rect 19014 44952 19074 45152
rect 19566 44952 19626 45152
rect 20118 44952 20178 45152
rect 20670 45010 20730 45152
rect 21222 45010 21282 45152
rect 21774 45010 21834 45152
rect 22326 45010 22386 45152
rect 22878 45010 22938 45152
rect 23430 45010 23490 45152
rect 23982 45010 24042 45152
rect 24534 45010 24594 45152
rect 25086 45010 25146 45152
rect 25638 45010 25698 45152
rect 20660 44900 20740 45010
rect 21212 44900 21292 45010
rect 21764 44900 21844 45010
rect 22316 44900 22396 45010
rect 22868 44900 22948 45010
rect 23420 44900 23500 45010
rect 23972 44900 24052 45010
rect 24524 44900 24604 45010
rect 25076 44900 25156 45010
rect 25628 44900 25708 45010
rect 26190 44952 26250 45152
rect 10704 44875 10824 44900
rect 10704 44805 10727 44875
rect 10797 44805 10824 44875
rect 10704 44780 10824 44805
rect 11256 44875 11376 44900
rect 11256 44805 11279 44875
rect 11349 44805 11376 44875
rect 11256 44780 11376 44805
rect 11808 44875 11928 44900
rect 11808 44805 11831 44875
rect 11901 44805 11928 44875
rect 11808 44780 11928 44805
rect 12360 44875 12480 44900
rect 12360 44805 12383 44875
rect 12453 44805 12480 44875
rect 12360 44780 12480 44805
rect 12912 44875 13032 44900
rect 12912 44805 12935 44875
rect 13005 44805 13032 44875
rect 12912 44780 13032 44805
rect 13464 44875 13584 44900
rect 13464 44805 13487 44875
rect 13557 44805 13584 44875
rect 13464 44780 13584 44805
rect 14016 44875 14136 44900
rect 14016 44805 14039 44875
rect 14109 44805 14136 44875
rect 14016 44780 14136 44805
rect 14568 44875 14688 44900
rect 14568 44805 14591 44875
rect 14661 44805 14688 44875
rect 14568 44780 14688 44805
rect 15120 44875 15240 44900
rect 15120 44805 15143 44875
rect 15213 44805 15240 44875
rect 15120 44780 15240 44805
rect 15672 44875 15792 44900
rect 15672 44805 15695 44875
rect 15765 44805 15792 44875
rect 15672 44780 15792 44805
rect 20640 44875 20760 44900
rect 20640 44805 20663 44875
rect 20733 44805 20760 44875
rect 20640 44780 20760 44805
rect 21192 44875 21312 44900
rect 21192 44805 21215 44875
rect 21285 44805 21312 44875
rect 21192 44780 21312 44805
rect 21744 44875 21864 44900
rect 21744 44805 21767 44875
rect 21837 44805 21864 44875
rect 21744 44780 21864 44805
rect 22296 44875 22416 44900
rect 22296 44805 22319 44875
rect 22389 44805 22416 44875
rect 22296 44780 22416 44805
rect 22848 44875 22968 44900
rect 22848 44805 22871 44875
rect 22941 44805 22968 44875
rect 22848 44780 22968 44805
rect 23400 44875 23520 44900
rect 23400 44805 23423 44875
rect 23493 44805 23520 44875
rect 23400 44780 23520 44805
rect 23952 44875 24072 44900
rect 23952 44805 23975 44875
rect 24045 44805 24072 44875
rect 23952 44780 24072 44805
rect 24504 44875 24624 44900
rect 24504 44805 24527 44875
rect 24597 44805 24624 44875
rect 24504 44780 24624 44805
rect 25056 44875 25176 44900
rect 25056 44805 25079 44875
rect 25149 44805 25176 44875
rect 25056 44780 25176 44805
rect 25608 44875 25728 44900
rect 25608 44805 25631 44875
rect 25701 44805 25728 44875
rect 25608 44780 25728 44805
rect 1073 44564 10316 44696
rect 1073 44557 1074 44564
rect 926 44556 1074 44557
rect 321 44442 479 44449
rect 321 44402 7092 44442
rect 321 44338 6316 44402
rect 6380 44338 6868 44402
rect 6932 44338 7092 44402
rect 321 44298 7092 44338
rect 321 44152 479 44298
rect 928 44152 1072 44160
rect 200 19750 600 44152
rect 200 19390 220 19750
rect 580 19390 600 19750
rect 200 1000 600 19390
rect 800 44064 1200 44152
rect 800 43916 926 44064
rect 1074 43916 1200 44064
rect 800 19189 1200 43916
rect 800 18791 801 19189
rect 1199 18791 1200 19189
rect 800 1000 1200 18791
rect 1400 1000 1800 44152
rect 3788 19769 4188 20880
rect 3788 19371 3789 19769
rect 4187 19371 4188 19769
rect 3788 19370 4188 19371
rect 1979 19190 2381 19191
rect 6788 19190 7188 20960
rect 9788 19750 10188 20880
rect 9788 19390 9810 19750
rect 10170 19390 10188 19750
rect 9788 19370 10188 19390
rect 12788 19190 13188 20960
rect 15788 19750 16188 20880
rect 15788 19390 15810 19750
rect 16170 19390 16188 19750
rect 15788 19370 16188 19390
rect 18788 19190 19188 20960
rect 21788 19750 22188 20880
rect 21788 19390 21810 19750
rect 22170 19390 22188 19750
rect 21788 19370 22188 19390
rect 24788 19190 25188 20960
rect 1979 18790 1980 19190
rect 2380 19189 25200 19190
rect 2380 18791 6789 19189
rect 7187 18791 12789 19189
rect 13187 18791 18789 19189
rect 19187 18791 24789 19189
rect 25187 18791 25200 19189
rect 2380 18790 25200 18791
rect 1979 18789 2381 18790
rect 8740 16800 8940 18790
rect 9120 17199 10040 17200
rect 9120 17001 9121 17199
rect 9319 17001 10040 17199
rect 9120 17000 10040 17001
rect 8740 16600 10050 16800
rect 20890 7330 27420 7530
rect 20930 6930 23560 7130
rect 20870 6530 21510 6730
rect 21310 6320 21510 6530
rect 19500 6120 21510 6320
rect 19518 200 19682 6120
rect 23376 200 23544 6930
rect 27238 200 27402 7330
rect 186 0 366 200
rect 4050 0 4230 200
rect 7914 0 8094 200
rect 11778 0 11958 200
rect 15642 0 15822 200
rect 19506 0 19686 200
rect 23370 0 23550 200
rect 27234 0 27414 200
use controller  controller_0
timestamp 1724102933
transform 1 0 2436 0 1 19984
box 386 0 23630 24000
use csdac_nom  green_dac
timestamp 1724037054
transform 1 0 9780 0 1 13000
box 0 -6470 11390 5396
<< labels >>
flabel metal4 s 25638 44952 25698 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 26190 44952 26250 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 27234 0 27414 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 23370 0 23550 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 19506 0 19686 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 15642 0 15822 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 11778 0 11958 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 7914 0 8094 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4050 0 4230 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 186 0 366 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 24534 44952 24594 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 23982 44952 24042 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 23430 44952 23490 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 22326 44952 22386 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 21774 44952 21834 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 21222 44952 21282 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 20118 44952 20178 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 19566 44952 19626 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 19014 44952 19074 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 17910 44952 17970 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 17358 44952 17418 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 16806 44952 16866 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 6870 44952 6930 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 6318 44952 6378 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 5766 44952 5826 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 4662 44952 4722 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 4110 44952 4170 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3558 44952 3618 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11286 44952 11346 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 10734 44952 10794 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10182 44952 10242 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 9078 44952 9138 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8526 44952 8586 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7974 44952 8034 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 15702 44952 15762 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 15150 44952 15210 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 14598 44952 14658 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 13494 44952 13554 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 12942 44952 13002 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 12390 44952 12450 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 1400 1000 1800 44152 1 FreeSans 400 0 0 0 VAPWR
port 53 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 29072 45152
<< end >>

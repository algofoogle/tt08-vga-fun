magic
tech sky130A
magscale 1 2
timestamp 1723353804
<< error_s >>
rect 17658 8263 17693 8297
rect 17659 8244 17693 8263
rect 298 1015 333 1032
rect 299 1014 333 1015
rect 299 978 369 1014
rect 129 947 187 953
rect 129 913 141 947
rect 316 944 387 978
rect 737 944 772 978
rect 129 907 187 913
rect 129 719 187 725
rect 129 685 141 719
rect 129 679 187 685
rect 316 583 386 944
rect 738 925 772 944
rect 316 547 369 583
rect 757 530 772 925
rect 791 891 826 925
rect 4276 891 4311 925
rect 791 530 825 891
rect 4277 872 4311 891
rect 791 496 806 530
rect 4296 477 4311 872
rect 4330 838 4365 872
rect 4645 838 4680 872
rect 4330 477 4364 838
rect 4646 819 4680 838
rect 4476 770 4534 776
rect 4476 736 4488 770
rect 4476 730 4534 736
rect 4476 560 4534 566
rect 4476 526 4488 560
rect 4476 520 4534 526
rect 4330 443 4345 477
rect 4665 424 4680 819
rect 4699 785 4734 819
rect 5014 785 5049 819
rect 4699 424 4733 785
rect 5015 766 5049 785
rect 4845 717 4903 723
rect 4845 683 4857 717
rect 4845 677 4903 683
rect 4845 507 4903 513
rect 4845 473 4857 507
rect 4845 467 4903 473
rect 4699 390 4714 424
rect 5034 371 5049 766
rect 5068 732 5103 766
rect 6953 732 6988 766
rect 5068 371 5102 732
rect 6954 713 6988 732
rect 5068 337 5083 371
rect 6973 318 6988 713
rect 7007 679 7042 713
rect 7322 679 7357 713
rect 7007 318 7041 679
rect 7323 660 7357 679
rect 7153 611 7211 617
rect 7153 577 7165 611
rect 7153 571 7211 577
rect 7153 401 7211 407
rect 7153 367 7165 401
rect 7153 361 7211 367
rect 7007 284 7022 318
rect 7342 265 7357 660
rect 7376 626 7411 660
rect 7691 626 7726 660
rect 7376 265 7410 626
rect 7692 607 7726 626
rect 7522 558 7580 564
rect 7522 524 7534 558
rect 7522 518 7580 524
rect 7522 348 7580 354
rect 7522 314 7534 348
rect 7522 308 7580 314
rect 7376 231 7391 265
rect 7711 212 7726 607
rect 7745 573 7780 607
rect 8830 573 8865 607
rect 7745 212 7779 573
rect 8831 554 8865 573
rect 7745 178 7760 212
rect 8850 159 8865 554
rect 8884 520 8919 554
rect 9199 520 9234 554
rect 8884 159 8918 520
rect 9200 501 9234 520
rect 9030 452 9088 458
rect 9030 418 9042 452
rect 9030 412 9088 418
rect 9030 242 9088 248
rect 9030 208 9042 242
rect 9030 202 9088 208
rect 8884 125 8899 159
rect 9219 106 9234 501
rect 9253 467 9288 501
rect 9568 467 9603 501
rect 9253 106 9287 467
rect 9569 448 9603 467
rect 9399 399 9457 405
rect 9399 365 9411 399
rect 9399 359 9457 365
rect 9399 189 9457 195
rect 9399 155 9411 189
rect 9399 149 9457 155
rect 9253 72 9268 106
rect 9588 53 9603 448
rect 9622 414 9657 448
rect 10327 414 10362 448
rect 9622 53 9656 414
rect 10328 395 10362 414
rect 9622 19 9637 53
rect 10347 0 10362 395
rect 10381 361 10416 395
rect 10696 361 10731 395
rect 10381 0 10415 361
rect 10697 342 10731 361
rect 10527 293 10585 299
rect 10527 259 10539 293
rect 10527 253 10585 259
rect 10527 83 10585 89
rect 10527 49 10539 83
rect 10527 43 10585 49
rect 10381 -34 10396 0
rect 10716 -53 10731 342
rect 10750 308 10785 342
rect 11065 308 11100 342
rect 10750 -53 10784 308
rect 11066 289 11100 308
rect 10896 240 10954 246
rect 10896 206 10908 240
rect 10896 200 10954 206
rect 10896 30 10954 36
rect 10896 -4 10908 30
rect 10896 -10 10954 -4
rect 10750 -87 10765 -53
rect 11085 -106 11100 289
rect 11119 255 11154 289
rect 11604 255 11639 289
rect 11119 -106 11153 255
rect 11605 236 11639 255
rect 11119 -140 11134 -106
rect 11624 -159 11639 236
rect 11658 202 11693 236
rect 11973 202 12008 236
rect 11658 -159 11692 202
rect 11974 183 12008 202
rect 11804 134 11862 140
rect 11804 100 11816 134
rect 11804 94 11862 100
rect 11804 -76 11862 -70
rect 11804 -110 11816 -76
rect 11804 -116 11862 -110
rect 11658 -193 11673 -159
rect 11993 -212 12008 183
rect 12027 149 12062 183
rect 12027 -212 12061 149
rect 12173 81 12231 87
rect 12173 47 12185 81
rect 12173 41 12231 47
rect 12173 -129 12231 -123
rect 12173 -163 12185 -129
rect 12173 -169 12231 -163
rect 12027 -246 12042 -212
rect 12362 -265 12377 183
rect 12396 -265 12430 237
rect 13142 177 13176 231
rect 15864 225 15899 259
rect 14687 184 14722 218
rect 15865 206 15899 225
rect 12396 -299 12411 -265
rect 13161 -318 13176 177
rect 13195 143 13230 177
rect 13510 143 13545 177
rect 14688 165 14722 184
rect 13195 -318 13229 143
rect 13511 124 13545 143
rect 13341 75 13399 81
rect 13341 41 13353 75
rect 13341 35 13399 41
rect 13341 -235 13399 -229
rect 13341 -269 13353 -235
rect 13341 -275 13399 -269
rect 13195 -352 13210 -318
rect 13530 -371 13545 124
rect 13564 90 13599 124
rect 13879 91 13914 124
rect 13564 -371 13598 90
rect 13710 22 13768 28
rect 13710 -12 13722 22
rect 13710 -18 13768 -12
rect 13710 -288 13768 -282
rect 13710 -322 13722 -288
rect 13710 -328 13768 -322
rect 13564 -405 13579 -371
rect 13899 -424 13914 91
rect 13933 57 13968 91
rect 13933 -424 13967 57
rect 13933 -458 13948 -424
rect 14338 -477 14353 91
rect 14372 -477 14406 145
rect 14518 116 14576 122
rect 14518 82 14530 116
rect 14518 76 14576 82
rect 14518 -394 14576 -388
rect 14518 -428 14530 -394
rect 14518 -434 14576 -428
rect 14372 -511 14387 -477
rect 14707 -530 14722 165
rect 14741 131 14776 165
rect 15056 132 15091 165
rect 14741 -530 14775 131
rect 14887 63 14945 69
rect 14887 29 14899 63
rect 14887 23 14945 29
rect 14887 -447 14945 -441
rect 14887 -481 14899 -447
rect 14887 -487 14945 -481
rect 14741 -564 14756 -530
rect 15076 -583 15091 132
rect 15110 98 15145 132
rect 15110 -583 15144 98
rect 15110 -617 15125 -583
rect 15515 -636 15530 132
rect 15549 -636 15583 186
rect 15695 157 15753 163
rect 15695 123 15707 157
rect 15695 117 15753 123
rect 15695 -553 15753 -547
rect 15695 -587 15707 -553
rect 15695 -593 15753 -587
rect 15549 -670 15564 -636
rect 15884 -689 15899 206
rect 15918 172 15953 206
rect 15918 -689 15952 172
rect 16064 104 16122 110
rect 16064 70 16076 104
rect 16064 64 16122 70
rect 16064 -606 16122 -600
rect 16064 -640 16076 -606
rect 16064 -646 16122 -640
rect 15918 -723 15933 -689
rect 16253 -742 16268 206
rect 16287 -742 16321 260
rect 16287 -776 16302 -742
rect 17678 -795 17693 8244
rect 17712 8210 17747 8244
rect 17712 -795 17746 8210
rect 17712 -829 17727 -795
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
rect 0 -4000 200 -3800
rect 0 -4400 200 -4200
rect 0 -4800 200 -4600
rect 0 -5200 200 -5000
rect 0 -5600 200 -5400
rect 0 -6000 200 -5800
rect 0 -6400 200 -6200
rect 0 -6800 200 -6600
rect 0 -7200 200 -7000
rect 0 -7600 200 -7400
rect 0 -8000 200 -7800
use csdac_nom__devices/sky130_fd_pr__nfet_01v8_HZS9GD  XMB0
timestamp 1723353804
transform 1 0 2551 0 1 701
box -1796 -260 1796 260
use csdac_nom__devices/sky130_fd_pr__nfet_01v8_FMHZDY  XMB1
timestamp 1723353804
transform 1 0 6028 0 1 542
box -996 -260 996 260
use csdac_nom__devices/sky130_fd_pr__nfet_01v8_AHZR5K  XMB2
timestamp 1723353804
transform 1 0 8305 0 1 383
box -596 -260 596 260
use csdac_nom__devices/sky130_fd_pr__nfet_01v8_BHEWB6  XMB3
timestamp 1723353804
transform 1 0 9992 0 1 224
box -406 -260 406 260
use csdac_nom__devices/sky130_fd_pr__nfet_01v8_FMMQLY  XMB4
timestamp 1723353804
transform 1 0 11379 0 1 65
box -296 -260 296 260
use csdac_nom__devices/sky130_fd_pr__nfet_01v8_C4RU6Y  XMB5
timestamp 1723353804
transform 1 0 12786 0 1 46
box -426 -400 426 400
use csdac_nom__devices/sky130_fd_pr__nfet_01v8_N5FCK4  XMB6
timestamp 1723353804
transform 1 0 14143 0 1 -193
box -246 -320 246 320
use csdac_nom__devices/sky130_fd_pr__nfet_01v8_8TEC39  XMB7
timestamp 1723353804
transform 1 0 15320 0 1 -252
box -246 -420 246 420
use csdac_nom__devices/sky130_fd_pr__nfet_01v8_SMGLWN  XMmirror
timestamp 1723353804
transform 1 0 562 0 1 754
box -246 -260 246 260
use csdac_nom__devices/sky130_fd_pr__nfet_01v8_L9ESAD  XMN0
timestamp 1723353804
transform 1 0 4874 0 1 595
box -211 -260 211 260
use csdac_nom__devices/sky130_fd_pr__nfet_01v8_L9ESAD  XMN1
timestamp 1723353804
transform 1 0 7551 0 1 436
box -211 -260 211 260
use csdac_nom__devices/sky130_fd_pr__nfet_01v8_L9ESAD  XMN2
timestamp 1723353804
transform 1 0 9428 0 1 277
box -211 -260 211 260
use csdac_nom__devices/sky130_fd_pr__nfet_01v8_L9ESAD  XMN3
timestamp 1723353804
transform 1 0 10925 0 1 118
box -211 -260 211 260
use csdac_nom__devices/sky130_fd_pr__nfet_01v8_L9ESAD  XMN4
timestamp 1723353804
transform 1 0 12202 0 1 -41
box -211 -260 211 260
use csdac_nom__devices/sky130_fd_pr__nfet_01v8_648S5X  XMN5
timestamp 1723353804
transform 1 0 13739 0 1 -150
box -211 -310 211 310
use csdac_nom__devices/sky130_fd_pr__nfet_01v8_ATLS57  XMN6
timestamp 1723353804
transform 1 0 14916 0 1 -209
box -211 -410 211 410
use csdac_nom__devices/sky130_fd_pr__nfet_01v8_J2SMEF  XMN7
timestamp 1723353804
transform 1 0 16093 0 1 -268
box -211 -510 211 510
use csdac_nom__devices/sky130_fd_pr__nfet_01v8_L9ESAD  XMP0
timestamp 1723353804
transform 1 0 4505 0 1 648
box -211 -260 211 260
use csdac_nom__devices/sky130_fd_pr__nfet_01v8_L9ESAD  XMP1
timestamp 1723353804
transform 1 0 7182 0 1 489
box -211 -260 211 260
use csdac_nom__devices/sky130_fd_pr__nfet_01v8_L9ESAD  XMP2
timestamp 1723353804
transform 1 0 9059 0 1 330
box -211 -260 211 260
use csdac_nom__devices/sky130_fd_pr__nfet_01v8_L9ESAD  XMP3
timestamp 1723353804
transform 1 0 10556 0 1 171
box -211 -260 211 260
use csdac_nom__devices/sky130_fd_pr__nfet_01v8_L9ESAD  XMP4
timestamp 1723353804
transform 1 0 11833 0 1 12
box -211 -260 211 260
use csdac_nom__devices/sky130_fd_pr__nfet_01v8_648S5X  XMP5
timestamp 1723353804
transform 1 0 13370 0 1 -97
box -211 -310 211 310
use csdac_nom__devices/sky130_fd_pr__nfet_01v8_ATLS57  XMP6
timestamp 1723353804
transform 1 0 14547 0 1 -156
box -211 -410 211 410
use csdac_nom__devices/sky130_fd_pr__nfet_01v8_J2SMEF  XMP7
timestamp 1723353804
transform 1 0 15724 0 1 -215
box -211 -510 211 510
use csdac_nom__devices/sky130_fd_pr__pfet_01v8_XJ7GBL  XMprog
timestamp 1723353804
transform 1 0 158 0 1 816
box -211 -269 211 269
use csdac_nom__devices/sky130_fd_pr__res_high_po_5p73_MRHKYZ  XR5
timestamp 1723353804
transform 1 0 16990 0 1 3751
box -739 -4582 739 4582
use csdac_nom__devices/sky130_fd_pr__res_high_po_5p73_MRHKYZ  XR6
timestamp 1723353804
transform 1 0 18415 0 1 3698
box -739 -4582 739 4582
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 vcc
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 vss
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 p0
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 n0
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 p1
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 n1
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 p2
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 n2
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 p3
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 n3
port 9 nsew
flabel metal1 0 -4000 200 -3800 0 FreeSans 256 0 0 0 p4
port 10 nsew
flabel metal1 0 -4400 200 -4200 0 FreeSans 256 0 0 0 n4
port 11 nsew
flabel metal1 0 -4800 200 -4600 0 FreeSans 256 0 0 0 p5
port 12 nsew
flabel metal1 0 -5200 200 -5000 0 FreeSans 256 0 0 0 n5
port 13 nsew
flabel metal1 0 -5600 200 -5400 0 FreeSans 256 0 0 0 p6
port 14 nsew
flabel metal1 0 -6000 200 -5800 0 FreeSans 256 0 0 0 n6
port 15 nsew
flabel metal1 0 -6400 200 -6200 0 FreeSans 256 0 0 0 p7
port 16 nsew
flabel metal1 0 -6800 200 -6600 0 FreeSans 256 0 0 0 n7
port 17 nsew
flabel metal1 0 -7200 200 -7000 0 FreeSans 256 0 0 0 Vpos
port 18 nsew
flabel metal1 0 -7600 200 -7400 0 FreeSans 256 0 0 0 Vneg
port 19 nsew
flabel metal1 0 -8000 200 -7800 0 FreeSans 256 0 0 0 Vbias
port 20 nsew
<< end >>

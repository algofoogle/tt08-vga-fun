magic
tech sky130A
magscale 1 2
timestamp 1725588957
<< error_s >>
rect 1840 5389 2020 5390
rect 1840 5171 1841 5389
rect 2019 5171 2020 5389
rect 1840 5170 2020 5171
rect 2450 5389 2630 5390
rect 2450 5171 2451 5389
rect 2629 5171 2630 5389
rect 2450 5170 2630 5171
rect 3060 5389 3240 5390
rect 3060 5171 3061 5389
rect 3239 5171 3240 5389
rect 3060 5170 3240 5171
rect -668 4299 -662 4300
rect -640 4271 -634 4300
rect 8775 408 8810 442
rect 11159 410 11194 444
rect 8776 389 8810 408
rect 11160 391 11194 410
rect 12336 391 12371 425
rect 8795 -106 8810 389
rect 8829 355 8864 389
rect 9214 355 9249 389
rect 8829 -106 8863 355
rect 9215 336 9249 355
rect 8829 -140 8844 -106
rect 9234 -159 9249 336
rect 9268 302 9303 336
rect 9268 -159 9302 302
rect 9268 -193 9283 -159
rect 9673 -212 9688 336
rect 9707 329 9742 363
rect 10022 329 10057 363
rect 9707 -212 9741 329
rect 10023 310 10057 329
rect 10975 342 11033 348
rect 9853 261 9911 267
rect 9853 227 9865 261
rect 9853 221 9911 227
rect 9853 -129 9911 -123
rect 9853 -163 9865 -129
rect 9853 -169 9911 -163
rect 9707 -246 9722 -212
rect 10042 -265 10057 310
rect 10076 276 10111 310
rect 10391 276 10426 310
rect 10076 -265 10110 276
rect 10392 257 10426 276
rect 10222 208 10280 214
rect 10222 174 10234 208
rect 10222 168 10280 174
rect 10222 -182 10280 -176
rect 10222 -216 10234 -182
rect 10222 -222 10280 -216
rect 10076 -299 10091 -265
rect 10411 -318 10426 257
rect 10445 223 10480 257
rect 10445 -318 10479 223
rect 10591 155 10649 161
rect 10591 121 10603 155
rect 10591 115 10649 121
rect 10591 -235 10649 -229
rect 10591 -269 10603 -235
rect 10591 -275 10649 -269
rect 10445 -352 10460 -318
rect 10780 -371 10795 257
rect 10814 -371 10848 311
rect 10975 308 10987 342
rect 10975 302 11033 308
rect 10975 -288 11033 -282
rect 10975 -322 10987 -288
rect 10975 -328 11033 -322
rect 10814 -405 10829 -371
rect 11179 -424 11194 391
rect 11213 357 11248 391
rect 11558 357 11593 391
rect 11213 -424 11247 357
rect 11559 338 11593 357
rect 11374 289 11432 295
rect 11374 255 11386 289
rect 11374 249 11432 255
rect 11374 -341 11432 -335
rect 11374 -375 11386 -341
rect 11374 -381 11432 -375
rect 11213 -458 11228 -424
rect 11578 -477 11593 338
rect 11612 304 11647 338
rect 11612 -477 11646 304
rect 11773 236 11831 242
rect 11773 202 11785 236
rect 11773 196 11831 202
rect 11773 -394 11831 -388
rect 11773 -428 11785 -394
rect 11773 -434 11831 -428
rect 11612 -511 11627 -477
rect 11977 -530 11992 338
rect 12011 -530 12045 391
rect 12337 372 12371 391
rect 12162 323 12220 329
rect 12162 289 12174 323
rect 12162 283 12220 289
rect 12162 -447 12220 -441
rect 12162 -481 12174 -447
rect 12162 -487 12220 -481
rect 12011 -564 12026 -530
rect 12356 -583 12371 372
rect 12390 338 12425 372
rect 12715 338 12750 372
rect 12390 -583 12424 338
rect 12716 319 12750 338
rect 12541 270 12599 276
rect 12541 236 12553 270
rect 12541 230 12599 236
rect 12541 -500 12599 -494
rect 12541 -534 12553 -500
rect 12541 -540 12599 -534
rect 12390 -617 12405 -583
rect 12735 -636 12750 319
rect 12769 285 12804 319
rect 12769 -636 12803 285
rect 12920 217 12978 223
rect 12920 183 12932 217
rect 12920 177 12978 183
rect 12920 -553 12978 -547
rect 12920 -587 12932 -553
rect 12920 -593 12978 -587
rect 12769 -670 12784 -636
<< viali >>
rect -1470 4720 -1420 4910
rect -510 4830 -450 4910
rect 320 4790 470 4830
rect 780 4790 880 4830
rect 1190 4800 1290 4840
rect -600 4310 -540 4390
rect 470 3890 620 4570
rect 980 3890 1130 4570
rect 1500 3920 1540 4640
rect 2260 4240 2300 4410
rect 2780 4240 2820 4410
rect 1650 4070 1700 4140
rect 2170 4080 2210 4140
rect 2870 4080 2910 4140
rect 3380 4070 3430 4140
rect -1280 3590 -1230 3860
rect 2200 3400 2280 3560
rect 2400 3420 2680 3480
rect 2820 3400 2900 3560
<< metal1 >>
rect 1510 5390 1680 5400
rect -1310 5380 -1190 5390
rect -1310 5280 -1300 5380
rect -1200 5280 -1190 5380
rect -1310 5270 -1190 5280
rect -1010 5380 -890 5390
rect -1010 5280 -1000 5380
rect -900 5280 -890 5380
rect 1510 5360 1520 5390
rect -1010 5270 -890 5280
rect 490 5270 1520 5360
rect -1300 4960 -1200 5270
rect -1010 5170 -670 5270
rect -1500 4910 -1310 4920
rect -1500 4720 -1470 4910
rect -1420 4820 -1310 4910
rect -1420 4720 -1400 4820
rect -1280 4740 -1230 4960
rect -1200 4820 -830 4920
rect -1500 3290 -1400 4720
rect -1170 4590 -1110 4820
rect -770 4740 -670 5170
rect 350 5170 430 5180
rect 350 5110 360 5170
rect 420 5110 430 5170
rect 490 5070 580 5270
rect 760 5170 840 5180
rect 760 5110 770 5170
rect 830 5110 840 5170
rect 772 5108 784 5110
rect 818 5108 830 5110
rect 772 5102 830 5108
rect 900 5070 990 5270
rect 1170 5180 1250 5190
rect 1170 5120 1180 5180
rect 1240 5120 1250 5180
rect 1182 5118 1194 5120
rect 1228 5118 1240 5120
rect 1182 5112 1240 5118
rect 1310 5080 1400 5270
rect 1510 5240 1520 5270
rect 1670 5240 1680 5390
rect 1510 5230 1680 5240
rect 1830 5390 2030 5400
rect 170 4980 370 5070
rect 420 4980 580 5070
rect -620 4910 -270 4920
rect -620 4830 -510 4910
rect -450 4830 -270 4910
rect -620 4820 -270 4830
rect -1220 4530 -1110 4590
rect -530 4540 -410 4550
rect -1220 4400 -1160 4530
rect -530 4500 -520 4540
rect -1100 4440 -520 4500
rect -420 4440 -410 4540
rect -1220 4300 -1120 4400
rect -1220 4060 -1160 4300
rect -950 4260 -870 4440
rect -530 4430 -410 4440
rect -370 4400 -270 4820
rect 170 4740 270 4980
rect 630 4970 780 5070
rect 822 5058 990 5070
rect 822 4982 828 5058
rect 830 4982 990 5058
rect 822 4980 990 4982
rect 1040 4980 1190 5080
rect 1232 5068 1400 5080
rect 1232 4992 1238 5068
rect 1240 4992 1400 5068
rect 1232 4980 1400 4992
rect 1830 5170 1840 5390
rect 2020 5170 2030 5390
rect 822 4970 840 4980
rect 350 4880 360 4940
rect 420 4880 430 4940
rect 350 4870 430 4880
rect 300 4830 520 4840
rect 300 4790 320 4830
rect 470 4790 520 4830
rect 300 4770 520 4790
rect 170 4640 340 4740
rect 240 4580 340 4640
rect 460 4590 520 4770
rect 630 4740 730 4970
rect 760 4880 770 4940
rect 830 4880 840 4940
rect 760 4870 840 4880
rect 760 4830 1010 4840
rect 760 4790 780 4830
rect 880 4790 1010 4830
rect 760 4770 1010 4790
rect 630 4640 850 4740
rect 750 4590 850 4640
rect 960 4590 1010 4770
rect 1040 4740 1140 4980
rect 1170 4890 1180 4950
rect 1240 4890 1250 4950
rect 1170 4880 1250 4890
rect 1170 4840 1560 4850
rect 1170 4800 1190 4840
rect 1290 4800 1560 4840
rect 1170 4780 1560 4800
rect 1040 4640 1360 4740
rect 1390 4680 1560 4780
rect -700 4390 -270 4400
rect -700 4310 -600 4390
rect -540 4310 -270 4390
rect -700 4300 -270 4310
rect 460 4570 630 4590
rect -1120 4210 -710 4260
rect -1220 4000 -1050 4060
rect -1500 3210 -1490 3290
rect -1410 3210 -1400 3290
rect -1500 3200 -1400 3210
rect -1310 3860 -1210 3880
rect -1310 3590 -1280 3860
rect -1230 3780 -1210 3860
rect -1110 3870 -1050 4000
rect -640 4040 -520 4300
rect -640 3914 -520 3920
rect 460 3890 470 4570
rect 620 3890 630 4570
rect 460 3870 630 3890
rect 970 4570 1140 4590
rect 1260 4580 1360 4640
rect 1480 4640 1560 4680
rect 970 3890 980 4570
rect 1130 3890 1140 4570
rect 1480 3990 1500 4640
rect 1540 4160 1560 4640
rect 1720 4280 1800 4290
rect 1720 4220 1730 4280
rect 1790 4220 1800 4280
rect 1720 4210 1800 4220
rect 1730 4190 1800 4210
rect 1830 4200 2030 5170
rect 2440 5390 2640 5400
rect 2440 5170 2450 5390
rect 2630 5170 2640 5390
rect 2170 4410 2320 4430
rect 2060 4280 2140 4290
rect 2060 4220 2070 4280
rect 2130 4220 2140 4280
rect 2060 4210 2140 4220
rect 2170 4240 2260 4410
rect 2300 4240 2320 4410
rect 1540 4140 1710 4160
rect 1540 4070 1650 4140
rect 1700 4070 1710 4140
rect 1740 4120 1800 4190
rect 2060 4190 2130 4210
rect 1540 4050 1710 4070
rect 1540 4000 1560 4050
rect 1540 3990 1590 4000
rect 1480 3900 1490 3990
rect 1580 3900 1590 3990
rect 1830 3960 2030 4130
rect 2060 4120 2120 4190
rect 2170 4170 2320 4240
rect 2170 4160 2190 4170
rect 2150 4140 2190 4160
rect 2150 4080 2170 4140
rect 2290 4120 2320 4170
rect 2350 4220 2410 4390
rect 2440 4370 2640 5170
rect 3050 5390 3250 5400
rect 3050 5170 3060 5390
rect 3240 5170 3250 5390
rect 2760 4410 2910 4430
rect 2350 4210 2430 4220
rect 2350 4150 2360 4210
rect 2420 4150 2430 4210
rect 2350 4140 2430 4150
rect 2150 4070 2190 4080
rect 2290 4070 2300 4120
rect 2150 4060 2300 4070
rect 1480 3890 1590 3900
rect 1660 3950 2030 3960
rect 970 3870 1140 3890
rect -1110 3810 -950 3870
rect 1660 3850 1670 3950
rect 1770 3850 2030 3950
rect 2480 3860 2600 4290
rect 2670 4220 2730 4390
rect 2650 4210 2730 4220
rect 2650 4150 2660 4210
rect 2720 4150 2730 4210
rect 2650 4140 2730 4150
rect 2760 4240 2780 4410
rect 2820 4240 2910 4410
rect 2760 4170 2910 4240
rect 2940 4280 3020 4290
rect 2940 4220 2950 4280
rect 3010 4220 3020 4280
rect 2940 4210 3020 4220
rect 2950 4190 3020 4210
rect 3050 4200 3250 5170
rect 3280 4280 3360 4290
rect 3280 4220 3290 4280
rect 3350 4220 3360 4280
rect 3280 4210 3360 4220
rect 2760 4120 2790 4170
rect 2890 4160 2910 4170
rect 2890 4140 2930 4160
rect 2780 4070 2790 4120
rect 2910 4080 2930 4140
rect 2960 4120 3020 4190
rect 3280 4190 3350 4210
rect 2890 4070 2930 4080
rect 2780 4060 2930 4070
rect 3050 3960 3250 4130
rect 3280 4120 3340 4190
rect 3370 4140 3450 4160
rect 3370 4070 3380 4140
rect 3430 4070 3450 4140
rect 3370 4050 3450 4070
rect 3050 3950 3420 3960
rect 1660 3840 2030 3850
rect 3050 3850 3310 3950
rect 3410 3850 3420 3950
rect 3050 3840 3420 3850
rect -1230 3680 -1120 3780
rect -1230 3590 -1210 3680
rect -1090 3650 3860 3810
rect -1110 3600 -950 3650
rect -1090 3590 -950 3600
rect 490 3590 600 3600
rect -1310 2690 -1210 3590
rect 240 3340 340 3570
rect 490 3500 500 3590
rect 590 3500 600 3590
rect 1000 3590 1110 3600
rect 490 3340 600 3500
rect 750 3340 850 3570
rect 1000 3500 1010 3590
rect 1100 3500 1110 3590
rect 1660 3580 1840 3600
rect 1000 3340 1110 3500
rect 1260 3480 1360 3570
rect 1660 3500 1680 3580
rect 1760 3500 1840 3580
rect 1660 3480 1840 3500
rect 1260 3470 1590 3480
rect 1260 3380 1490 3470
rect 1580 3380 1590 3470
rect 1920 3420 2040 3650
rect 2120 3590 2300 3600
rect 2120 3490 2190 3590
rect 2290 3540 2300 3590
rect 2780 3590 2960 3600
rect 2480 3540 2600 3560
rect 2780 3540 2790 3590
rect 2890 3560 2960 3590
rect 2290 3490 2790 3540
rect 2120 3480 2200 3490
rect 1260 3340 1590 3380
rect 2180 3400 2200 3480
rect 2280 3480 2820 3490
rect 2280 3420 2400 3480
rect 2680 3420 2820 3480
rect 2280 3400 2820 3420
rect 2900 3480 2960 3560
rect 2900 3400 2920 3480
rect 3060 3420 3180 3650
rect 3260 3580 3440 3600
rect 3260 3500 3340 3580
rect 3420 3500 3440 3580
rect 3260 3480 3440 3500
rect 2180 3360 2920 3400
rect 240 3210 1590 3340
rect -1310 2610 -1300 2690
rect -1220 2610 -1210 2690
rect -1310 2600 -1210 2610
rect 700 2690 900 3210
rect 700 2510 710 2690
rect 890 2510 900 2690
rect 700 2500 900 2510
rect 2320 2690 2760 3360
rect 2320 2310 2330 2690
rect 2750 2310 2760 2690
rect 2320 2300 2760 2310
rect 3700 2091 3860 3650
rect -1901 1929 3861 2091
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3600 200 -3400
rect 0 -4000 200 -3800
rect 0 -4400 200 -4200
rect 0 -4800 200 -4600
rect 0 -5200 200 -5000
rect 0 -5600 200 -5400
rect 0 -6000 200 -5800
rect 0 -6400 200 -6200
rect 0 -6800 200 -6600
rect 0 -7200 200 -7000
rect 2600 -7600 2800 -7400
<< via1 >>
rect -1300 5280 -1200 5380
rect -1000 5280 -900 5380
rect 360 5110 420 5170
rect 770 5110 830 5170
rect 1180 5120 1240 5180
rect 1520 5240 1670 5390
rect -520 4440 -420 4540
rect 1840 5170 2020 5390
rect 360 4880 420 4940
rect 770 4880 830 4940
rect 1180 4890 1240 4950
rect -1490 3210 -1410 3290
rect -640 3920 -520 4040
rect 500 3940 590 4030
rect 1010 3940 1100 4030
rect 1730 4220 1790 4280
rect 2450 5170 2630 5390
rect 2070 4220 2130 4280
rect 1490 3920 1500 3990
rect 1500 3920 1540 3990
rect 1540 3920 1580 3990
rect 1490 3900 1580 3920
rect 2190 4140 2290 4170
rect 2190 4080 2210 4140
rect 2210 4080 2290 4140
rect 3060 5170 3240 5390
rect 2360 4150 2420 4210
rect 2190 4070 2290 4080
rect 1670 3850 1770 3950
rect 2660 4150 2720 4210
rect 2950 4220 3010 4280
rect 3290 4220 3350 4280
rect 2790 4140 2890 4170
rect 2790 4080 2870 4140
rect 2870 4080 2890 4140
rect 2790 4070 2890 4080
rect 3310 3850 3410 3950
rect 500 3500 590 3590
rect 1010 3500 1100 3590
rect 1680 3500 1760 3580
rect 1490 3380 1580 3470
rect 2190 3560 2290 3590
rect 2190 3490 2200 3560
rect 2200 3490 2280 3560
rect 2280 3490 2290 3560
rect 2790 3560 2890 3590
rect 2790 3490 2820 3560
rect 2820 3490 2890 3560
rect 3340 3500 3420 3580
rect -1300 2610 -1220 2690
rect 710 2510 890 2690
rect 2330 2310 2750 2690
<< metal2 >>
rect 340 5500 440 5600
rect 750 5500 850 5600
rect 1160 5500 1260 5600
rect 1700 5500 1800 5600
rect 2050 5500 2150 5600
rect 2310 5500 2410 5600
rect -1310 5380 -1190 5390
rect -1310 5280 -1300 5380
rect -1200 5280 -1190 5380
rect -1310 5270 -1190 5280
rect -1010 5380 -890 5390
rect -1010 5280 -1000 5380
rect -900 5280 -890 5380
rect -1010 5270 -890 5280
rect 350 5170 430 5500
rect 350 5110 360 5170
rect 420 5110 430 5170
rect 350 4940 430 5110
rect 350 4880 360 4940
rect 420 4880 430 4940
rect 350 4870 430 4880
rect 760 5170 840 5500
rect 760 5110 770 5170
rect 830 5110 840 5170
rect 760 4940 840 5110
rect 760 4880 770 4940
rect 830 4880 840 4940
rect 1170 5180 1250 5500
rect 1510 5390 1680 5400
rect 1510 5240 1520 5390
rect 1670 5240 1680 5390
rect 1510 5230 1680 5240
rect 1170 5120 1180 5180
rect 1240 5120 1250 5180
rect 1170 4950 1250 5120
rect 1170 4890 1180 4950
rect 1240 4890 1250 4950
rect 1170 4880 1250 4890
rect 760 4870 840 4880
rect -530 4540 -410 4550
rect -530 4440 -520 4540
rect -420 4440 -410 4540
rect -530 4430 -410 4440
rect 1710 4290 1790 5500
rect 1830 5390 2030 5400
rect 1830 5170 1840 5390
rect 2020 5170 2030 5390
rect 1830 5160 2030 5170
rect 2060 4700 2140 5500
rect 2320 4850 2400 5500
rect 2440 5390 2640 5400
rect 2440 5170 2450 5390
rect 2630 5170 2640 5390
rect 2440 5160 2640 5170
rect 3050 5390 3250 5400
rect 3050 5170 3060 5390
rect 3240 5170 3250 5390
rect 3050 5160 3250 5170
rect 2320 4770 3020 4850
rect 2060 4620 2400 4700
rect 1710 4280 2140 4290
rect 1710 4220 1730 4280
rect 1790 4220 2070 4280
rect 2130 4220 2140 4280
rect 1710 4210 2140 4220
rect 2320 4220 2400 4620
rect 2940 4290 3020 4770
rect 2940 4280 3360 4290
rect 2940 4220 2950 4280
rect 3010 4220 3290 4280
rect 3350 4220 3360 4280
rect 2320 4210 2730 4220
rect 2940 4210 3360 4220
rect 2180 4170 2300 4180
rect 2180 4070 2190 4170
rect 2290 4070 2300 4170
rect 2330 4150 2360 4210
rect 2420 4150 2660 4210
rect 2720 4150 2730 4210
rect 2330 4140 2730 4150
rect 2780 4170 2900 4180
rect -646 3920 -640 4040
rect -520 3920 -514 4040
rect 490 4030 600 4040
rect 490 3940 500 4030
rect 590 3940 600 4030
rect -1500 3290 -1400 3300
rect -1500 3210 -1490 3290
rect -1410 3210 -1400 3290
rect -1500 3200 -1400 3210
rect -640 3290 -520 3920
rect 490 3590 600 3940
rect 490 3500 500 3590
rect 590 3500 600 3590
rect 490 3490 600 3500
rect 1000 4030 1110 4040
rect 1000 3940 1010 4030
rect 1100 3940 1110 4030
rect 1000 3590 1110 3940
rect 1000 3500 1010 3590
rect 1100 3500 1110 3590
rect 1000 3490 1110 3500
rect 1480 3990 1590 4000
rect 1480 3900 1490 3990
rect 1580 3900 1590 3990
rect 1480 3470 1590 3900
rect 1660 3950 1780 3960
rect 1660 3850 1670 3950
rect 1770 3850 1780 3950
rect 1660 3580 1780 3850
rect 1660 3500 1680 3580
rect 1760 3500 1780 3580
rect 1660 3480 1780 3500
rect 2180 3590 2300 4070
rect 2180 3490 2190 3590
rect 2290 3490 2300 3590
rect 2180 3480 2300 3490
rect 2780 4070 2790 4170
rect 2890 4070 2900 4170
rect 2780 3590 2900 4070
rect 3300 3950 3440 3960
rect 3300 3850 3310 3950
rect 3410 3850 3440 3950
rect 3300 3840 3440 3850
rect 2780 3490 2790 3590
rect 2890 3490 2900 3590
rect 2780 3480 2900 3490
rect 3320 3580 3440 3840
rect 3320 3500 3340 3580
rect 3420 3500 3440 3580
rect 3320 3480 3440 3500
rect 1480 3380 1490 3470
rect 1580 3380 1590 3470
rect 1480 3370 1590 3380
rect -640 3160 -630 3290
rect -530 3160 -520 3290
rect -640 3150 -520 3160
rect -1310 2690 -1210 2700
rect -1310 2610 -1300 2690
rect -1220 2610 -1210 2690
rect -1310 2600 -1210 2610
rect 700 2690 900 2700
rect 700 2510 710 2690
rect 890 2510 900 2690
rect 700 2500 900 2510
rect 2320 2690 2760 2700
rect 2320 2310 2330 2690
rect 2750 2310 2760 2690
rect 2320 2300 2760 2310
<< via2 >>
rect -1295 5285 -1205 5375
rect -995 5285 -905 5375
rect 1520 5240 1670 5390
rect -515 4445 -425 4535
rect 1840 5170 2020 5390
rect 2450 5170 2630 5390
rect 3060 5170 3240 5390
rect -1490 3210 -1410 3290
rect -630 3160 -530 3290
rect -1300 2610 -1220 2690
rect 710 2510 890 2690
rect 2330 2310 2750 2690
<< metal3 >>
rect -1300 5390 -1200 5600
rect -1000 5390 -900 5600
rect -700 5410 -600 5600
rect -1310 5375 -1190 5390
rect -1310 5285 -1295 5375
rect -1205 5285 -1190 5375
rect -1310 5270 -1190 5285
rect -1010 5375 -890 5390
rect -1010 5285 -995 5375
rect -905 5285 -890 5375
rect -700 5310 -420 5410
rect -1010 5270 -890 5285
rect -520 4550 -420 5310
rect 1510 5390 4160 5400
rect 1510 5240 1520 5390
rect 1670 5240 1840 5390
rect 1510 5170 1840 5240
rect 2020 5170 2450 5390
rect 2630 5170 3060 5390
rect 3240 5170 4160 5390
rect 1510 5160 4160 5170
rect -530 4535 -410 4550
rect -530 4445 -515 4535
rect -425 4445 -410 4535
rect -530 4430 -410 4445
rect -1500 3290 -1400 3300
rect -1500 3210 -1490 3290
rect -1410 3210 -1400 3290
rect -1500 3200 -1400 3210
rect -640 3290 -520 3300
rect -640 3160 -630 3290
rect -530 3160 -520 3290
rect -640 3150 -520 3160
rect -1310 2690 -1210 2700
rect -1310 2610 -1300 2690
rect -1220 2610 -1210 2690
rect -1310 2600 -1210 2610
rect 700 2690 900 2700
rect 700 2510 710 2690
rect 890 2510 900 2690
rect 700 2500 900 2510
rect 2320 2690 2760 2700
rect 2320 2310 2330 2690
rect 2750 2310 2760 2690
rect 2320 2300 2760 2310
rect 3920 -360 4160 5160
rect -1520 -1040 4160 -360
rect 3480 -1360 4160 -1040
<< via3 >>
rect 1840 5170 2020 5390
rect 2450 5170 2630 5390
rect 3060 5170 3240 5390
rect -1490 3210 -1410 3290
rect -630 3160 -530 3290
rect -1300 2610 -1220 2690
rect 710 2510 890 2690
rect 2330 2310 2750 2690
<< metal4 >>
rect -490 8280 5410 8590
rect -1900 3290 3680 3300
rect -1900 3210 -1490 3290
rect -1410 3210 -630 3290
rect -1900 3160 -630 3210
rect -530 3160 3680 3290
rect -1900 2900 3680 3160
rect -1900 2690 3680 2700
rect -1900 2610 -1300 2690
rect -1220 2610 710 2690
rect -1900 2510 710 2610
rect 890 2510 2330 2690
rect -1900 2310 2330 2510
rect 2750 2310 3680 2690
rect -1900 2300 3680 2310
rect 3300 -7600 3700 -7200
use sky130_fd_pr__pfet_01v8_JE7DK3  XM1
timestamp 1725517196
transform 1 0 -1254 0 1 4869
box -246 -269 246 269
use sky130_fd_pr__pfet_01v8_QBPJZQ  XM2
timestamp 1725517196
transform 1 0 -724 0 1 4869
box -296 -269 296 269
use sky130_fd_pr__pfet_01v8_8JDY5S  XM3
timestamp 1725517196
transform 1 0 -914 0 1 4349
box -396 -269 396 269
use sky130_fd_pr__nfet_01v8_DB7J7C  XMia1
timestamp 1725517196
transform 0 1 290 -1 0 4076
box -696 -260 696 260
use sky130_fd_pr__nfet_01v8_DB7J7C  XMia2
timestamp 1725517196
transform 0 1 800 -1 0 4076
box -696 -260 696 260
use sky130_fd_pr__nfet_01v8_DB7J7C  XMia3
timestamp 1725517196
transform 0 1 1310 -1 0 4076
box -696 -260 696 260
use sky130_fd_pr__nfet_01v8_33M553  XMib1
timestamp 1725517196
transform 1 0 1976 0 1 3540
box -316 -260 316 260
use sky130_fd_pr__nfet_01v8_33M553  XMib2
timestamp 1725517196
transform 0 1 2540 -1 0 3716
box -316 -260 316 260
use sky130_fd_pr__nfet_01v8_33M553  XMib3
timestamp 1725517196
transform 1 0 3116 0 1 3540
box -316 -260 316 260
use sky130_fd_pr__nfet_01v8_7DN82Q  XMic1
timestamp 1725517196
transform 1 0 8600 0 1 168
box -246 -310 246 310
use sky130_fd_pr__nfet_01v8_7DN82Q  XMic2
timestamp 1725517196
transform 1 0 9039 0 1 115
box -246 -310 246 310
use sky130_fd_pr__nfet_01v8_7DN82Q  XMic3
timestamp 1725517196
transform 1 0 9478 0 1 62
box -246 -310 246 310
use sky130_fd_pr__nfet_01v8_3ZUKNL  XMid1
timestamp 1725517196
transform 1 0 11004 0 1 10
box -226 -470 226 470
use sky130_fd_pr__nfet_01v8_3ZUKNL  XMid2
timestamp 1725517196
transform 1 0 11403 0 1 -43
box -226 -470 226 470
use sky130_fd_pr__nfet_01v8_3ZUKNL  XMid3
timestamp 1725517196
transform 1 0 11802 0 1 -96
box -226 -470 226 470
use sky130_fd_pr__nfet_01v8_VRHU84  XMmirror
timestamp 1725517196
transform 1 0 -1064 0 1 3730
box -246 -260 246 260
use sky130_fd_pr__nfet_01v8_AJ3M4R  XMsa1
timestamp 1725517196
transform 1 0 391 0 1 5020
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_AJ3M4R  XMsa2
timestamp 1725517196
transform 1 0 801 0 1 5020
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_AJ3M4R  XMsa3
timestamp 1725517196
transform 1 0 1211 0 1 5030
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_V8CAV6  XMsb1
timestamp 1725517196
transform 0 1 1930 -1 0 4161
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_V8CAV6  XMsb2
timestamp 1725517196
transform 0 1 2540 -1 0 4331
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_V8CAV6  XMsb3
timestamp 1725517196
transform 0 1 3150 -1 0 4161
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_V8CYR7  XMsc1
timestamp 1725517196
transform 1 0 9882 0 1 49
box -211 -350 211 350
use sky130_fd_pr__nfet_01v8_V8CYR7  XMsc2
timestamp 1725517196
transform 1 0 10251 0 1 -4
box -211 -350 211 350
use sky130_fd_pr__nfet_01v8_V8CYR7  XMsc3
timestamp 1725517196
transform 1 0 10620 0 1 -57
box -211 -350 211 350
use sky130_fd_pr__nfet_01v8_2BSVCH  XMsd1
timestamp 1725517196
transform 1 0 12191 0 1 -79
box -216 -540 216 540
use sky130_fd_pr__nfet_01v8_2BSVCH  XMsd2
timestamp 1725517196
transform 1 0 12570 0 1 -132
box -216 -540 216 540
use sky130_fd_pr__nfet_01v8_2BSVCH  XMsd3
timestamp 1725517196
transform 1 0 12949 0 1 -185
box -216 -540 216 540
<< labels >>
flabel metal1 0 -2400 200 -2200 0 FreeSans 1280 0 0 0 sb1
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 1280 0 0 0 sb2
port 7 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 1280 0 0 0 sb3
port 9 nsew
flabel metal1 0 -4000 200 -3800 0 FreeSans 1280 0 0 0 sc1
port 10 nsew
flabel metal1 0 -4400 200 -4200 0 FreeSans 1280 0 0 0 sc2
port 11 nsew
flabel metal1 0 -4800 200 -4600 0 FreeSans 1280 0 0 0 sc3
port 12 nsew
flabel metal1 0 -5200 200 -5000 0 FreeSans 1280 0 0 0 sd1
port 13 nsew
flabel metal1 0 -5600 200 -5400 0 FreeSans 1280 0 0 0 sd2
port 14 nsew
flabel metal1 0 -6000 200 -5800 0 FreeSans 1280 0 0 0 sd3
port 15 nsew
flabel metal1 0 -6400 200 -6200 0 FreeSans 1280 0 0 0 bias1
port 16 nsew
flabel metal1 0 -6800 200 -6600 0 FreeSans 1280 0 0 0 bias2
port 17 nsew
flabel metal1 0 -7200 200 -7000 0 FreeSans 1280 0 0 0 bias3
port 18 nsew
flabel metal4 3300 -7600 3700 -7200 0 FreeSans 1280 0 0 0 Vout
port 23 nsew
flabel metal1 2600 -7600 2800 -7400 0 FreeSans 1280 0 0 0 Vbias
port 8 nsew
flabel metal4 -1900 2900 -1500 3300 0 FreeSans 1600 0 0 0 vcc
port 19 nsew
flabel metal3 -1300 5500 -1200 5600 0 FreeSans 480 0 0 0 bias1
port 21 nsew
flabel metal3 -1000 5500 -900 5600 0 FreeSans 480 0 0 0 bias2
port 22 nsew
flabel metal3 -700 5500 -600 5600 0 FreeSans 480 0 0 0 bias3
port 24 nsew
flabel metal4 -1900 2300 -1500 2700 0 FreeSans 1600 0 0 0 vss
port 20 nsew
flabel metal2 340 5500 440 5600 0 FreeSans 480 0 0 0 sa1
port 25 nsew
flabel metal2 750 5500 850 5600 0 FreeSans 480 0 0 0 sa2
port 26 nsew
flabel metal2 1160 5500 1260 5600 0 FreeSans 480 0 0 0 sa3
port 27 nsew
flabel metal1 -1901 1929 -1739 2091 0 FreeSans 480 0 0 0 Vbias
port 28 nsew
flabel metal3 3480 -1360 4160 -680 0 FreeSans 1600 0 0 0 Vout
port 29 nsew
flabel metal2 1700 5500 1800 5600 0 FreeSans 480 0 0 0 sb1
port 30 nsew
flabel metal2 2050 5500 2150 5600 0 FreeSans 480 0 0 0 sb2
port 31 nsew
flabel metal2 2310 5500 2410 5600 0 FreeSans 480 0 0 0 sb3
port 32 nsew
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1724306358
<< pwell >>
rect 5780 1530 5860 1570
rect 5980 1540 6080 1590
rect 1360 -1760 1420 -1700
rect 1220 -2140 1310 -2050
rect 1230 -2710 1300 -2550
rect 1600 -2840 1690 -2770
rect 1600 -3070 1690 -3000
rect 1230 -3160 1300 -3090
rect 1230 -3390 1300 -3320
rect 1970 -3600 2050 -3520
rect 1230 -3880 1300 -3730
rect 1230 -4320 1300 -4250
rect 1230 -4550 1300 -4480
rect 1230 -4980 1300 -4910
<< locali >>
rect 880 4410 930 4420
<< viali >>
rect 540 4700 720 4750
rect 980 4690 1230 4740
rect 450 4360 500 4650
rect 880 4600 930 4650
rect 880 4370 930 4410
rect 1280 4370 1320 4640
rect 540 4270 720 4320
rect 1120 4280 1230 4320
rect 1720 3170 2030 3220
rect 1470 2880 1520 3130
rect 1570 2690 1770 2830
rect 5290 2500 5470 2550
rect 5900 2510 6160 2550
rect 5290 2090 5470 2140
rect 5300 1830 5460 1880
rect 1570 1680 1730 1810
rect 5800 1510 5840 1560
rect 6210 1510 6260 2460
rect 5300 1420 5460 1470
rect 5900 1420 6160 1460
rect 5340 970 5500 1020
rect 6160 980 6280 1030
rect 1570 750 1730 800
rect 1570 510 1740 570
rect 5340 560 5500 610
rect 5340 170 5500 220
rect 2220 -50 2460 0
rect 1570 -200 1740 -160
rect 1570 -430 1740 -390
rect 2500 -490 2560 -90
rect 5340 -240 5500 -190
rect 2220 -580 2460 -530
rect 5910 -810 5960 -140
rect 6320 -810 6380 920
rect 6010 -910 6270 -860
rect 1570 -1160 1740 -1100
rect 1480 -1330 1650 -1280
rect 5340 -1390 5500 -1340
rect 6030 -1380 6270 -1340
rect 2050 -1620 2660 -1570
rect 1480 -1850 1650 -1800
rect 1480 -2110 1650 -2060
rect 2690 -2230 2750 -1650
rect 5340 -1800 5500 -1750
rect 5340 -2190 5500 -2140
rect 2050 -2310 2660 -2260
rect 1480 -2620 1650 -2570
rect 5340 -2600 5500 -2550
rect 1750 -2730 1910 -2690
rect 2480 -3060 2660 -3010
rect 1750 -3150 1910 -3110
rect 1750 -3370 1910 -3330
rect 2700 -3380 2760 -3100
rect 2480 -3470 2660 -3420
rect 1750 -3790 1910 -3750
rect 1550 -3880 1710 -3840
rect 2140 -4220 2700 -4160
rect 1550 -4300 1710 -4260
rect 1550 -4540 1710 -4500
rect 2740 -4540 2800 -4260
rect 2140 -4640 2700 -4580
rect 5900 -4780 5960 -2500
rect 6320 -4780 6380 -1430
rect 1550 -4960 1710 -4920
rect 1480 -6070 5080 -6020
rect 174 -6584 1304 -6168
rect 3900 -6586 5030 -6170
rect 30 -7890 80 -6750
rect 5130 -7890 5180 -6120
rect 120 -7980 5080 -7930
<< metal1 >>
rect 1400 4920 1492 5196
rect 1768 4920 1860 5196
rect 2136 4920 2228 5196
rect 2504 4920 2596 5196
rect 2872 4920 2964 5196
rect 3240 4920 3332 5196
rect 3608 4920 3700 5196
rect 3976 4920 4068 5196
rect 4344 4920 4436 5196
rect 4712 4920 4804 5196
rect 5080 4920 5172 5196
rect 5448 4920 5540 5196
rect 5816 4920 5908 5196
rect 6184 4920 6276 5196
rect 6552 4920 6644 5196
rect 6920 4920 7012 5196
rect 1410 4860 1620 4920
rect 420 4750 740 4780
rect 420 4700 540 4750
rect 720 4700 740 4750
rect 420 4690 740 4700
rect 870 4740 1470 4750
rect 870 4690 980 4740
rect 1230 4690 1470 4740
rect 420 4650 530 4690
rect 870 4680 1470 4690
rect 870 4660 950 4680
rect 420 4360 450 4650
rect 500 4570 530 4650
rect 590 4600 880 4660
rect 940 4600 950 4660
rect 1190 4640 1470 4680
rect 710 4590 950 4600
rect 980 4590 1160 4640
rect 500 4450 610 4570
rect 980 4560 1070 4590
rect 1190 4560 1280 4640
rect 650 4460 1070 4560
rect 1160 4460 1280 4560
rect 500 4360 530 4450
rect 710 4420 940 4430
rect 590 4360 850 4420
rect 420 4330 530 4360
rect 840 4350 850 4360
rect 930 4350 940 4420
rect 840 4340 940 4350
rect 970 4420 1070 4460
rect 1170 4450 1280 4460
rect 970 4370 1160 4420
rect 1190 4370 1280 4450
rect 1320 4370 1470 4640
rect 420 4320 740 4330
rect 420 4270 540 4320
rect 720 4270 740 4320
rect 420 4180 740 4270
rect 970 4210 1070 4370
rect 1190 4340 1470 4370
rect 420 4020 440 4180
rect 720 4020 740 4180
rect 420 4000 740 4020
rect 890 3970 1070 4210
rect 1100 4320 1470 4340
rect 1100 4280 1120 4320
rect 1230 4280 1470 4320
rect 1100 4150 1470 4280
rect 1560 4320 1620 4860
rect 1780 4440 1840 4920
rect 2155 4545 2205 4920
rect 2525 4645 2575 4920
rect 2895 4735 2945 4920
rect 3265 4755 3315 4920
rect 2895 4685 3185 4735
rect 3265 4705 3355 4755
rect 2525 4595 2995 4645
rect 2155 4495 2695 4545
rect 1780 4380 2540 4440
rect 1560 4260 2390 4320
rect 1100 4100 1530 4150
rect 890 3950 1100 3970
rect 890 3850 910 3950
rect 1080 3850 1100 3950
rect 890 3830 1100 3850
rect 1160 3800 1530 4100
rect 1160 3600 1180 3800
rect 1470 3600 1530 3800
rect 1160 3490 1530 3600
rect 1220 3130 1530 3490
rect 1710 3780 2040 3800
rect 1710 3620 1730 3780
rect 2020 3620 2040 3780
rect 1560 3460 1660 3470
rect 1560 3350 1570 3460
rect 1650 3350 1660 3460
rect 1560 3340 1660 3350
rect 1220 2880 1470 3130
rect 1520 2880 1530 3130
rect 1570 2950 1620 3340
rect 1710 3220 2040 3620
rect 2090 3460 2190 3470
rect 2090 3350 2100 3460
rect 2180 3350 2190 3460
rect 2090 3340 2190 3350
rect 1710 3170 1720 3220
rect 2030 3170 2040 3220
rect 1710 3120 2040 3170
rect 1650 3060 2070 3120
rect 2100 2950 2150 3340
rect 2330 3250 2390 4260
rect 2480 3250 2540 4380
rect 2645 3250 2695 4495
rect 2945 3250 2995 4595
rect 2324 3190 2330 3250
rect 2390 3190 2396 3250
rect 2474 3190 2480 3250
rect 2540 3190 2546 3250
rect 2630 3246 2710 3250
rect 2630 3194 2644 3246
rect 2696 3194 2710 3246
rect 2630 3190 2710 3194
rect 2930 3246 3010 3250
rect 3135 3246 3185 4685
rect 3305 3246 3355 4705
rect 3635 4645 3685 4920
rect 3465 4595 3685 4645
rect 3465 3246 3515 4595
rect 3995 4545 4045 4920
rect 3625 4495 4045 4545
rect 3625 3246 3675 4495
rect 4375 4435 4425 4920
rect 3765 4385 4425 4435
rect 3765 3246 3815 4385
rect 4735 4315 4785 4920
rect 3915 4265 4785 4315
rect 3915 3246 3965 4265
rect 2930 3194 2944 3246
rect 2996 3194 3010 3246
rect 3128 3194 3134 3246
rect 3186 3194 3192 3246
rect 3298 3194 3304 3246
rect 3356 3194 3362 3246
rect 3458 3194 3464 3246
rect 3516 3194 3522 3246
rect 3618 3194 3624 3246
rect 3676 3194 3682 3246
rect 3758 3194 3764 3246
rect 3816 3194 3822 3246
rect 3908 3194 3914 3246
rect 3966 3194 3972 3246
rect 2930 3190 3010 3194
rect 1650 2890 2070 2950
rect 1220 2850 1530 2880
rect 1220 2830 1790 2850
rect 1220 2810 1570 2830
rect 1220 2700 1240 2810
rect 1350 2700 1570 2810
rect 1220 2690 1570 2700
rect 1770 2690 1790 2830
rect 1220 2680 1790 2690
rect 1610 2580 1710 2640
rect 1770 2580 1780 2640
rect 1850 2540 2060 2890
rect 5095 2845 5145 4920
rect 5465 2966 5515 4920
rect 5830 3520 5890 4920
rect 6200 3660 6260 4920
rect 6570 4200 6630 4920
rect 6940 4200 7000 4920
rect 6570 4140 6888 4200
rect 6940 4140 7026 4200
rect 6200 3600 6480 3660
rect 5830 3460 6340 3520
rect 6280 3250 6340 3460
rect 6420 3250 6480 3600
rect 6274 3190 6280 3250
rect 6340 3190 6346 3250
rect 6414 3190 6420 3250
rect 6480 3190 6486 3250
rect 6828 3248 6888 4140
rect 6966 3248 7026 4140
rect 6822 3188 6828 3248
rect 6888 3188 6894 3248
rect 6960 3188 6966 3248
rect 7026 3188 7032 3248
rect 5458 2914 5464 2966
rect 5516 2914 5522 2966
rect 5095 2795 5680 2845
rect 610 2520 1630 2540
rect 610 1980 630 2520
rect 790 1980 1630 2520
rect 610 1960 1630 1980
rect 1670 1960 2060 2540
rect 4900 2560 5490 2570
rect 4900 2490 4910 2560
rect 5030 2550 5490 2560
rect 5030 2500 5290 2550
rect 5470 2500 5490 2550
rect 5030 2490 5490 2500
rect 4900 2480 5490 2490
rect 5630 2450 5680 2795
rect 5880 2550 6750 2570
rect 5270 2400 5680 2450
rect 5730 2510 5830 2520
rect 5730 2430 5740 2510
rect 5820 2470 5830 2510
rect 5880 2510 5900 2550
rect 6160 2510 6570 2550
rect 5880 2500 6570 2510
rect 5820 2430 6080 2470
rect 5730 2420 6080 2430
rect 4050 2360 5360 2370
rect 4050 2280 4060 2360
rect 4240 2280 5360 2360
rect 4050 2270 5360 2280
rect 5400 2360 5590 2370
rect 5400 2280 5510 2360
rect 5580 2280 5590 2360
rect 5400 2270 5590 2280
rect 5630 2240 5680 2400
rect 5980 2390 6080 2420
rect 6200 2460 6570 2500
rect 5340 2190 5680 2240
rect 4900 2150 5490 2160
rect 4900 2080 4910 2150
rect 5030 2140 5490 2150
rect 5030 2090 5290 2140
rect 5470 2090 5490 2140
rect 5030 2080 5490 2090
rect 4900 2070 5490 2080
rect 1610 1860 1710 1920
rect 1770 1860 1780 1920
rect 1220 1810 1790 1820
rect 1220 1800 1570 1810
rect 1220 1690 1240 1800
rect 1350 1690 1570 1800
rect 1220 1680 1570 1690
rect 1730 1680 1790 1810
rect 1220 1670 1790 1680
rect 1610 1570 1710 1630
rect 1770 1570 1780 1630
rect 1850 1530 2060 1960
rect 4620 2020 6165 2030
rect 4620 1950 4630 2020
rect 4810 1950 6165 2020
rect 4620 1940 6165 1950
rect 4900 1890 5490 1900
rect 4900 1820 4910 1890
rect 5030 1880 5490 1890
rect 5030 1830 5300 1880
rect 5460 1830 5490 1880
rect 5030 1820 5490 1830
rect 4900 1810 5490 1820
rect 5629 1876 5681 1882
rect 5629 1818 5681 1824
rect 5630 1780 5680 1818
rect 5280 1730 5680 1780
rect 4330 1630 5360 1700
rect 4330 1550 4350 1630
rect 4510 1600 5360 1630
rect 5400 1690 5590 1700
rect 5400 1610 5510 1690
rect 5580 1610 5590 1690
rect 5400 1600 5590 1610
rect 4510 1550 4600 1600
rect 5630 1570 5680 1730
rect 4330 1530 4600 1550
rect 290 1510 1630 1530
rect 290 970 310 1510
rect 470 970 1630 1510
rect 290 950 1630 970
rect 1670 950 2060 1530
rect 5340 1520 5680 1570
rect 5780 1560 5860 1570
rect 5780 1510 5800 1560
rect 5840 1550 5860 1560
rect 5980 1550 6080 1590
rect 6200 1550 6210 2460
rect 5840 1510 6210 1550
rect 6260 1510 6570 2460
rect 4900 1480 5490 1490
rect 4900 1410 4910 1480
rect 5030 1470 5490 1480
rect 5030 1420 5300 1470
rect 5460 1420 5490 1470
rect 5030 1410 5490 1420
rect 4900 1400 5490 1410
rect 5780 1460 6570 1510
rect 5780 1420 5900 1460
rect 6160 1420 6570 1460
rect 6730 1420 6750 2550
rect 5780 1400 6750 1420
rect 4900 1030 5520 1040
rect 4900 970 4910 1030
rect 5030 1020 5520 1030
rect 5030 970 5340 1020
rect 5500 970 5520 1020
rect 6140 1030 6750 1050
rect 4900 960 5520 970
rect 5990 980 6110 990
rect 5620 930 5700 940
rect 5620 920 5630 930
rect 1220 870 1370 890
rect 1220 760 1240 870
rect 1350 810 1370 870
rect 1610 850 1710 910
rect 1770 850 1780 910
rect 5390 870 5630 920
rect 5690 870 5700 930
rect 5990 900 6000 980
rect 6080 940 6110 980
rect 6140 980 6160 1030
rect 6280 980 6570 1030
rect 6140 970 6570 980
rect 6080 900 6190 940
rect 5990 890 6190 900
rect 5620 860 5700 870
rect 6090 860 6190 890
rect 6310 920 6570 970
rect 4050 830 4250 850
rect 1350 800 1790 810
rect 1350 760 1570 800
rect 1220 750 1570 760
rect 1730 750 1790 800
rect 1220 740 1790 750
rect 4050 750 4070 830
rect 4220 750 5400 830
rect 5440 820 5980 830
rect 5440 760 5890 820
rect 5970 760 5980 820
rect 5440 750 5980 760
rect 4050 730 4250 750
rect 5620 710 5700 720
rect 5390 660 5630 710
rect 5620 650 5630 660
rect 5690 650 5700 710
rect 5620 640 5700 650
rect 4900 610 5520 620
rect 1220 580 2830 590
rect 1220 510 1230 580
rect 1300 570 2830 580
rect 1300 520 1570 570
rect 1300 510 1310 520
rect 1220 500 1310 510
rect 1550 510 1570 520
rect 1740 560 2830 570
rect 1740 510 2650 560
rect 1550 500 2650 510
rect 2630 490 2650 500
rect 2810 490 2830 560
rect 4900 550 4910 610
rect 5030 560 5340 610
rect 5500 560 5520 610
rect 5030 550 5520 560
rect 4900 540 5520 550
rect 1350 480 1430 490
rect 1350 420 1360 480
rect 1420 460 1430 480
rect 2630 470 2830 490
rect 2273 460 2279 461
rect 1420 420 2279 460
rect 1350 410 2279 420
rect 2273 409 2279 410
rect 2331 409 2337 461
rect 4620 440 6280 450
rect 610 360 1620 380
rect 610 10 630 360
rect 790 10 1620 360
rect 610 -10 1620 10
rect 1670 360 1870 370
rect 1670 0 1780 360
rect 1860 0 1870 360
rect 4620 350 4630 440
rect 4810 350 6280 440
rect 4620 340 6280 350
rect 4900 230 5520 240
rect 4900 170 4910 230
rect 5030 220 5520 230
rect 5030 170 5340 220
rect 5500 170 5520 220
rect 4900 160 5520 170
rect 5620 130 5700 140
rect 5620 120 5630 130
rect 5390 70 5630 120
rect 5690 70 5700 130
rect 5620 60 5700 70
rect 4330 30 4530 50
rect 1670 -10 1870 0
rect 2200 10 2830 30
rect 2200 0 2650 10
rect 2200 -50 2220 0
rect 2460 -50 2650 0
rect 1350 -60 1680 -50
rect 2200 -60 2650 -50
rect 1350 -120 1360 -60
rect 1420 -100 1680 -60
rect 2480 -90 2650 -60
rect 1420 -120 1430 -100
rect 1350 -130 1430 -120
rect 1220 -140 1300 -130
rect 1220 -200 1230 -140
rect 1290 -170 1300 -140
rect 1910 -150 2380 -100
rect 1550 -160 1760 -150
rect 1550 -170 1570 -160
rect 1290 -200 1570 -170
rect 1740 -200 1760 -160
rect 1220 -210 1760 -200
rect 890 -250 1090 -230
rect 1910 -250 1960 -150
rect 2480 -180 2500 -90
rect 890 -340 910 -250
rect 1070 -340 1960 -250
rect 890 -360 1090 -340
rect 1220 -390 1760 -380
rect 1220 -450 1230 -390
rect 1290 -420 1570 -390
rect 1290 -450 1300 -420
rect 1550 -430 1570 -420
rect 1740 -430 1760 -390
rect 1550 -440 1760 -430
rect 1910 -430 1960 -340
rect 2000 -200 2280 -190
rect 2000 -380 2010 -200
rect 2140 -380 2280 -200
rect 2000 -390 2280 -380
rect 2390 -400 2500 -180
rect 1220 -460 1300 -450
rect 1350 -470 1430 -460
rect 1350 -530 1360 -470
rect 1420 -490 1430 -470
rect 1910 -480 2380 -430
rect 2480 -490 2500 -400
rect 2560 -490 2650 -90
rect 1420 -530 1680 -490
rect 2480 -520 2650 -490
rect 1350 -540 1680 -530
rect 2200 -530 2650 -520
rect 290 -590 1620 -570
rect 2200 -580 2220 -530
rect 2460 -580 2650 -530
rect 290 -940 310 -590
rect 470 -940 1620 -590
rect 290 -960 1620 -940
rect 1670 -590 1870 -580
rect 1670 -950 1780 -590
rect 1860 -950 1870 -590
rect 2200 -590 2650 -580
rect 2810 -590 2830 10
rect 4330 -50 4350 30
rect 4510 -50 5400 30
rect 5440 20 5980 30
rect 5440 -40 5890 20
rect 5970 -40 5980 20
rect 5440 -50 5980 -40
rect 4330 -70 4530 -50
rect 5620 -90 5700 -80
rect 5390 -140 5630 -90
rect 5620 -150 5630 -140
rect 5690 -150 5700 -90
rect 5620 -160 5700 -150
rect 5890 -140 5980 -110
rect 4900 -190 5520 -180
rect 4900 -250 4910 -190
rect 5030 -240 5340 -190
rect 5500 -240 5520 -190
rect 5030 -250 5520 -240
rect 4900 -260 5520 -250
rect 2200 -610 2830 -590
rect 5890 -810 5910 -140
rect 5960 -780 5980 -140
rect 6090 -780 6190 -750
rect 6310 -780 6320 920
rect 5960 -810 6320 -780
rect 6380 -810 6570 920
rect 5890 -860 6570 -810
rect 5890 -910 6010 -860
rect 6270 -910 6570 -860
rect 6730 -910 6750 1030
rect 5890 -930 6750 -910
rect 1670 -960 1870 -950
rect 2273 -1000 2279 -999
rect 1350 -1010 2279 -1000
rect 1350 -1070 1360 -1010
rect 1420 -1050 2279 -1010
rect 1420 -1070 1430 -1050
rect 2273 -1051 2279 -1050
rect 2331 -1051 2337 -999
rect 1350 -1080 1430 -1070
rect 2630 -1080 2830 -1060
rect 2630 -1090 2650 -1080
rect 1220 -1100 1310 -1090
rect 1220 -1170 1230 -1100
rect 1300 -1110 1310 -1100
rect 1550 -1100 2650 -1090
rect 1550 -1110 1570 -1100
rect 1300 -1160 1570 -1110
rect 1740 -1160 2650 -1100
rect 1300 -1170 2650 -1160
rect 1220 -1180 2650 -1170
rect 1460 -1280 2650 -1180
rect 1460 -1330 1480 -1280
rect 1650 -1320 2650 -1280
rect 2810 -1320 2830 -1080
rect 1650 -1330 2830 -1320
rect 1460 -1340 2830 -1330
rect 4900 -1330 5520 -1320
rect 1350 -1360 1430 -1350
rect 1350 -1420 1360 -1360
rect 1420 -1380 1430 -1360
rect 2273 -1380 2279 -1379
rect 1420 -1420 2279 -1380
rect 1350 -1430 2279 -1420
rect 2273 -1431 2279 -1430
rect 2331 -1431 2337 -1379
rect 4900 -1390 4910 -1330
rect 5030 -1340 5520 -1330
rect 5030 -1390 5340 -1340
rect 5500 -1390 5520 -1340
rect 6010 -1340 6750 -1320
rect 4900 -1400 5520 -1390
rect 5880 -1380 5980 -1370
rect 5620 -1430 5700 -1420
rect 5620 -1440 5630 -1430
rect 610 -1480 1540 -1460
rect 610 -1640 630 -1480
rect 790 -1640 1540 -1480
rect 610 -1660 1540 -1640
rect 1580 -1470 1770 -1460
rect 1580 -1650 1690 -1470
rect 1760 -1650 1770 -1470
rect 5390 -1490 5630 -1440
rect 5690 -1490 5700 -1430
rect 5880 -1440 5890 -1380
rect 5970 -1420 5980 -1380
rect 6010 -1380 6030 -1340
rect 6270 -1380 6570 -1340
rect 6010 -1390 6570 -1380
rect 5970 -1440 6190 -1420
rect 5880 -1480 6190 -1440
rect 6310 -1430 6570 -1390
rect 5620 -1500 5700 -1490
rect 4050 -1530 4250 -1510
rect 2030 -1570 3030 -1560
rect 2030 -1620 2050 -1570
rect 2660 -1580 3030 -1570
rect 2660 -1620 2850 -1580
rect 2030 -1630 2850 -1620
rect 1580 -1660 1770 -1650
rect 2680 -1650 2850 -1630
rect 1350 -1700 1600 -1690
rect 1350 -1760 1360 -1700
rect 1420 -1740 1600 -1700
rect 1800 -1720 2570 -1670
rect 1420 -1760 1430 -1740
rect 1350 -1770 1430 -1760
rect 1220 -1780 1310 -1770
rect 1220 -1850 1230 -1780
rect 1300 -1800 1310 -1780
rect 1460 -1800 1670 -1790
rect 1300 -1850 1480 -1800
rect 1650 -1850 1670 -1800
rect 1220 -1860 1670 -1850
rect 890 -1870 1090 -1860
rect 890 -2020 910 -1870
rect 1070 -1890 1090 -1870
rect 1800 -1890 1850 -1720
rect 2680 -1750 2690 -1650
rect 1070 -2010 1850 -1890
rect 1070 -2020 1090 -2010
rect 890 -2040 1090 -2020
rect 1220 -2060 1670 -2040
rect 1220 -2130 1230 -2060
rect 1300 -2100 1480 -2060
rect 1300 -2130 1310 -2100
rect 1460 -2110 1480 -2100
rect 1650 -2110 1670 -2060
rect 1460 -2120 1670 -2110
rect 1220 -2140 1310 -2130
rect 1350 -2140 1430 -2130
rect 1350 -2200 1360 -2140
rect 1420 -2160 1430 -2140
rect 1800 -2160 1850 -2010
rect 1890 -1770 2110 -1760
rect 1890 -2110 1900 -1770
rect 1990 -2110 2110 -1770
rect 1890 -2120 2110 -2110
rect 2580 -2130 2690 -1750
rect 1420 -2200 1600 -2160
rect 1350 -2210 1600 -2200
rect 1800 -2210 2570 -2160
rect 2680 -2230 2690 -2130
rect 2750 -2230 2850 -1650
rect 290 -2260 1540 -2240
rect 290 -2420 310 -2260
rect 470 -2420 1540 -2260
rect 290 -2440 1540 -2420
rect 1580 -2250 1770 -2240
rect 2680 -2250 2850 -2230
rect 1580 -2430 1690 -2250
rect 1760 -2430 1770 -2250
rect 2030 -2260 2850 -2250
rect 2030 -2310 2050 -2260
rect 2660 -2300 2850 -2260
rect 3010 -2300 3030 -1580
rect 4050 -1610 4070 -1530
rect 4220 -1610 5400 -1530
rect 5440 -1540 5980 -1530
rect 5440 -1600 5890 -1540
rect 5970 -1600 5980 -1540
rect 5440 -1610 5980 -1600
rect 4050 -1630 4250 -1610
rect 5620 -1650 5700 -1640
rect 5390 -1700 5630 -1650
rect 5620 -1710 5630 -1700
rect 5690 -1710 5700 -1650
rect 5620 -1720 5700 -1710
rect 4900 -1750 5520 -1740
rect 4900 -1810 4910 -1750
rect 5030 -1800 5340 -1750
rect 5500 -1800 5520 -1750
rect 5030 -1810 5520 -1800
rect 4900 -1820 5520 -1810
rect 4620 -1920 6280 -1910
rect 4620 -2020 4630 -1920
rect 4810 -2020 6280 -1920
rect 4620 -2030 6280 -2020
rect 4900 -2130 5520 -2120
rect 4900 -2190 4910 -2130
rect 5030 -2140 5520 -2130
rect 5030 -2190 5340 -2140
rect 5500 -2190 5520 -2140
rect 4900 -2200 5520 -2190
rect 5620 -2230 5700 -2220
rect 5620 -2240 5630 -2230
rect 5390 -2290 5630 -2240
rect 5690 -2290 5700 -2230
rect 5620 -2300 5700 -2290
rect 2660 -2310 3030 -2300
rect 2030 -2320 3030 -2310
rect 4330 -2330 4530 -2310
rect 4330 -2410 4350 -2330
rect 4510 -2410 5400 -2330
rect 5440 -2340 5980 -2330
rect 5440 -2400 5890 -2340
rect 5970 -2400 5980 -2340
rect 5440 -2410 5980 -2400
rect 4330 -2430 4530 -2410
rect 1580 -2440 1770 -2430
rect 5620 -2450 5700 -2440
rect 2273 -2470 2279 -2469
rect 1350 -2480 2279 -2470
rect 1350 -2540 1360 -2480
rect 1420 -2520 2279 -2480
rect 1420 -2540 1430 -2520
rect 2273 -2521 2279 -2520
rect 2331 -2521 2337 -2469
rect 5390 -2500 5630 -2450
rect 5620 -2510 5630 -2500
rect 5690 -2510 5700 -2450
rect 5620 -2520 5700 -2510
rect 5890 -2500 5970 -2480
rect 1220 -2550 1310 -2540
rect 1350 -2550 1430 -2540
rect 4900 -2550 5520 -2540
rect 1220 -2710 1230 -2550
rect 1300 -2580 1310 -2550
rect 1460 -2570 3030 -2560
rect 1460 -2580 1480 -2570
rect 1300 -2620 1480 -2580
rect 1650 -2580 3030 -2570
rect 1650 -2620 2850 -2580
rect 1300 -2690 2850 -2620
rect 1300 -2710 1750 -2690
rect 1220 -2720 1750 -2710
rect 1730 -2730 1750 -2720
rect 1910 -2700 2850 -2690
rect 3010 -2700 3030 -2580
rect 4900 -2610 4910 -2550
rect 5030 -2600 5340 -2550
rect 5500 -2600 5520 -2550
rect 5030 -2610 5520 -2600
rect 4900 -2620 5520 -2610
rect 1910 -2720 3030 -2700
rect 1910 -2730 1930 -2720
rect 1730 -2750 1930 -2730
rect 1600 -2830 1610 -2770
rect 1680 -2790 1690 -2770
rect 2303 -2790 2309 -2789
rect 1680 -2830 2309 -2790
rect 610 -2850 810 -2830
rect 1600 -2840 2309 -2830
rect 2303 -2841 2309 -2840
rect 2361 -2841 2367 -2789
rect 610 -2990 630 -2850
rect 790 -2870 810 -2850
rect 790 -2970 1810 -2870
rect 1860 -2880 2060 -2870
rect 1860 -2960 1970 -2880
rect 2050 -2960 2060 -2880
rect 1860 -2970 2060 -2960
rect 790 -2990 810 -2970
rect 610 -3010 810 -2990
rect 1600 -3010 1880 -3000
rect 1600 -3070 1610 -3010
rect 1680 -3050 1880 -3010
rect 2460 -3010 3030 -3000
rect 1680 -3070 1690 -3050
rect 2460 -3060 2480 -3010
rect 2660 -3020 3030 -3010
rect 2660 -3060 2850 -3020
rect 2460 -3070 2850 -3060
rect 1220 -3090 1310 -3080
rect 1220 -3160 1230 -3090
rect 1300 -3100 1310 -3090
rect 1730 -3100 1940 -3090
rect 1300 -3110 1940 -3100
rect 1300 -3150 1750 -3110
rect 1910 -3150 1940 -3110
rect 1300 -3160 1940 -3150
rect 1220 -3170 1940 -3160
rect 2060 -3110 2430 -3080
rect 2620 -3100 2850 -3070
rect 2060 -3120 2580 -3110
rect 890 -3190 1090 -3170
rect 890 -3290 910 -3190
rect 1070 -3200 1090 -3190
rect 2060 -3200 2100 -3120
rect 1070 -3280 2100 -3200
rect 1070 -3290 1090 -3280
rect 890 -3310 1090 -3290
rect 1220 -3320 1940 -3310
rect 1220 -3390 1230 -3320
rect 1300 -3330 1940 -3320
rect 1300 -3370 1750 -3330
rect 1910 -3370 1940 -3330
rect 1300 -3380 1940 -3370
rect 1300 -3390 1310 -3380
rect 1730 -3390 1940 -3380
rect 2060 -3360 2100 -3280
rect 2130 -3160 2360 -3150
rect 2390 -3160 2580 -3120
rect 2130 -3320 2140 -3160
rect 2270 -3180 2360 -3160
rect 2620 -3180 2700 -3100
rect 2270 -3200 2370 -3180
rect 2600 -3200 2700 -3180
rect 2270 -3280 2380 -3200
rect 2590 -3280 2700 -3200
rect 2270 -3300 2370 -3280
rect 2600 -3300 2700 -3280
rect 2270 -3320 2360 -3300
rect 2130 -3330 2360 -3320
rect 2390 -3360 2580 -3320
rect 2060 -3370 2580 -3360
rect 1220 -3400 1310 -3390
rect 2060 -3400 2430 -3370
rect 2620 -3380 2700 -3300
rect 2760 -3380 2850 -3100
rect 2620 -3410 2850 -3380
rect 1600 -3470 1610 -3410
rect 1680 -3430 1690 -3410
rect 2460 -3420 2850 -3410
rect 1680 -3470 1880 -3430
rect 1600 -3480 1880 -3470
rect 2460 -3470 2480 -3420
rect 2660 -3460 2850 -3420
rect 3010 -3460 3030 -3020
rect 2660 -3470 3030 -3460
rect 2460 -3480 3030 -3470
rect 290 -3510 490 -3490
rect 290 -3610 310 -3510
rect 470 -3610 1810 -3510
rect 1860 -3520 2060 -3510
rect 1860 -3600 1970 -3520
rect 2050 -3600 2060 -3520
rect 1860 -3610 2060 -3600
rect 290 -3630 490 -3610
rect 2298 -3640 2304 -3639
rect 1600 -3650 2304 -3640
rect 1600 -3710 1610 -3650
rect 1680 -3690 2304 -3650
rect 1680 -3710 1690 -3690
rect 2298 -3691 2304 -3690
rect 2356 -3691 2362 -3639
rect 1220 -3730 1310 -3720
rect 1220 -3880 1230 -3730
rect 1300 -3740 1310 -3730
rect 1730 -3740 1940 -3730
rect 1300 -3750 3030 -3740
rect 1300 -3790 1750 -3750
rect 1910 -3760 3030 -3750
rect 1910 -3790 2850 -3760
rect 1300 -3840 2850 -3790
rect 1300 -3870 1550 -3840
rect 1220 -3890 1300 -3880
rect 1530 -3880 1550 -3870
rect 1710 -3880 2850 -3840
rect 3010 -3880 3030 -3760
rect 1530 -3900 3030 -3880
rect 1420 -3920 1500 -3910
rect 1420 -3980 1430 -3920
rect 1490 -3940 1500 -3920
rect 2303 -3940 2309 -3939
rect 1490 -3980 2309 -3940
rect 1420 -3990 2309 -3980
rect 2303 -3991 2309 -3990
rect 2361 -3991 2367 -3939
rect 610 -4020 810 -4000
rect 610 -4120 630 -4020
rect 790 -4120 1610 -4020
rect 1650 -4030 1870 -4020
rect 1650 -4110 1790 -4030
rect 1650 -4120 1870 -4110
rect 610 -4140 810 -4120
rect 1420 -4160 1670 -4150
rect 1420 -4220 1430 -4160
rect 1490 -4200 1670 -4160
rect 2120 -4160 3030 -4150
rect 1490 -4220 1500 -4200
rect 1420 -4230 1500 -4220
rect 2120 -4220 2140 -4160
rect 2700 -4170 3030 -4160
rect 2700 -4220 2850 -4170
rect 2120 -4230 2850 -4220
rect 1220 -4250 1300 -4240
rect 1220 -4320 1230 -4250
rect 1530 -4260 1740 -4240
rect 1530 -4270 1550 -4260
rect 1300 -4300 1550 -4270
rect 1710 -4300 1740 -4260
rect 2730 -4260 2850 -4230
rect 1300 -4320 1740 -4300
rect 1860 -4320 2620 -4270
rect 890 -4350 1090 -4330
rect 1860 -4350 1900 -4320
rect 2730 -4350 2740 -4260
rect 890 -4450 910 -4350
rect 1070 -4450 1900 -4350
rect 1930 -4360 2210 -4350
rect 1930 -4440 1940 -4360
rect 2020 -4440 2210 -4360
rect 1930 -4450 2210 -4440
rect 2630 -4450 2740 -4350
rect 890 -4470 1090 -4450
rect 1860 -4480 1900 -4450
rect 1220 -4550 1230 -4480
rect 1300 -4500 1740 -4480
rect 1300 -4540 1550 -4500
rect 1710 -4540 1740 -4500
rect 1860 -4530 2620 -4480
rect 1220 -4560 1300 -4550
rect 1530 -4560 1740 -4540
rect 2730 -4540 2740 -4450
rect 2800 -4540 2850 -4260
rect 2730 -4570 2850 -4540
rect 1420 -4580 1500 -4570
rect 1420 -4640 1430 -4580
rect 1490 -4600 1500 -4580
rect 2120 -4580 2850 -4570
rect 1490 -4640 1670 -4600
rect 1420 -4650 1670 -4640
rect 2120 -4640 2140 -4580
rect 2700 -4630 2850 -4580
rect 3010 -4630 3030 -4170
rect 2700 -4640 3030 -4630
rect 2120 -4650 3030 -4640
rect 290 -4680 490 -4660
rect 290 -4780 310 -4680
rect 470 -4780 1610 -4680
rect 1650 -4690 1870 -4680
rect 1650 -4770 1790 -4690
rect 1650 -4780 1870 -4770
rect 5890 -4780 5900 -2500
rect 5960 -4740 5970 -2500
rect 6090 -4740 6190 -4710
rect 6310 -4740 6320 -1430
rect 5960 -4780 6320 -4740
rect 6380 -4780 6570 -1430
rect 290 -4800 490 -4780
rect 2303 -4810 2309 -4809
rect 1420 -4820 2309 -4810
rect 1420 -4880 1430 -4820
rect 1490 -4860 2309 -4820
rect 1490 -4880 1500 -4860
rect 2303 -4861 2309 -4860
rect 2361 -4861 2367 -4809
rect 1420 -4890 1500 -4880
rect 5890 -4870 6570 -4780
rect 6730 -4870 6750 -1340
rect 5890 -4890 6750 -4870
rect 1220 -4910 1300 -4900
rect 1220 -4980 1230 -4910
rect 1530 -4920 3030 -4900
rect 1530 -4930 1550 -4920
rect 1300 -4960 1550 -4930
rect 1710 -4960 2850 -4920
rect 1300 -4980 2850 -4960
rect 2830 -5040 2850 -4980
rect 3010 -5040 3030 -4920
rect 2830 -5060 3030 -5040
rect 5080 -5900 5300 -5890
rect 5080 -5990 5090 -5900
rect 1460 -6020 5090 -5990
rect 1460 -6070 1480 -6020
rect 5080 -6070 5090 -6020
rect 1460 -6100 5090 -6070
rect 5290 -6100 5300 -5900
rect 1460 -6110 5300 -6100
rect 1460 -6120 5210 -6110
rect 150 -6150 1330 -6140
rect 150 -6600 160 -6150
rect 1320 -6600 1330 -6150
rect 150 -6610 1330 -6600
rect 3880 -6160 5050 -6150
rect 3880 -6600 3890 -6160
rect 5040 -6600 5050 -6160
rect 3880 -6610 5050 -6600
rect 0 -6750 130 -6730
rect 0 -7890 30 -6750
rect 80 -7880 130 -6750
rect 5080 -7880 5130 -6120
rect 80 -7890 5130 -7880
rect 5180 -7890 5210 -6120
rect 0 -7930 5210 -7890
rect 0 -7980 120 -7930
rect 5080 -7980 5210 -7930
rect 0 -8010 5210 -7980
<< via1 >>
rect 880 4650 940 4660
rect 880 4600 930 4650
rect 930 4600 940 4650
rect 850 4410 930 4420
rect 850 4370 880 4410
rect 880 4370 930 4410
rect 850 4350 930 4370
rect 440 4020 720 4180
rect 910 3850 1080 3950
rect 1180 3600 1470 3800
rect 1730 3620 2020 3780
rect 1570 3350 1650 3460
rect 2100 3350 2180 3460
rect 2330 3190 2390 3250
rect 2480 3190 2540 3250
rect 2644 3194 2696 3246
rect 2944 3194 2996 3246
rect 3134 3194 3186 3246
rect 3304 3194 3356 3246
rect 3464 3194 3516 3246
rect 3624 3194 3676 3246
rect 3764 3194 3816 3246
rect 3914 3194 3966 3246
rect 1240 2700 1350 2810
rect 1710 2580 1770 2640
rect 6280 3190 6340 3250
rect 6420 3190 6480 3250
rect 6828 3188 6888 3248
rect 6966 3188 7026 3248
rect 5464 2914 5516 2966
rect 630 1980 790 2520
rect 4910 2490 5030 2560
rect 5740 2430 5820 2510
rect 4060 2280 4240 2360
rect 5510 2280 5580 2360
rect 4910 2080 5030 2150
rect 1710 1860 1770 1920
rect 1240 1690 1350 1800
rect 1710 1570 1770 1630
rect 4630 1950 4810 2020
rect 4910 1820 5030 1890
rect 5629 1824 5681 1876
rect 4350 1550 4510 1630
rect 5510 1610 5580 1690
rect 310 970 470 1510
rect 4910 1410 5030 1480
rect 6570 1420 6730 2550
rect 4910 970 5030 1030
rect 1240 760 1350 870
rect 1710 850 1770 910
rect 5630 870 5690 930
rect 6000 900 6080 980
rect 4070 750 4220 830
rect 5890 760 5970 820
rect 5630 650 5690 710
rect 1230 510 1300 580
rect 2650 490 2810 560
rect 4910 550 5030 610
rect 1360 420 1420 480
rect 2279 409 2331 461
rect 630 10 790 360
rect 1780 0 1860 360
rect 4630 350 4810 440
rect 4910 170 5030 230
rect 5630 70 5690 130
rect 1360 -120 1420 -60
rect 1230 -200 1290 -140
rect 910 -340 1070 -250
rect 1230 -450 1290 -390
rect 2010 -380 2140 -200
rect 1360 -530 1420 -470
rect 310 -940 470 -590
rect 1780 -950 1860 -590
rect 2650 -590 2810 10
rect 4350 -50 4510 30
rect 5890 -40 5970 20
rect 5630 -150 5690 -90
rect 4910 -250 5030 -190
rect 6570 -910 6730 1030
rect 1360 -1070 1420 -1010
rect 2279 -1051 2331 -999
rect 1230 -1170 1300 -1100
rect 2650 -1320 2810 -1080
rect 1360 -1420 1420 -1360
rect 2279 -1431 2331 -1379
rect 4910 -1390 5030 -1330
rect 630 -1640 790 -1480
rect 1690 -1650 1760 -1470
rect 5630 -1490 5690 -1430
rect 5890 -1440 5970 -1380
rect 1360 -1760 1420 -1700
rect 1230 -1850 1300 -1780
rect 910 -2020 1070 -1870
rect 1230 -2130 1300 -2060
rect 1360 -2200 1420 -2140
rect 1900 -2110 1990 -1770
rect 310 -2420 470 -2260
rect 1690 -2430 1760 -2250
rect 2850 -2300 3010 -1580
rect 4070 -1610 4220 -1530
rect 5890 -1600 5970 -1540
rect 5630 -1710 5690 -1650
rect 4910 -1810 5030 -1750
rect 4630 -2020 4810 -1920
rect 4910 -2190 5030 -2130
rect 5630 -2290 5690 -2230
rect 4350 -2410 4510 -2330
rect 5890 -2400 5970 -2340
rect 1360 -2540 1420 -2480
rect 2279 -2521 2331 -2469
rect 5630 -2510 5690 -2450
rect 1230 -2710 1300 -2550
rect 2850 -2700 3010 -2580
rect 4910 -2610 5030 -2550
rect 1610 -2830 1680 -2770
rect 2309 -2841 2361 -2789
rect 630 -2990 790 -2850
rect 1970 -2960 2050 -2880
rect 1610 -3070 1680 -3010
rect 1230 -3160 1300 -3090
rect 910 -3290 1070 -3190
rect 1230 -3390 1300 -3320
rect 2140 -3320 2270 -3160
rect 1610 -3470 1680 -3410
rect 2850 -3460 3010 -3020
rect 310 -3610 470 -3510
rect 1970 -3600 2050 -3520
rect 1610 -3710 1680 -3650
rect 2304 -3691 2356 -3639
rect 1230 -3880 1300 -3730
rect 2850 -3880 3010 -3760
rect 1430 -3980 1490 -3920
rect 2309 -3991 2361 -3939
rect 630 -4120 790 -4020
rect 1790 -4110 1870 -4030
rect 1430 -4220 1490 -4160
rect 1230 -4320 1300 -4250
rect 910 -4450 1070 -4350
rect 1940 -4440 2020 -4360
rect 1230 -4550 1300 -4480
rect 1430 -4640 1490 -4580
rect 2850 -4630 3010 -4170
rect 310 -4780 470 -4680
rect 1790 -4770 1870 -4690
rect 1430 -4880 1490 -4820
rect 2309 -4861 2361 -4809
rect 6570 -4870 6730 -1340
rect 1230 -4980 1300 -4910
rect 2850 -5040 3010 -4920
rect 5090 -6100 5290 -5900
rect 160 -6168 1320 -6150
rect 160 -6584 174 -6168
rect 174 -6584 1304 -6168
rect 1304 -6584 1320 -6168
rect 160 -6600 1320 -6584
rect 3890 -6170 5040 -6160
rect 3890 -6586 3900 -6170
rect 3900 -6586 5030 -6170
rect 5030 -6586 5040 -6170
rect 3890 -6600 5040 -6586
<< metal2 >>
rect 870 4660 950 4670
rect 870 4600 880 4660
rect 940 4600 950 4660
rect 870 4440 950 4600
rect 840 4420 950 4440
rect 840 4350 850 4420
rect 930 4350 950 4420
rect 840 4340 950 4350
rect 420 4180 740 4200
rect 420 4020 440 4180
rect 720 4020 740 4180
rect 420 4000 740 4020
rect 890 3950 1100 3970
rect 890 3850 910 3950
rect 1080 3850 1100 3950
rect 890 3470 1100 3850
rect 1160 3800 1490 3820
rect 1160 3600 1180 3800
rect 1470 3600 1490 3800
rect 1710 3780 2040 3800
rect 1710 3620 1730 3780
rect 2020 3620 2040 3780
rect 1710 3600 2040 3620
rect 1160 3580 1490 3600
rect 890 3460 4820 3470
rect 890 3350 1570 3460
rect 1650 3350 2100 3460
rect 2180 3350 4820 3460
rect 890 3340 4820 3350
rect 610 2520 810 2540
rect 610 1980 630 2520
rect 790 1980 810 2520
rect 610 1960 810 1980
rect 290 1510 490 1530
rect 290 970 310 1510
rect 470 970 490 1510
rect 290 950 490 970
rect 610 360 810 380
rect 610 10 630 360
rect 790 10 810 360
rect 610 -10 810 10
rect 890 -250 1090 3340
rect 2330 3250 2390 3256
rect 1220 2810 1370 2830
rect 1220 2700 1240 2810
rect 1350 2700 1370 2810
rect 1220 1800 1370 2700
rect 2330 2640 2390 3190
rect 1700 2580 1710 2640
rect 1770 2580 2390 2640
rect 2480 3250 2540 3256
rect 2120 1920 2180 2580
rect 2480 2490 2540 3190
rect 2644 3246 2696 3252
rect 2644 3188 2696 3194
rect 2944 3246 2996 3252
rect 2944 3188 2996 3194
rect 3134 3246 3186 3252
rect 3134 3188 3186 3194
rect 3304 3246 3356 3252
rect 3304 3188 3356 3194
rect 3464 3246 3516 3252
rect 3464 3188 3516 3194
rect 3624 3246 3676 3252
rect 3624 3188 3676 3194
rect 3764 3246 3816 3252
rect 3764 3188 3816 3194
rect 3914 3246 3966 3252
rect 3914 3188 3966 3194
rect 1700 1860 1710 1920
rect 1770 1860 2180 1920
rect 2260 2430 2540 2490
rect 1220 1690 1240 1800
rect 1350 1690 1370 1800
rect 1220 870 1370 1690
rect 2260 1630 2320 2430
rect 2645 2275 2695 3188
rect 1700 1570 1710 1630
rect 1770 1570 2320 1630
rect 2455 2225 2695 2275
rect 2120 910 2180 1570
rect 1220 760 1240 870
rect 1350 760 1370 870
rect 1700 850 1710 910
rect 1770 850 2180 910
rect 1220 740 1370 760
rect 890 -340 910 -250
rect 1070 -340 1090 -250
rect 290 -590 490 -570
rect 290 -940 310 -590
rect 470 -940 490 -590
rect 290 -960 490 -940
rect 610 -1480 810 -1460
rect 610 -1640 630 -1480
rect 790 -1640 810 -1480
rect 610 -1660 810 -1640
rect 890 -1870 1090 -340
rect 890 -2020 910 -1870
rect 1070 -2020 1090 -1870
rect 290 -2260 490 -2240
rect 290 -2420 310 -2260
rect 470 -2420 490 -2260
rect 290 -2440 490 -2420
rect 610 -2850 810 -2830
rect 610 -2990 630 -2850
rect 790 -2990 810 -2850
rect 610 -3010 810 -2990
rect 890 -3190 1090 -2020
rect 890 -3290 910 -3190
rect 1070 -3290 1090 -3190
rect 290 -3510 490 -3490
rect 290 -3610 310 -3510
rect 470 -3610 490 -3510
rect 290 -3630 490 -3610
rect 610 -4020 810 -4000
rect 610 -4120 630 -4020
rect 790 -4120 810 -4020
rect 610 -4140 810 -4120
rect 890 -4350 1090 -3290
rect 890 -4450 910 -4350
rect 1070 -4450 1090 -4350
rect 290 -4680 490 -4660
rect 290 -4780 310 -4680
rect 470 -4780 490 -4680
rect 290 -4800 490 -4780
rect 890 -5150 1090 -4450
rect 1220 580 1300 590
rect 1220 510 1230 580
rect 1220 -140 1300 510
rect 1350 480 1430 490
rect 1350 420 1360 480
rect 1420 420 1430 480
rect 1350 -60 1430 420
rect 2279 461 2331 467
rect 2455 460 2505 2225
rect 2630 560 2830 580
rect 2630 490 2650 560
rect 2810 490 2830 560
rect 2630 470 2830 490
rect 2331 410 2505 460
rect 2279 403 2331 409
rect 1770 360 2150 370
rect 1770 0 1780 360
rect 1860 0 2150 360
rect 1770 -10 2150 0
rect 1350 -120 1360 -60
rect 1420 -120 1430 -60
rect 1350 -130 1430 -120
rect 1220 -200 1230 -140
rect 1290 -200 1300 -140
rect 1220 -390 1300 -200
rect 1220 -450 1230 -390
rect 1290 -450 1300 -390
rect 1220 -1100 1300 -450
rect 2000 -200 2150 -10
rect 2000 -380 2010 -200
rect 2140 -380 2150 -200
rect 1350 -470 1430 -460
rect 1350 -530 1360 -470
rect 1420 -530 1430 -470
rect 1350 -1010 1430 -530
rect 2000 -580 2150 -380
rect 1770 -590 2150 -580
rect 1770 -950 1780 -590
rect 1860 -950 2150 -590
rect 2630 10 2830 30
rect 2630 -590 2650 10
rect 2810 -590 2830 10
rect 2630 -610 2830 -590
rect 1770 -960 2150 -950
rect 2945 -970 2995 3188
rect 1350 -1070 1360 -1010
rect 1420 -1070 1430 -1010
rect 2279 -999 2331 -993
rect 2520 -1000 2995 -970
rect 2331 -1020 2995 -1000
rect 2331 -1050 2570 -1020
rect 2279 -1057 2331 -1051
rect 1350 -1080 1430 -1070
rect 2630 -1080 2830 -1060
rect 1220 -1170 1230 -1100
rect 1220 -1780 1300 -1170
rect 2630 -1320 2650 -1080
rect 2810 -1320 2830 -1080
rect 2630 -1340 2830 -1320
rect 1350 -1360 1430 -1350
rect 1350 -1420 1360 -1360
rect 1420 -1420 1430 -1360
rect 1350 -1700 1430 -1420
rect 2279 -1379 2331 -1373
rect 3135 -1380 3185 3188
rect 2331 -1430 3185 -1380
rect 2279 -1437 2331 -1431
rect 1680 -1470 2000 -1460
rect 1680 -1650 1690 -1470
rect 1760 -1650 2000 -1470
rect 1680 -1660 2000 -1650
rect 1350 -1760 1360 -1700
rect 1420 -1760 1430 -1700
rect 1350 -1770 1430 -1760
rect 1890 -1770 2000 -1660
rect 1220 -1850 1230 -1780
rect 1220 -2060 1300 -1850
rect 1220 -2130 1230 -2060
rect 1890 -2110 1900 -1770
rect 1990 -2110 2000 -1770
rect 1220 -2550 1300 -2130
rect 1350 -2140 1430 -2130
rect 1350 -2200 1360 -2140
rect 1420 -2200 1430 -2140
rect 1350 -2480 1430 -2200
rect 1890 -2240 2000 -2110
rect 1680 -2250 2000 -2240
rect 1680 -2430 1690 -2250
rect 1760 -2430 2000 -2250
rect 2830 -1580 3030 -1560
rect 2830 -2300 2850 -1580
rect 3010 -2300 3030 -1580
rect 2830 -2320 3030 -2300
rect 1680 -2440 2000 -2430
rect 1350 -2540 1360 -2480
rect 1420 -2540 1430 -2480
rect 2279 -2469 2331 -2463
rect 3305 -2470 3355 3188
rect 2331 -2520 3355 -2470
rect 2279 -2527 2331 -2521
rect 1350 -2550 1430 -2540
rect 1220 -2710 1230 -2550
rect 1220 -3090 1300 -2710
rect 2830 -2580 3030 -2560
rect 2830 -2700 2850 -2580
rect 3010 -2700 3030 -2580
rect 2830 -2720 3030 -2700
rect 1600 -2830 1610 -2770
rect 1680 -2830 1690 -2770
rect 1600 -3010 1690 -2830
rect 2309 -2789 2361 -2783
rect 3465 -2790 3515 3188
rect 2361 -2840 3515 -2790
rect 2309 -2847 2361 -2841
rect 1960 -2880 2280 -2870
rect 1960 -2960 1970 -2880
rect 2050 -2960 2280 -2880
rect 1960 -2970 2280 -2960
rect 1600 -3070 1610 -3010
rect 1680 -3070 1690 -3010
rect 1220 -3160 1230 -3090
rect 1220 -3320 1300 -3160
rect 1220 -3390 1230 -3320
rect 1220 -3730 1300 -3390
rect 2130 -3160 2280 -2970
rect 2130 -3320 2140 -3160
rect 2270 -3320 2280 -3160
rect 1600 -3470 1610 -3410
rect 1680 -3470 1690 -3410
rect 1600 -3650 1690 -3470
rect 2130 -3510 2280 -3320
rect 2830 -3020 3030 -3000
rect 2830 -3460 2850 -3020
rect 3010 -3460 3030 -3020
rect 2830 -3480 3030 -3460
rect 1960 -3520 2280 -3510
rect 1960 -3600 1970 -3520
rect 2050 -3600 2280 -3520
rect 1960 -3610 2280 -3600
rect 1600 -3710 1610 -3650
rect 1680 -3710 1690 -3650
rect 2304 -3639 2356 -3633
rect 3625 -3640 3675 3188
rect 2356 -3690 3675 -3640
rect 2304 -3697 2356 -3691
rect 1220 -3880 1230 -3730
rect 1220 -4250 1300 -3880
rect 2830 -3760 3030 -3740
rect 2830 -3880 2850 -3760
rect 3010 -3880 3030 -3760
rect 2830 -3900 3030 -3880
rect 1420 -3920 1500 -3910
rect 1420 -3980 1430 -3920
rect 1490 -3980 1500 -3920
rect 1420 -4160 1500 -3980
rect 2309 -3939 2361 -3933
rect 3765 -3940 3815 3188
rect 2361 -3990 3815 -3940
rect 2309 -3997 2361 -3991
rect 1780 -4030 2030 -4020
rect 1780 -4110 1790 -4030
rect 1870 -4110 2030 -4030
rect 1780 -4120 2030 -4110
rect 1420 -4220 1430 -4160
rect 1490 -4220 1500 -4160
rect 1420 -4230 1500 -4220
rect 1220 -4320 1230 -4250
rect 1220 -4480 1300 -4320
rect 1220 -4550 1230 -4480
rect 1220 -4910 1300 -4550
rect 1930 -4360 2030 -4120
rect 1930 -4440 1940 -4360
rect 2020 -4440 2030 -4360
rect 1420 -4580 1500 -4570
rect 1420 -4640 1430 -4580
rect 1490 -4640 1500 -4580
rect 1420 -4820 1500 -4640
rect 1930 -4680 2030 -4440
rect 2830 -4170 3030 -4150
rect 2830 -4630 2850 -4170
rect 3010 -4630 3030 -4170
rect 2830 -4650 3030 -4630
rect 1780 -4690 2030 -4680
rect 1780 -4770 1790 -4690
rect 1870 -4770 2030 -4690
rect 1780 -4780 2030 -4770
rect 1420 -4880 1430 -4820
rect 1490 -4880 1500 -4820
rect 2309 -4809 2361 -4803
rect 3915 -4810 3965 3188
rect 4050 2360 4250 2370
rect 4050 2280 4060 2360
rect 4240 2280 4250 2360
rect 4050 2270 4250 2280
rect 4620 2020 4820 3340
rect 6280 3250 6340 3256
rect 4620 1950 4630 2020
rect 4810 1950 4820 2020
rect 4330 1630 4530 1650
rect 4330 1550 4350 1630
rect 4510 1550 4530 1630
rect 4330 1530 4530 1550
rect 4050 830 4250 850
rect 4050 750 4070 830
rect 4230 750 4250 830
rect 4050 730 4250 750
rect 4620 440 4820 1950
rect 4620 350 4630 440
rect 4810 350 4820 440
rect 4330 30 4530 50
rect 4330 -50 4350 30
rect 4510 -50 4530 30
rect 4330 -70 4530 -50
rect 4050 -1530 4250 -1510
rect 4050 -1610 4070 -1530
rect 4230 -1610 4250 -1530
rect 4050 -1630 4250 -1610
rect 4620 -1920 4820 350
rect 4620 -2020 4630 -1920
rect 4810 -2020 4820 -1920
rect 4330 -2330 4530 -2310
rect 4330 -2410 4350 -2330
rect 4510 -2410 4530 -2330
rect 4330 -2430 4530 -2410
rect 2361 -4860 3965 -4810
rect 2309 -4867 2361 -4861
rect 1420 -4890 1500 -4880
rect 1220 -4980 1230 -4910
rect 1220 -4990 1300 -4980
rect 2830 -4920 3030 -4900
rect 2830 -5040 2850 -4920
rect 3010 -5040 3030 -4920
rect 2830 -5060 3030 -5040
rect 4620 -5150 4820 -2020
rect 4900 3149 5040 3160
rect 4900 3031 4911 3149
rect 5029 3031 5040 3149
rect 4900 2560 5040 3031
rect 5464 2966 5516 2972
rect 5464 2908 5516 2914
rect 5465 2715 5515 2908
rect 4900 2490 4910 2560
rect 5030 2490 5040 2560
rect 4900 2150 5040 2490
rect 4900 2080 4910 2150
rect 5030 2080 5040 2150
rect 4900 1890 5040 2080
rect 5075 2665 5515 2715
rect 5075 1965 5125 2665
rect 5730 2510 5830 2520
rect 5730 2430 5740 2510
rect 5820 2430 5830 2510
rect 5730 2370 5830 2430
rect 5500 2360 5830 2370
rect 5500 2280 5510 2360
rect 5580 2280 5830 2360
rect 5500 2270 5830 2280
rect 5075 1915 5680 1965
rect 4900 1820 4910 1890
rect 5030 1820 5040 1890
rect 5630 1876 5680 1915
rect 5623 1824 5629 1876
rect 5681 1824 5687 1876
rect 4900 1480 5040 1820
rect 5730 1700 5830 2270
rect 5500 1690 5830 1700
rect 5500 1610 5510 1690
rect 5580 1610 5830 1690
rect 5500 1600 5830 1610
rect 4900 1410 4910 1480
rect 5030 1410 5040 1480
rect 4900 1030 5040 1410
rect 6280 1300 6340 3190
rect 4900 970 4910 1030
rect 5030 970 5040 1030
rect 4900 610 5040 970
rect 5630 1240 6340 1300
rect 6420 3250 6480 3256
rect 5630 940 5690 1240
rect 6420 1170 6480 3190
rect 6828 3248 6888 3254
rect 6550 2550 6750 2570
rect 6550 1420 6570 2550
rect 6730 1420 6750 2550
rect 6550 1400 6750 1420
rect 5760 1110 6480 1170
rect 5620 930 5700 940
rect 5620 870 5630 930
rect 5690 870 5700 930
rect 5620 860 5700 870
rect 5630 720 5690 860
rect 5620 710 5700 720
rect 5620 650 5630 710
rect 5690 650 5700 710
rect 5620 640 5700 650
rect 4900 550 4910 610
rect 5030 550 5040 610
rect 4900 230 5040 550
rect 5760 270 5820 1110
rect 6550 1030 6750 1050
rect 4900 170 4910 230
rect 5030 170 5040 230
rect 4900 -190 5040 170
rect 5630 210 5820 270
rect 5880 980 6090 990
rect 5880 900 6000 980
rect 6080 900 6090 980
rect 5880 890 6090 900
rect 5880 820 5980 890
rect 5880 760 5890 820
rect 5970 760 5980 820
rect 5630 140 5690 210
rect 5620 130 5700 140
rect 5620 70 5630 130
rect 5690 70 5700 130
rect 5620 60 5700 70
rect 5630 -80 5690 60
rect 5880 20 5980 760
rect 5880 -40 5890 20
rect 5970 -40 5980 20
rect 5880 -50 5980 -40
rect 5620 -90 5700 -80
rect 5620 -150 5630 -90
rect 5690 -150 5700 -90
rect 5620 -160 5700 -150
rect 4900 -250 4910 -190
rect 5030 -250 5040 -190
rect 4900 -1330 5040 -250
rect 6550 -910 6570 1030
rect 6730 -910 6750 1030
rect 6550 -930 6750 -910
rect 6828 -1060 6888 3188
rect 4900 -1390 4910 -1330
rect 5030 -1390 5040 -1330
rect 4900 -1750 5040 -1390
rect 5630 -1120 6888 -1060
rect 6966 3248 7026 3254
rect 5630 -1420 5690 -1120
rect 6966 -1190 7026 3188
rect 5760 -1250 7026 -1190
rect 5620 -1430 5700 -1420
rect 5620 -1490 5630 -1430
rect 5690 -1490 5700 -1430
rect 5620 -1500 5700 -1490
rect 5630 -1640 5690 -1500
rect 5620 -1650 5700 -1640
rect 5620 -1710 5630 -1650
rect 5690 -1710 5700 -1650
rect 5620 -1720 5700 -1710
rect 4900 -1810 4910 -1750
rect 5030 -1810 5040 -1750
rect 4900 -2130 5040 -1810
rect 5760 -2090 5820 -1250
rect 6550 -1340 6750 -1320
rect 4900 -2190 4910 -2130
rect 5030 -2190 5040 -2130
rect 4900 -2550 5040 -2190
rect 5630 -2150 5820 -2090
rect 5880 -1380 5980 -1370
rect 5880 -1440 5890 -1380
rect 5970 -1440 5980 -1380
rect 5880 -1540 5980 -1440
rect 5880 -1600 5890 -1540
rect 5970 -1600 5980 -1540
rect 5630 -2220 5690 -2150
rect 5620 -2230 5700 -2220
rect 5620 -2290 5630 -2230
rect 5690 -2290 5700 -2230
rect 5620 -2300 5700 -2290
rect 5630 -2440 5690 -2300
rect 5880 -2340 5980 -1600
rect 5880 -2400 5890 -2340
rect 5970 -2400 5980 -2340
rect 5880 -2410 5980 -2400
rect 5620 -2450 5700 -2440
rect 5620 -2510 5630 -2450
rect 5690 -2510 5700 -2450
rect 5620 -2520 5700 -2510
rect 4900 -2610 4910 -2550
rect 5030 -2610 5040 -2550
rect 4900 -2620 5040 -2610
rect 6550 -4870 6570 -1340
rect 6730 -4870 6750 -1340
rect 6550 -4890 6750 -4870
rect 890 -5155 6390 -5150
rect 890 -5345 6175 -5155
rect 6365 -5345 6390 -5155
rect 890 -5350 6390 -5345
rect 5080 -5900 5300 -5890
rect 5080 -6100 5090 -5900
rect 5290 -6100 5300 -5900
rect 5080 -6110 5300 -6100
rect 150 -6150 1330 -6140
rect 150 -6600 160 -6150
rect 1320 -6600 1330 -6150
rect 150 -6610 1330 -6600
rect 3880 -6160 5050 -6150
rect 3880 -6600 3890 -6160
rect 5040 -6600 5050 -6160
rect 3880 -6610 5050 -6600
<< via2 >>
rect 440 4020 720 4180
rect 1180 3600 1470 3800
rect 1730 3620 2020 3780
rect 630 1980 790 2520
rect 310 970 470 1510
rect 630 10 790 360
rect 310 -940 470 -590
rect 630 -1640 790 -1480
rect 310 -2420 470 -2260
rect 630 -2990 790 -2850
rect 310 -3610 470 -3510
rect 630 -4120 790 -4020
rect 310 -4780 470 -4680
rect 2650 490 2810 560
rect 2650 -590 2810 10
rect 2650 -1320 2810 -1080
rect 2850 -2300 3010 -1580
rect 2850 -2700 3010 -2580
rect 2850 -3460 3010 -3020
rect 2850 -3880 3010 -3760
rect 2850 -4630 3010 -4170
rect 4060 2280 4240 2360
rect 4350 1550 4510 1630
rect 4070 750 4220 830
rect 4220 750 4230 830
rect 4350 -50 4510 30
rect 4070 -1610 4220 -1530
rect 4220 -1610 4230 -1530
rect 4350 -2410 4510 -2330
rect 2850 -5040 3010 -4920
rect 4911 3031 5029 3149
rect 6570 1420 6730 2550
rect 6570 -910 6730 1030
rect 6570 -4870 6730 -1340
rect 6175 -5345 6365 -5155
rect 5095 -6095 5285 -5905
rect 160 -6600 1320 -6150
rect 3890 -6600 5040 -6160
<< metal3 >>
rect 420 4180 740 4200
rect 420 4020 440 4180
rect 720 4020 740 4180
rect 420 3400 740 4020
rect 1160 3800 1490 3820
rect 1160 3600 1180 3800
rect 1470 3780 6750 3800
rect 1470 3620 1730 3780
rect 2020 3620 6750 3780
rect 1470 3600 6750 3620
rect 1160 3580 1490 3600
rect 420 3240 440 3400
rect 720 3240 740 3400
rect 420 3220 740 3240
rect 610 2520 810 2540
rect 610 1980 630 2520
rect 790 1980 810 2520
rect 290 1510 490 1530
rect 290 970 310 1510
rect 470 970 490 1510
rect 290 950 490 970
rect 610 360 810 1980
rect 610 10 630 360
rect 790 10 810 360
rect 290 -590 490 -570
rect 290 -940 310 -590
rect 470 -940 490 -590
rect 290 -960 490 -940
rect 610 -1480 810 10
rect 2630 560 2830 3600
rect 4906 3149 5034 3600
rect 4906 3031 4911 3149
rect 5029 3031 5034 3149
rect 4906 3026 5034 3031
rect 6550 2550 6750 3600
rect 2630 490 2650 560
rect 2810 490 2830 560
rect 2630 10 2830 490
rect 2630 -590 2650 10
rect 2810 -590 2830 10
rect 2630 -1080 2830 -590
rect 2630 -1320 2650 -1080
rect 2810 -1280 2830 -1080
rect 4050 2360 4250 2370
rect 4050 2280 4060 2360
rect 4240 2280 4250 2360
rect 4050 830 4250 2280
rect 4330 1630 4530 1650
rect 4330 1550 4350 1630
rect 4510 1550 4530 1630
rect 4330 1530 4530 1550
rect 4050 750 4070 830
rect 4230 750 4250 830
rect 2810 -1320 3030 -1280
rect 2630 -1480 3030 -1320
rect 610 -1640 630 -1480
rect 790 -1640 810 -1480
rect 290 -2260 490 -2240
rect 290 -2420 310 -2260
rect 470 -2420 490 -2260
rect 290 -2440 490 -2420
rect 610 -2850 810 -1640
rect 610 -2990 630 -2850
rect 790 -2990 810 -2850
rect 290 -3510 490 -3490
rect 290 -3610 310 -3510
rect 470 -3610 490 -3510
rect 290 -3630 490 -3610
rect 610 -4020 810 -2990
rect 610 -4120 630 -4020
rect 790 -4120 810 -4020
rect 290 -4680 490 -4660
rect 290 -4780 310 -4680
rect 470 -4780 490 -4680
rect 290 -4800 490 -4780
rect 610 -5430 810 -4120
rect 2830 -1580 3030 -1480
rect 2830 -2300 2850 -1580
rect 3010 -2300 3030 -1580
rect 2830 -2580 3030 -2300
rect 2830 -2700 2850 -2580
rect 3010 -2700 3030 -2580
rect 2830 -3020 3030 -2700
rect 2830 -3460 2850 -3020
rect 3010 -3460 3030 -3020
rect 2830 -3760 3030 -3460
rect 2830 -3880 2850 -3760
rect 3010 -3880 3030 -3760
rect 2830 -4170 3030 -3880
rect 2830 -4630 2850 -4170
rect 3010 -4630 3030 -4170
rect 2830 -4920 3030 -4630
rect 2830 -5040 2850 -4920
rect 3010 -5040 3030 -4920
rect 2830 -5060 3030 -5040
rect 4050 -1530 4250 750
rect 6550 1420 6570 2550
rect 6730 1420 6750 2550
rect 6550 1030 6750 1420
rect 4330 30 4530 50
rect 4330 -50 4350 30
rect 4510 -50 4530 30
rect 4330 -70 4530 -50
rect 4050 -1610 4070 -1530
rect 4230 -1610 4250 -1530
rect 4050 -5430 4250 -1610
rect 6550 -910 6570 1030
rect 6730 -910 6750 1030
rect 6550 -1340 6750 -910
rect 4330 -2330 4530 -2310
rect 4330 -2410 4350 -2330
rect 4510 -2410 4530 -2330
rect 4330 -2430 4530 -2410
rect 6550 -4870 6570 -1340
rect 6730 -4870 6750 -1340
rect 6171 -5150 6369 -5145
rect 6170 -5151 6370 -5150
rect 6170 -5349 6171 -5151
rect 6369 -5349 6370 -5151
rect 6170 -5350 6370 -5349
rect 6171 -5355 6369 -5350
rect 610 -5630 5880 -5430
rect 6080 -5630 6086 -5430
rect 6550 -5900 6750 -4870
rect 5090 -5905 6750 -5900
rect 5090 -6095 5095 -5905
rect 5285 -6095 6750 -5905
rect 5090 -6100 6750 -6095
rect 150 -6150 1330 -6140
rect 150 -6600 160 -6150
rect 1320 -6600 1330 -6150
rect 150 -6610 1330 -6600
rect 3880 -6160 5050 -6150
rect 3880 -6600 3890 -6160
rect 5040 -6600 5050 -6160
rect 3880 -6610 5050 -6600
<< via3 >>
rect 440 4020 720 4180
rect 1180 3600 1470 3800
rect 440 3240 720 3400
rect 310 970 470 1510
rect 310 -940 470 -590
rect 4350 1550 4510 1630
rect 310 -2420 470 -2260
rect 310 -3610 470 -3510
rect 310 -4780 470 -4680
rect 4350 -50 4510 30
rect 4350 -2410 4510 -2330
rect 6171 -5155 6369 -5151
rect 6171 -5345 6175 -5155
rect 6175 -5345 6365 -5155
rect 6365 -5345 6369 -5155
rect 6171 -5349 6369 -5345
rect 5880 -5630 6080 -5430
rect 160 -6600 1320 -6150
rect 3890 -6600 5040 -6160
<< metal4 >>
rect 0 4180 740 4200
rect 0 4020 440 4180
rect 720 4020 740 4180
rect 0 4000 740 4020
rect 1160 3800 1490 3820
rect 0 3600 1180 3800
rect 1470 3600 1490 3800
rect 1160 3580 1490 3600
rect 0 3400 740 3420
rect 0 3240 440 3400
rect 720 3240 740 3400
rect 0 3220 740 3240
rect 0 -6110 200 3220
rect 4330 1630 4530 1650
rect 4330 1550 4350 1630
rect 4510 1550 4530 1630
rect 290 1510 490 1530
rect 290 970 310 1510
rect 470 970 490 1510
rect 290 -590 490 970
rect 290 -940 310 -590
rect 470 -940 490 -590
rect 290 -2260 490 -940
rect 290 -2420 310 -2260
rect 470 -2420 490 -2260
rect 290 -3510 490 -2420
rect 290 -3610 310 -3510
rect 470 -3610 490 -3510
rect 290 -4680 490 -3610
rect 290 -4780 310 -4680
rect 470 -4780 490 -4680
rect 290 -5710 490 -4780
rect 4330 30 4530 1550
rect 4330 -50 4350 30
rect 4510 -50 4530 30
rect 4330 -2330 4530 -50
rect 4330 -2410 4350 -2330
rect 4510 -2410 4530 -2330
rect 4330 -5710 4530 -2410
rect 6170 -5151 6500 -5150
rect 6170 -5349 6171 -5151
rect 6369 -5349 6500 -5151
rect 6170 -5350 6500 -5349
rect 5879 -5430 6081 -5429
rect 5879 -5630 5880 -5430
rect 6080 -5630 6081 -5430
rect 5879 -5631 6081 -5630
rect 290 -5910 4530 -5710
rect 0 -6150 1360 -6110
rect 4330 -6150 4530 -5910
rect 0 -6600 160 -6150
rect 1320 -6600 1360 -6150
rect 0 -6650 1360 -6600
rect 3880 -6160 5050 -6150
rect 3880 -6600 3890 -6160
rect 5040 -6320 5050 -6160
rect 5040 -6520 5660 -6320
rect 5040 -6600 5050 -6520
rect 3880 -6610 5050 -6600
rect 5460 -8010 5660 -6520
rect 5880 -8010 6080 -5631
rect 6300 -8010 6500 -5350
use sky130_fd_pr__nfet_01v8_ATLS57  sky130_fd_pr__nfet_01v8_ATLS57_0 csdac_nom__devices
timestamp 1723780759
transform -1 0 1651 0 -1 -770
box -211 -410 211 410
use sky130_fd_pr__nfet_01v8_HZS9GD  XMB0 csdac_nom__devices
timestamp 1723780759
transform 0 1 6140 -1 0 -3104
box -1796 -260 1796 260
use sky130_fd_pr__nfet_01v8_FMHZDY  XMB1 csdac_nom__devices
timestamp 1723780759
transform 0 1 6140 -1 0 56
box -996 -260 996 260
use sky130_fd_pr__nfet_01v8_AHZR5K  XMB2 csdac_nom__devices
timestamp 1723780759
transform 0 1 6030 -1 0 1986
box -596 -260 596 260
use sky130_fd_pr__nfet_01v8_BHEWB6  XMB3 csdac_nom__devices
timestamp 1723780759
transform 1 0 2416 0 1 -4400
box -406 -260 406 260
use sky130_fd_pr__nfet_01v8_FMMQLY  XMB4 csdac_nom__devices
timestamp 1723780759
transform 1 0 2486 0 1 -3240
box -296 -260 296 260
use sky130_fd_pr__nfet_01v8_C4RU6Y  XMB5 csdac_nom__devices
timestamp 1723780759
transform 1 0 2346 0 1 -1940
box -426 -400 426 400
use sky130_fd_pr__nfet_01v8_N5FCK4  XMB6 csdac_nom__devices
timestamp 1723780759
transform 1 0 2336 0 1 -290
box -246 -320 246 320
use sky130_fd_pr__nfet_01v8_8TEC39  XMB7 csdac_nom__devices
timestamp 1723780759
transform 0 -1 1860 1 0 3006
box -246 -420 246 420
use sky130_fd_pr__nfet_01v8_SMGLWN  XMmirror csdac_nom__devices
timestamp 1723780759
transform 1 0 1105 0 1 4507
box -246 -260 246 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMN0 csdac_nom__devices
timestamp 1723780759
transform 1 0 5421 0 1 -1570
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMN1
timestamp 1723780759
transform 1 0 5421 0 1 790
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMN2
timestamp 1723780759
transform 1 0 5381 0 1 2320
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMN3
timestamp 1723780759
transform 1 0 1631 0 1 -4070
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMN4
timestamp 1723780759
transform 1 0 1831 0 1 -2920
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_648S5X  XMN5 csdac_nom__devices
timestamp 1723780759
transform 1 0 1561 0 1 -1560
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_ATLS57  XMN6
timestamp 1723780759
transform -1 0 1651 0 -1 180
box -211 -410 211 410
use sky130_fd_pr__nfet_01v8_J2SMEF  XMN7 csdac_nom__devices
timestamp 1723780759
transform 1 0 1651 0 1 2250
box -211 -510 211 510
use sky130_fd_pr__nfet_01v8_L9ESAD  XMP0
timestamp 1723780759
transform 1 0 5421 0 1 -2370
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMP1
timestamp 1723780759
transform 1 0 5421 0 1 -10
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMP2
timestamp 1723780759
transform 1 0 5381 0 1 1650
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMP3
timestamp 1723780759
transform 1 0 1631 0 1 -4730
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMP4
timestamp 1723780759
transform 1 0 1831 0 1 -3560
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_648S5X  XMP5
timestamp 1723780759
transform 1 0 1561 0 1 -2340
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_J2SMEF  XMP7
timestamp 1723780759
transform 1 0 1651 0 1 1240
box -211 -510 211 510
use sky130_fd_pr__pfet_01v8_XJ7GBL  XMprog csdac_nom__devices
timestamp 1723780759
transform 1 0 631 0 1 4509
box -211 -269 211 269
use sky130_fd_pr__res_high_po_5p73_3RZNGL  XR5
timestamp 1724299458
transform 1 0 2602 0 -1 -7003
box -2602 -1007 2602 1007
<< labels >>
flabel metal4 0 4000 300 4200 0 FreeSans 1120 0 0 0 vcc
port 21 nsew
flabel metal4 0 3600 300 3800 0 FreeSans 1120 0 0 0 vss
port 22 nsew
flabel metal1 1400 4920 1492 5196 0 FreeSans 640 0 0 0 n7
port 26 nsew
flabel metal1 3976 4920 4068 5196 0 FreeSans 640 0 0 0 p4
port 33 nsew
flabel metal1 4344 4920 4436 5196 0 FreeSans 640 0 0 0 n3
port 34 nsew
flabel metal1 4712 4920 4804 5196 0 FreeSans 640 0 0 0 p3
port 35 nsew
flabel metal1 5080 4920 5172 5196 0 FreeSans 640 0 0 0 n2
port 36 nsew
flabel metal1 5448 4920 5540 5196 0 FreeSans 640 0 0 0 p2
port 37 nsew
flabel metal1 6552 4920 6644 5196 0 FreeSans 640 0 0 0 n0
port 40 nsew
flabel metal1 6920 4920 7012 5196 0 FreeSans 640 0 0 0 p0
port 41 nsew
flabel metal1 6184 4920 6276 5196 0 FreeSans 640 0 0 0 p1
port 39 nsew
flabel metal1 5816 4920 5908 5196 0 FreeSans 640 0 0 0 n1
port 38 nsew
flabel metal1 3608 4920 3700 5196 0 FreeSans 640 0 0 0 n4
port 32 nsew
flabel metal1 3240 4920 3332 5196 0 FreeSans 640 0 0 0 p5
port 31 nsew
flabel metal1 2872 4920 2964 5196 0 FreeSans 640 0 0 0 n5
port 30 nsew
flabel metal1 2504 4920 2596 5196 0 FreeSans 640 0 0 0 p6
port 29 nsew
flabel metal1 2136 4920 2228 5196 0 FreeSans 640 0 0 0 n6
port 28 nsew
flabel metal1 1768 4920 1860 5196 0 FreeSans 640 0 0 0 p7
port 27 nsew
flabel metal1 1850 950 2060 2950 0 FreeSans 800 0 0 0 IS7
flabel metal2 2000 -200 2150 370 0 FreeSans 800 0 0 0 IS6
flabel metal2 1760 -1660 2000 -1460 0 FreeSans 800 0 0 0 IS5
flabel metal2 2130 -3160 2280 -2870 0 FreeSans 800 0 0 0 IS4
flabel metal2 1930 -4360 2030 -4020 0 FreeSans 800 0 0 0 IS3
flabel metal2 5880 -2340 5980 -1600 0 FreeSans 800 0 0 0 IS0
flabel metal2 5880 20 5980 760 0 FreeSans 800 0 0 0 IS1
flabel metal2 5580 2270 5830 2370 0 FreeSans 800 0 0 0 IS2
flabel metal4 5880 -8010 6080 -7810 0 FreeSans 640 0 0 0 Vneg
port 42 nsew
flabel metal4 5460 -8010 5660 -7810 0 FreeSans 640 0 0 0 Vpos
port 43 nsew
flabel metal4 6300 -8010 6500 -7810 0 FreeSans 640 0 0 0 Vbias
port 44 nsew
<< end >>

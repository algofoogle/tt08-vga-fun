magic
tech sky130A
magscale 1 2
timestamp 1725599052
<< viali >>
rect -1470 4780 -1420 4970
rect -510 4890 -450 4970
rect 40 4790 190 4830
rect 500 4790 600 4830
rect 910 4800 1010 4840
rect -600 4370 -540 4450
rect -1280 3690 -1230 3960
rect 190 3890 340 4570
rect 700 3890 850 4570
rect 1220 3920 1260 4640
rect 1980 4240 2020 4410
rect 2500 4240 2540 4410
rect 1370 4070 1420 4140
rect 1890 3980 1930 4140
rect 2590 3970 2630 4140
rect 1920 3400 2000 3560
rect 2120 3420 2400 3480
rect 2540 3400 2620 3560
rect -1110 2240 -630 2280
rect 350 2240 830 2280
rect 1480 2250 1660 2290
rect 2090 2250 2270 2290
rect 2700 2250 2880 2290
rect 1810 1950 1940 2010
rect 2420 1950 2550 2010
rect -380 1790 100 1830
rect 1770 1450 1900 1610
rect 2460 1450 2590 1610
rect -1400 1100 -1360 1290
rect 1080 1110 1120 1280
rect -650 910 -480 1060
rect 200 910 370 1060
<< metal1 >>
rect 1230 5390 1400 5400
rect -1310 5380 -1190 5390
rect -1310 5280 -1300 5380
rect -1200 5280 -1190 5380
rect -1310 5270 -1190 5280
rect -1010 5380 -890 5390
rect -1010 5280 -1000 5380
rect -900 5280 -890 5380
rect 1230 5360 1240 5390
rect -1010 5270 -890 5280
rect 210 5270 1240 5360
rect -1300 5020 -1200 5270
rect -1010 5170 -670 5270
rect -1500 4970 -1310 4980
rect -1500 4780 -1470 4970
rect -1420 4880 -1310 4970
rect -1420 4780 -1400 4880
rect -1280 4800 -1230 5020
rect -1200 4880 -830 4980
rect -1500 3530 -1400 4780
rect -1170 4650 -1110 4880
rect -770 4800 -670 5170
rect 70 5170 150 5180
rect 70 5110 80 5170
rect 140 5110 150 5170
rect 210 5070 300 5270
rect 480 5170 560 5180
rect 480 5110 490 5170
rect 550 5110 560 5170
rect 492 5108 504 5110
rect 538 5108 550 5110
rect 492 5102 550 5108
rect 620 5070 710 5270
rect 890 5180 970 5190
rect 890 5120 900 5180
rect 960 5120 970 5180
rect 902 5118 914 5120
rect 948 5118 960 5120
rect 902 5112 960 5118
rect 1030 5080 1120 5270
rect 1230 5240 1240 5270
rect 1390 5240 1400 5390
rect 1230 5230 1400 5240
rect 1550 5390 1750 5400
rect -110 4980 90 5070
rect 140 4980 300 5070
rect -620 4970 -270 4980
rect -620 4890 -510 4970
rect -450 4890 -270 4970
rect -620 4880 -270 4890
rect -1220 4590 -1110 4650
rect -530 4600 -410 4610
rect -1220 4460 -1160 4590
rect -530 4560 -520 4600
rect -1100 4500 -520 4560
rect -420 4500 -410 4600
rect -1220 4360 -1120 4460
rect -1220 4160 -1160 4360
rect -950 4320 -870 4500
rect -530 4490 -410 4500
rect -370 4460 -270 4880
rect -110 4740 -10 4980
rect 350 4970 500 5070
rect 542 5058 710 5070
rect 542 4982 548 5058
rect 550 4982 710 5058
rect 542 4980 710 4982
rect 760 4980 910 5080
rect 952 5068 1120 5080
rect 952 4992 958 5068
rect 960 4992 1120 5068
rect 952 4980 1120 4992
rect 1550 5170 1560 5390
rect 1740 5170 1750 5390
rect 542 4970 560 4980
rect 70 4880 80 4940
rect 140 4880 150 4940
rect 70 4870 150 4880
rect 20 4830 240 4840
rect 20 4790 40 4830
rect 190 4790 240 4830
rect 20 4770 240 4790
rect -110 4640 60 4740
rect -40 4580 60 4640
rect 180 4590 240 4770
rect 350 4740 450 4970
rect 480 4880 490 4940
rect 550 4880 560 4940
rect 480 4870 560 4880
rect 480 4830 730 4840
rect 480 4790 500 4830
rect 600 4790 730 4830
rect 480 4770 730 4790
rect 350 4640 570 4740
rect 470 4590 570 4640
rect 680 4590 730 4770
rect 760 4740 860 4980
rect 890 4890 900 4950
rect 960 4890 970 4950
rect 890 4880 970 4890
rect 890 4840 1280 4850
rect 890 4800 910 4840
rect 1010 4800 1280 4840
rect 890 4780 1280 4800
rect 760 4640 1080 4740
rect 1110 4680 1280 4780
rect -700 4450 -270 4460
rect -700 4370 -600 4450
rect -540 4370 -270 4450
rect -700 4360 -270 4370
rect 180 4570 350 4590
rect -670 4330 -520 4360
rect -1120 4270 -710 4320
rect -1220 4100 -1050 4160
rect -1500 3450 -1490 3530
rect -1410 3450 -1400 3530
rect -1500 3440 -1400 3450
rect -1310 3960 -1210 3980
rect -1310 3690 -1280 3960
rect -1230 3880 -1210 3960
rect -1110 3970 -1050 4100
rect -640 4140 -520 4330
rect -640 4014 -520 4020
rect -1110 3910 -950 3970
rect -1230 3780 -1120 3880
rect -1090 3810 -240 3910
rect 180 3890 190 4570
rect 340 3890 350 4570
rect 180 3870 350 3890
rect 690 4570 860 4590
rect 980 4580 1080 4640
rect 1200 4640 1280 4680
rect 690 3890 700 4570
rect 850 3890 860 4570
rect 1200 3990 1220 4640
rect 1260 4160 1280 4640
rect 1440 4280 1520 4290
rect 1440 4220 1450 4280
rect 1510 4220 1520 4280
rect 1440 4210 1520 4220
rect 1450 4190 1520 4210
rect 1550 4200 1750 5170
rect 2160 5390 2360 5400
rect 2160 5170 2170 5390
rect 2350 5170 2360 5390
rect 1890 4410 2040 4430
rect 1780 4280 1860 4290
rect 1780 4220 1790 4280
rect 1850 4220 1860 4280
rect 1780 4210 1860 4220
rect 1890 4240 1980 4410
rect 2020 4240 2040 4410
rect 1260 4140 1430 4160
rect 1260 4070 1370 4140
rect 1420 4070 1430 4140
rect 1460 4120 1520 4190
rect 1780 4190 1850 4210
rect 1260 4050 1430 4070
rect 1260 4000 1280 4050
rect 1260 3990 1310 4000
rect 1200 3900 1210 3990
rect 1300 3900 1310 3990
rect 1550 3960 1750 4130
rect 1780 4120 1840 4190
rect 1890 4170 2040 4240
rect 1890 4160 1910 4170
rect 1870 4140 1910 4160
rect 1200 3890 1310 3900
rect 1380 3950 1750 3960
rect 1870 3980 1890 4140
rect 2010 4120 2040 4170
rect 2070 4220 2130 4390
rect 2160 4370 2360 5170
rect 2770 5390 2970 5400
rect 2770 5170 2780 5390
rect 2960 5170 2970 5390
rect 2480 4410 2630 4430
rect 2070 4210 2150 4220
rect 2070 4150 2080 4210
rect 2140 4150 2150 4210
rect 2070 4140 2150 4150
rect 2010 4070 2020 4120
rect 1930 4060 2020 4070
rect 1930 3980 1990 4060
rect 1870 3950 1990 3980
rect 690 3870 860 3890
rect 1380 3850 1390 3950
rect 1490 3850 1750 3950
rect 2200 3860 2320 4290
rect 2390 4220 2450 4390
rect 2370 4210 2450 4220
rect 2370 4150 2380 4210
rect 2440 4150 2450 4210
rect 2370 4140 2450 4150
rect 2480 4240 2500 4410
rect 2540 4240 2630 4410
rect 2480 4170 2630 4240
rect 2660 4280 2740 4290
rect 2660 4220 2670 4280
rect 2730 4220 2740 4280
rect 2660 4210 2740 4220
rect 2670 4190 2740 4210
rect 2770 4200 2970 5170
rect 3000 4280 3080 4290
rect 3000 4220 3010 4280
rect 3070 4220 3080 4280
rect 3000 4210 3080 4220
rect 2480 4120 2510 4170
rect 2610 4160 2630 4170
rect 2610 4140 2650 4160
rect 2500 4070 2510 4120
rect 2500 4060 2590 4070
rect 2560 3970 2590 4060
rect 2630 3970 2650 4140
rect 2680 4120 2740 4190
rect 3000 4190 3070 4210
rect 2560 3950 2650 3970
rect 2770 3960 2970 4130
rect 3000 4120 3060 4190
rect 2770 3950 3140 3960
rect 1380 3840 1750 3850
rect 2770 3850 3030 3950
rect 3130 3850 3140 3950
rect 2770 3840 3140 3850
rect -1230 3690 -1210 3780
rect -1090 3750 3860 3810
rect -1110 3700 -950 3750
rect -1090 3690 -950 3700
rect -1310 3010 -1210 3690
rect -410 3650 3860 3750
rect 210 3590 320 3600
rect -40 3340 60 3570
rect 210 3500 220 3590
rect 310 3500 320 3590
rect 720 3590 830 3600
rect 210 3340 320 3500
rect 470 3340 570 3570
rect 720 3500 730 3590
rect 820 3500 830 3590
rect 1380 3580 1560 3600
rect 720 3340 830 3500
rect 980 3480 1080 3570
rect 1380 3500 1400 3580
rect 1480 3500 1560 3580
rect 1380 3480 1560 3500
rect 980 3470 1310 3480
rect 980 3380 1210 3470
rect 1300 3380 1310 3470
rect 1640 3420 1760 3650
rect 1840 3590 2020 3600
rect 1840 3490 1910 3590
rect 2010 3540 2020 3590
rect 2500 3590 2680 3600
rect 2200 3540 2320 3560
rect 2500 3540 2510 3590
rect 2610 3560 2680 3590
rect 2010 3490 2510 3540
rect 1840 3480 1920 3490
rect 980 3340 1310 3380
rect 1900 3400 1920 3480
rect 2000 3480 2540 3490
rect 2000 3420 2120 3480
rect 2400 3420 2540 3480
rect 2000 3400 2540 3420
rect 2620 3480 2680 3560
rect 2620 3400 2640 3480
rect 2780 3420 2900 3650
rect 2980 3580 3160 3600
rect 2980 3500 3060 3580
rect 3140 3500 3160 3580
rect 2980 3480 3160 3500
rect 1900 3360 2640 3400
rect -40 3210 1310 3340
rect -1310 2930 -1300 3010
rect -1220 2930 -1210 3010
rect -1310 2920 -1210 2930
rect 420 3010 620 3210
rect 420 2830 430 3010
rect 610 2830 620 3010
rect 420 2820 620 2830
rect 2040 3010 2480 3360
rect 2040 2630 2050 3010
rect 2470 2630 2480 3010
rect 2040 2620 2480 2630
rect 3700 2511 3860 3650
rect -1901 2349 3861 2511
rect -1210 2050 -1160 2349
rect -1130 2300 -610 2310
rect -1130 2230 -1120 2300
rect -620 2230 -610 2300
rect -1130 2140 -610 2230
rect -1430 1310 -1350 1320
rect -1430 1080 -1420 1310
rect -1360 1080 -1350 1310
rect -1130 1250 -610 2030
rect -581 1680 -529 2349
rect -400 1850 120 1860
rect -400 1780 -390 1850
rect 110 1780 120 1850
rect -400 1690 120 1780
rect 250 1680 300 2349
rect 330 2300 850 2310
rect 330 2230 340 2300
rect 840 2230 850 2300
rect 330 2140 850 2230
rect 880 2050 930 2349
rect 1460 2300 1680 2310
rect 1460 2230 1470 2300
rect 1670 2230 1680 2300
rect 1460 2150 1680 2230
rect 1845 2100 1895 2349
rect 2070 2300 2290 2310
rect 2070 2230 2080 2300
rect 2280 2230 2290 2300
rect 2070 2150 2290 2230
rect 2455 2100 2505 2349
rect 2680 2300 2900 2310
rect 2680 2230 2690 2300
rect 2890 2230 2900 2300
rect 2680 2150 2900 2230
rect 1390 2050 2960 2100
rect -581 1594 -430 1680
rect -580 1590 -430 1594
rect -1320 1230 -1250 1240
rect -1320 1160 -1310 1230
rect -1320 1150 -1250 1160
rect -530 1230 -460 1240
rect -470 1160 -460 1230
rect -530 1150 -460 1160
rect -1430 1070 -1350 1080
rect -1210 360 -690 1140
rect -660 1080 -450 1090
rect -460 890 -450 1080
rect -660 880 -450 890
rect -400 830 120 1610
rect 150 1590 300 1680
rect 250 1585 300 1590
rect 330 1250 850 2030
rect 1790 2010 1960 2020
rect 1460 1850 1680 2000
rect 1790 1950 1800 2010
rect 1940 1950 1960 2010
rect 2400 2010 2570 2020
rect 1790 1940 1960 1950
rect 1370 1740 1680 1850
rect 1250 1560 1320 1580
rect 1370 1570 1610 1740
rect 1760 1610 1910 1630
rect 1250 1500 1260 1560
rect 1250 1480 1320 1500
rect 1660 1560 1730 1580
rect 1720 1500 1730 1560
rect 1070 1300 1150 1310
rect 170 1230 250 1240
rect 170 1160 190 1230
rect 170 1150 250 1160
rect 970 1230 1040 1240
rect 1030 1160 1040 1230
rect 970 1150 1040 1160
rect 170 1080 380 1090
rect 170 890 180 1080
rect 170 880 380 890
rect -570 810 -500 820
rect -570 740 -560 810
rect -570 730 -500 740
rect 220 810 290 820
rect 280 740 290 810
rect 220 730 290 740
rect -1210 -20 -1190 360
rect -710 -20 -690 360
rect -1210 -40 -690 -20
rect -400 360 120 720
rect -400 -20 -380 360
rect 100 -20 120 360
rect -400 -40 120 -20
rect 410 360 930 1140
rect 1070 1090 1080 1300
rect 1140 1090 1150 1300
rect 1070 1080 1150 1090
rect 410 -20 430 360
rect 910 -20 930 360
rect 410 -40 930 -20
rect 1370 360 1610 1490
rect 1660 1480 1730 1500
rect 1760 1450 1770 1610
rect 1900 1450 1910 1610
rect 1940 1560 2010 1580
rect 2080 1570 2280 2000
rect 2400 1950 2420 2010
rect 2560 1950 2570 2010
rect 2400 1940 2570 1950
rect 2680 1850 2900 2000
rect 2680 1740 2990 1850
rect 2450 1610 2600 1630
rect 1940 1500 1950 1560
rect 1940 1480 2010 1500
rect 2350 1560 2420 1580
rect 2410 1500 2420 1560
rect 2350 1480 2420 1500
rect 1760 1430 1910 1450
rect 1370 -20 1390 360
rect 1590 -20 1610 360
rect 1370 -40 1610 -20
rect 2060 360 2300 1480
rect 2450 1450 2460 1610
rect 2590 1450 2600 1610
rect 2630 1560 2700 1580
rect 2750 1570 2990 1740
rect 2630 1500 2640 1560
rect 2630 1480 2700 1500
rect 3040 1560 3110 1580
rect 3100 1500 3110 1560
rect 3040 1480 3110 1500
rect 2450 1430 2600 1450
rect 2060 -20 2080 360
rect 2280 -20 2300 360
rect 2060 -40 2300 -20
rect 2750 360 2990 1480
rect 2750 -20 2770 360
rect 2970 -20 2990 360
rect 2750 -40 2990 -20
<< via1 >>
rect -1300 5280 -1200 5380
rect -1000 5280 -900 5380
rect 80 5110 140 5170
rect 490 5110 550 5170
rect 900 5120 960 5180
rect 1240 5240 1390 5390
rect -520 4500 -420 4600
rect 1560 5170 1740 5390
rect 80 4880 140 4940
rect 490 4880 550 4940
rect 900 4890 960 4950
rect -1490 3450 -1410 3530
rect -640 4020 -520 4140
rect 220 3940 310 4030
rect 730 3940 820 4030
rect 1450 4220 1510 4280
rect 2170 5170 2350 5390
rect 1790 4220 1850 4280
rect 1210 3920 1220 3990
rect 1220 3920 1260 3990
rect 1260 3920 1300 3990
rect 1210 3900 1300 3920
rect 1910 4140 2010 4170
rect 1910 4070 1930 4140
rect 1930 4070 2010 4140
rect 2780 5170 2960 5390
rect 2080 4150 2140 4210
rect 1390 3850 1490 3950
rect 2380 4150 2440 4210
rect 2670 4220 2730 4280
rect 3010 4220 3070 4280
rect 2510 4140 2610 4170
rect 2510 4070 2590 4140
rect 2590 4070 2610 4140
rect 3030 3850 3130 3950
rect 220 3500 310 3590
rect 730 3500 820 3590
rect 1400 3500 1480 3580
rect 1210 3380 1300 3470
rect 1910 3560 2010 3590
rect 1910 3490 1920 3560
rect 1920 3490 2000 3560
rect 2000 3490 2010 3560
rect 2510 3560 2610 3590
rect 2510 3490 2540 3560
rect 2540 3490 2610 3560
rect 3060 3500 3140 3580
rect -1300 2930 -1220 3010
rect 430 2830 610 3010
rect 2050 2630 2470 3010
rect -1120 2280 -620 2300
rect -1120 2240 -1110 2280
rect -1110 2240 -630 2280
rect -630 2240 -620 2280
rect -1120 2230 -620 2240
rect -1420 1290 -1360 1310
rect -1420 1100 -1400 1290
rect -1400 1100 -1360 1290
rect -1420 1080 -1360 1100
rect -390 1830 110 1850
rect -390 1790 -380 1830
rect -380 1790 100 1830
rect 100 1790 110 1830
rect -390 1780 110 1790
rect 340 2280 840 2300
rect 340 2240 350 2280
rect 350 2240 830 2280
rect 830 2240 840 2280
rect 340 2230 840 2240
rect 1470 2290 1670 2300
rect 1470 2250 1480 2290
rect 1480 2250 1660 2290
rect 1660 2250 1670 2290
rect 1470 2230 1670 2250
rect 2080 2290 2280 2300
rect 2080 2250 2090 2290
rect 2090 2250 2270 2290
rect 2270 2250 2280 2290
rect 2080 2230 2280 2250
rect 2690 2290 2890 2300
rect 2690 2250 2700 2290
rect 2700 2250 2880 2290
rect 2880 2250 2890 2290
rect 2690 2230 2890 2250
rect -1310 1160 -1250 1230
rect -530 1160 -470 1230
rect -660 1060 -460 1080
rect -660 910 -650 1060
rect -650 910 -480 1060
rect -480 910 -460 1060
rect -660 890 -460 910
rect 1800 1950 1810 2010
rect 1810 1950 1870 2010
rect 1260 1500 1320 1560
rect 1660 1500 1720 1560
rect 190 1160 250 1230
rect 970 1160 1030 1230
rect 180 1060 380 1080
rect 180 910 200 1060
rect 200 910 370 1060
rect 370 910 380 1060
rect 180 890 380 910
rect -560 740 -500 810
rect 220 740 280 810
rect -1190 -20 -710 360
rect -380 -20 100 360
rect 1080 1280 1140 1300
rect 1080 1110 1120 1280
rect 1120 1110 1140 1280
rect 1080 1090 1140 1110
rect 430 -20 910 360
rect 1780 1450 1890 1610
rect 2490 1950 2550 2010
rect 2550 1950 2560 2010
rect 1950 1500 2010 1560
rect 2350 1500 2410 1560
rect 1390 -20 1590 360
rect 2470 1450 2580 1610
rect 2640 1500 2700 1560
rect 3040 1500 3100 1560
rect 2080 -20 2280 360
rect 2770 -20 2970 360
<< metal2 >>
rect 60 5500 160 5600
rect 470 5500 570 5600
rect 880 5500 980 5600
rect 1420 5500 1520 5600
rect 1770 5500 1870 5600
rect 2030 5500 2130 5600
rect 3210 5500 3310 5600
rect 3370 5500 3470 5600
rect 3530 5500 3630 5600
rect 3690 5500 3790 5600
rect 3850 5500 3950 5600
rect 4010 5500 4110 5600
rect -1310 5380 -1190 5390
rect -1310 5280 -1300 5380
rect -1200 5280 -1190 5380
rect -1310 5270 -1190 5280
rect -1010 5380 -890 5390
rect -1010 5280 -1000 5380
rect -900 5280 -890 5380
rect -1010 5270 -890 5280
rect 70 5170 150 5500
rect 70 5110 80 5170
rect 140 5110 150 5170
rect 70 4940 150 5110
rect 70 4880 80 4940
rect 140 4880 150 4940
rect 70 4870 150 4880
rect 480 5170 560 5500
rect 480 5110 490 5170
rect 550 5110 560 5170
rect 480 4940 560 5110
rect 480 4880 490 4940
rect 550 4880 560 4940
rect 890 5180 970 5500
rect 1230 5390 1400 5400
rect 1230 5240 1240 5390
rect 1390 5240 1400 5390
rect 1230 5230 1400 5240
rect 890 5120 900 5180
rect 960 5120 970 5180
rect 890 4950 970 5120
rect 890 4890 900 4950
rect 960 4890 970 4950
rect 890 4880 970 4890
rect 480 4870 560 4880
rect -530 4600 -410 4610
rect -530 4500 -520 4600
rect -420 4500 -410 4600
rect -530 4490 -410 4500
rect 1430 4290 1510 5500
rect 1550 5390 1750 5400
rect 1550 5170 1560 5390
rect 1740 5170 1750 5390
rect 1550 5160 1750 5170
rect 1780 4700 1860 5500
rect 2040 4850 2120 5500
rect 2160 5390 2360 5400
rect 2160 5170 2170 5390
rect 2350 5170 2360 5390
rect 2160 5160 2360 5170
rect 2770 5390 2970 5400
rect 2770 5170 2780 5390
rect 2960 5170 2970 5390
rect 2770 5160 2970 5170
rect 2040 4770 2740 4850
rect 1780 4620 2120 4700
rect 1430 4280 1860 4290
rect 1430 4220 1450 4280
rect 1510 4220 1790 4280
rect 1850 4220 1860 4280
rect 1430 4210 1860 4220
rect 2040 4220 2120 4620
rect 2660 4290 2740 4770
rect 2660 4280 3080 4290
rect 2660 4220 2670 4280
rect 2730 4220 3010 4280
rect 3070 4220 3080 4280
rect 2040 4210 2450 4220
rect 2660 4210 3080 4220
rect 1900 4170 2020 4180
rect -646 4020 -640 4140
rect -520 4020 -514 4140
rect 1900 4070 1910 4170
rect 2010 4070 2020 4170
rect 2050 4150 2080 4210
rect 2140 4150 2380 4210
rect 2440 4150 2450 4210
rect 2050 4140 2450 4150
rect 2500 4170 2620 4180
rect 210 4030 320 4040
rect -1500 3530 -1400 3540
rect -1500 3450 -1490 3530
rect -1410 3450 -1400 3530
rect -1500 3440 -1400 3450
rect -640 3530 -520 4020
rect -640 3400 -630 3530
rect -530 3400 -520 3530
rect 210 3940 220 4030
rect 310 3940 320 4030
rect 210 3590 320 3940
rect 210 3500 220 3590
rect 310 3500 320 3590
rect 210 3490 320 3500
rect 720 4030 830 4040
rect 720 3940 730 4030
rect 820 3940 830 4030
rect 720 3590 830 3940
rect 720 3500 730 3590
rect 820 3500 830 3590
rect 720 3490 830 3500
rect 1200 3990 1310 4000
rect 1200 3900 1210 3990
rect 1300 3900 1310 3990
rect -640 3390 -520 3400
rect 1200 3470 1310 3900
rect 1380 3950 1500 3960
rect 1380 3850 1390 3950
rect 1490 3850 1500 3950
rect 1380 3580 1500 3850
rect 1380 3500 1400 3580
rect 1480 3500 1500 3580
rect 1380 3480 1500 3500
rect 1900 3590 2020 4070
rect 1900 3490 1910 3590
rect 2010 3490 2020 3590
rect 1900 3480 2020 3490
rect 2500 4070 2510 4170
rect 2610 4070 2620 4170
rect 2500 3590 2620 4070
rect 3020 3950 3160 3960
rect 3020 3850 3030 3950
rect 3130 3850 3160 3950
rect 3020 3840 3160 3850
rect 2500 3490 2510 3590
rect 2610 3490 2620 3590
rect 2500 3480 2620 3490
rect 3040 3580 3160 3840
rect 3040 3500 3060 3580
rect 3140 3500 3160 3580
rect 3040 3480 3160 3500
rect 1200 3380 1210 3470
rect 1300 3380 1310 3470
rect 1200 3370 1310 3380
rect -1310 3010 -1210 3020
rect -1310 2930 -1300 3010
rect -1220 2930 -1210 3010
rect -1310 2920 -1210 2930
rect -1130 3010 -610 3020
rect -1130 2630 -1120 3010
rect -620 2630 -610 3010
rect -1130 2300 -610 2630
rect -1130 2230 -1120 2300
rect -620 2230 -610 2300
rect -1130 2220 -610 2230
rect -400 3010 120 3020
rect -400 2630 -390 3010
rect 110 2630 120 3010
rect -400 1850 120 2630
rect 330 3010 850 3020
rect 330 2630 340 3010
rect 840 2630 850 3010
rect 2040 3010 2480 3020
rect 330 2300 850 2630
rect 330 2230 340 2300
rect 840 2230 850 2300
rect 330 2220 850 2230
rect 1460 2750 1680 2760
rect 1460 2630 1470 2750
rect 1670 2630 1680 2750
rect 1460 2320 1680 2630
rect 2040 2630 2050 3010
rect 2470 2630 2480 3010
rect 2040 2620 2480 2630
rect 2680 2750 2900 2760
rect 2680 2630 2690 2750
rect 2890 2630 2900 2750
rect 2070 2320 2290 2620
rect 2680 2320 2900 2630
rect 1460 2300 2900 2320
rect 1460 2230 1470 2300
rect 1670 2230 2080 2300
rect 2280 2230 2690 2300
rect 2890 2230 2900 2300
rect 1460 2220 2900 2230
rect -400 1780 -390 1850
rect 110 1780 120 1850
rect -400 1770 120 1780
rect 1790 2010 1880 2220
rect 1790 1950 1800 2010
rect 1870 1950 1880 2010
rect 1790 1630 1880 1950
rect 2480 2010 2570 2220
rect 2480 1950 2490 2010
rect 2560 1950 2570 2010
rect 2480 1630 2570 1950
rect 1750 1610 1920 1630
rect 1260 1560 1340 1570
rect 1320 1500 1340 1560
rect -1430 1310 -1350 1320
rect -1430 1080 -1420 1310
rect -1360 1080 -1350 1310
rect 1070 1300 1150 1310
rect -1430 1070 -1350 1080
rect -1320 1230 -460 1240
rect -1320 1160 -1310 1230
rect -1250 1160 -530 1230
rect -470 1160 -460 1230
rect 180 1230 1040 1240
rect 180 1160 190 1230
rect 250 1160 970 1230
rect 1030 1160 1040 1230
rect -1320 1150 -460 1160
rect -1320 580 -1240 1150
rect -680 1080 -450 1090
rect -680 890 -660 1080
rect -460 890 -450 1080
rect -680 880 -450 890
rect 170 1080 400 1090
rect 170 890 180 1080
rect 380 890 400 1080
rect 960 1050 1040 1160
rect 1070 1090 1080 1300
rect 1140 1090 1150 1300
rect 1260 1230 1340 1500
rect 1640 1560 1720 1570
rect 1640 1500 1660 1560
rect 1640 1230 1720 1500
rect 1750 1450 1780 1610
rect 1890 1450 1920 1610
rect 2440 1610 2610 1630
rect 1750 1430 1920 1450
rect 1950 1560 2030 1570
rect 2010 1500 2030 1560
rect 1950 1380 2030 1500
rect 2330 1560 2410 1570
rect 2330 1500 2350 1560
rect 2330 1380 2410 1500
rect 2440 1450 2470 1610
rect 2580 1450 2610 1610
rect 3220 1570 3300 5500
rect 2640 1560 3300 1570
rect 2700 1500 3040 1560
rect 3100 1500 3300 1560
rect 2640 1490 3300 1500
rect 2440 1430 2610 1450
rect 3380 1380 3460 5500
rect 1950 1300 3460 1380
rect 3540 1230 3620 5500
rect 1260 1150 3620 1230
rect 1070 1080 1150 1090
rect 3700 1050 3780 5500
rect 960 970 3780 1050
rect 170 880 400 890
rect 3860 820 3940 5500
rect -570 810 3940 820
rect -570 740 -560 810
rect -500 740 220 810
rect 280 740 3940 810
rect -570 730 290 740
rect 4020 580 4100 5500
rect -1320 500 4100 580
rect -1210 360 -690 380
rect -1210 -20 -1190 360
rect -710 -20 -690 360
rect -1210 -40 -690 -20
rect -400 360 120 380
rect -400 -20 -380 360
rect 100 -20 120 360
rect -400 -40 120 -20
rect 410 360 930 380
rect 410 -20 430 360
rect 910 -20 930 360
rect 410 -40 930 -20
rect 1370 360 1610 380
rect 1370 -20 1390 360
rect 1590 -20 1610 360
rect 1370 -40 1610 -20
rect 2060 360 2300 380
rect 2060 -20 2080 360
rect 2280 -20 2300 360
rect 2060 -40 2300 -20
rect 2750 360 2990 380
rect 2750 -20 2770 360
rect 2970 -20 2990 360
rect 2750 -40 2990 -20
<< via2 >>
rect -1295 5285 -1205 5375
rect -995 5285 -905 5375
rect 1240 5240 1390 5390
rect -515 4505 -425 4595
rect 1560 5170 1740 5390
rect 2170 5170 2350 5390
rect 2780 5170 2960 5390
rect -1490 3450 -1410 3530
rect -630 3400 -530 3530
rect -1300 2930 -1220 3010
rect -1120 2630 -620 3010
rect -390 2630 110 3010
rect 340 2830 430 3010
rect 430 2830 610 3010
rect 610 2830 840 3010
rect 340 2630 840 2830
rect 1470 2630 1670 2750
rect 2050 2630 2470 3010
rect 2690 2630 2890 2750
rect -1420 1080 -1360 1310
rect -660 900 -470 1070
rect 190 900 380 1070
rect 1080 1090 1140 1300
rect -1190 -20 -710 360
rect -380 -20 100 360
rect 430 -20 910 360
rect 1390 -20 1590 360
rect 2080 -20 2280 360
rect 2770 -20 2970 360
<< metal3 >>
rect -1300 5390 -1200 5600
rect -1000 5390 -900 5600
rect -700 5410 -600 5600
rect -1310 5375 -1190 5390
rect -1310 5285 -1295 5375
rect -1205 5285 -1190 5375
rect -1310 5270 -1190 5285
rect -1010 5375 -890 5390
rect -1010 5285 -995 5375
rect -905 5285 -890 5375
rect -700 5310 -420 5410
rect -1010 5270 -890 5285
rect -520 4610 -420 5310
rect 1230 5390 4160 5400
rect 1230 5240 1240 5390
rect 1390 5240 1560 5390
rect 1230 5170 1560 5240
rect 1740 5170 2170 5390
rect 2350 5170 2780 5390
rect 2960 5170 4160 5390
rect 1230 5160 4160 5170
rect -530 4595 -410 4610
rect -530 4505 -515 4595
rect -425 4505 -410 4595
rect -530 4490 -410 4505
rect -1500 3530 -1400 3540
rect -1500 3450 -1490 3530
rect -1410 3450 -1400 3530
rect -1500 3440 -1400 3450
rect -640 3530 -520 3540
rect -640 3400 -630 3530
rect -530 3400 -520 3530
rect -640 3390 -520 3400
rect -1310 3010 -1210 3020
rect -1310 2930 -1300 3010
rect -1220 2930 -1210 3010
rect -1310 2920 -1210 2930
rect -1130 3010 -610 3020
rect -1430 2820 -1310 2840
rect -1430 2640 -1410 2820
rect -1330 2640 -1310 2820
rect -1430 1310 -1310 2640
rect -1130 2630 -1120 3010
rect -620 2630 -610 3010
rect -1130 2620 -610 2630
rect -400 3010 120 3020
rect -400 2630 -390 3010
rect 110 2630 120 3010
rect -400 2620 120 2630
rect 330 3010 850 3020
rect 330 2630 340 3010
rect 840 2630 850 3010
rect 2040 3010 2480 3020
rect 330 2620 850 2630
rect 1030 2820 1150 2840
rect 1030 2640 1050 2820
rect 1130 2640 1150 2820
rect -1430 1080 -1420 1310
rect -1360 1080 -1310 1310
rect 1030 1300 1150 2640
rect 1460 2750 1680 2760
rect 1460 2630 1470 2750
rect 1670 2630 1680 2750
rect 1460 2620 1680 2630
rect 2040 2630 2050 3010
rect 2470 2630 2480 3010
rect 2040 2620 2480 2630
rect 2680 2750 2900 2760
rect 2680 2630 2690 2750
rect 2890 2630 2900 2750
rect 2680 2620 2900 2630
rect 1030 1090 1080 1300
rect 1140 1090 1150 1300
rect -1430 1000 -1310 1080
rect -680 1070 -450 1090
rect -680 1000 -660 1070
rect -1430 900 -660 1000
rect -470 1000 -450 1070
rect 170 1070 400 1090
rect 170 1000 190 1070
rect -470 900 190 1000
rect 380 1000 400 1070
rect 1030 1000 1150 1090
rect 380 900 1150 1000
rect -1430 880 1150 900
rect 3920 380 4160 5160
rect -1280 360 4160 380
rect -1280 -20 -1190 360
rect -710 -20 -380 360
rect 100 -20 430 360
rect 910 -20 1390 360
rect 1590 -20 2080 360
rect 2280 -20 2770 360
rect 2970 -20 4160 360
rect -1280 -40 4160 -20
rect 3480 -360 4160 -40
<< via3 >>
rect -1490 3450 -1410 3530
rect -630 3400 -530 3530
rect -1300 2930 -1220 3010
rect -1410 2640 -1330 2820
rect -1120 2630 -620 3010
rect -390 2630 110 3010
rect 340 2630 840 3010
rect 1050 2640 1130 2820
rect 1470 2630 1670 2750
rect 2050 2630 2470 3010
rect 2690 2630 2890 2750
<< metal4 >>
rect -1900 3530 -460 3540
rect -1900 3450 -1490 3530
rect -1410 3450 -630 3530
rect -1900 3400 -630 3450
rect -530 3400 -460 3530
rect -1900 3140 -460 3400
rect -1900 3010 2980 3020
rect -1900 2930 -1300 3010
rect -1220 2930 -1120 3010
rect -1900 2820 -1120 2930
rect -1900 2640 -1410 2820
rect -1330 2640 -1120 2820
rect -1900 2630 -1120 2640
rect -620 2630 -390 3010
rect 110 2630 340 3010
rect 840 2820 2050 3010
rect 840 2640 1050 2820
rect 1130 2750 2050 2820
rect 1130 2640 1470 2750
rect 840 2630 1470 2640
rect 1670 2630 2050 2750
rect 2470 2750 2980 3010
rect 2470 2630 2690 2750
rect 2890 2630 2980 2750
rect -1900 2620 2980 2630
use sky130_fd_pr__pfet_01v8_JE7DK3  XM1 segdac__devices
timestamp 1725599052
transform 1 0 -1254 0 1 4929
box -246 -269 246 269
use sky130_fd_pr__pfet_01v8_QBPJZQ  XM2 segdac__devices
timestamp 1725599052
transform 1 0 -724 0 1 4929
box -296 -269 296 269
use sky130_fd_pr__pfet_01v8_8JDY5S  XM3 segdac__devices
timestamp 1725599052
transform 1 0 -914 0 1 4409
box -396 -269 396 269
use sky130_fd_pr__nfet_01v8_DB7J7C  XMia1 segdac__devices
timestamp 1725599052
transform 0 1 10 -1 0 4076
box -696 -260 696 260
use sky130_fd_pr__nfet_01v8_DB7J7C  XMia2
timestamp 1725599052
transform 0 1 520 -1 0 4076
box -696 -260 696 260
use sky130_fd_pr__nfet_01v8_DB7J7C  XMia3
timestamp 1725599052
transform 0 1 1030 -1 0 4076
box -696 -260 696 260
use sky130_fd_pr__nfet_01v8_33M553  XMib1 segdac__devices
timestamp 1725599052
transform 1 0 1696 0 1 3540
box -316 -260 316 260
use sky130_fd_pr__nfet_01v8_33M553  XMib2
timestamp 1725599052
transform 0 1 2260 -1 0 3716
box -316 -260 316 260
use sky130_fd_pr__nfet_01v8_33M553  XMib3
timestamp 1725599052
transform 1 0 2836 0 1 3540
box -316 -260 316 260
use sky130_fd_pr__nfet_01v8_7DN82Q  XMic1 segdac__devices
timestamp 1725599052
transform 0 1 2790 -1 0 2076
box -246 -310 246 310
use sky130_fd_pr__nfet_01v8_7DN82Q  XMic2
timestamp 1725599052
transform 0 1 2180 -1 0 2076
box -246 -310 246 310
use sky130_fd_pr__nfet_01v8_7DN82Q  XMic3
timestamp 1725599052
transform 0 1 1570 -1 0 2076
box -246 -310 246 310
use sky130_fd_pr__nfet_01v8_3ZUKNL  XMid1 segdac__devices
timestamp 1725599052
transform 0 1 590 -1 0 2086
box -226 -470 226 470
use sky130_fd_pr__nfet_01v8_3ZUKNL  XMid2
timestamp 1725599052
transform 0 1 -140 -1 0 1636
box -226 -470 226 470
use sky130_fd_pr__nfet_01v8_3ZUKNL  XMid3
timestamp 1725599052
transform 0 1 -870 -1 0 2086
box -226 -470 226 470
use sky130_fd_pr__nfet_01v8_VRHU84  XMmirror segdac__devices
timestamp 1725599052
transform 1 0 -1064 0 1 3830
box -246 -260 246 260
use sky130_fd_pr__nfet_01v8_AJ3M4R  XMsa1 segdac__devices
timestamp 1725599052
transform 1 0 111 0 1 5020
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_AJ3M4R  XMsa2
timestamp 1725599052
transform 1 0 521 0 1 5020
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_AJ3M4R  XMsa3
timestamp 1725599052
transform 1 0 931 0 1 5030
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_V8CAV6  XMsb1 segdac__devices
timestamp 1725599052
transform 0 1 1650 -1 0 4161
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_V8CAV6  XMsb2
timestamp 1725599052
transform 0 1 2260 -1 0 4331
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_V8CAV6  XMsb3
timestamp 1725599052
transform 0 1 2870 -1 0 4161
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_V8CYR7  XMsc1 segdac__devices
timestamp 1725599052
transform 0 1 2870 -1 0 1531
box -211 -350 211 350
use sky130_fd_pr__nfet_01v8_V8CYR7  XMsc2
timestamp 1725599052
transform 0 1 2180 -1 0 1531
box -211 -350 211 350
use sky130_fd_pr__nfet_01v8_V8CYR7  XMsc3
timestamp 1725599052
transform 0 1 1490 -1 0 1531
box -211 -350 211 350
use sky130_fd_pr__nfet_01v8_2BSVCH  XMsd1 segdac__devices
timestamp 1725599052
transform 0 1 610 -1 0 1196
box -216 -540 216 540
use sky130_fd_pr__nfet_01v8_2BSVCH  XMsd2
timestamp 1725599052
transform 0 1 -140 -1 0 776
box -216 -540 216 540
use sky130_fd_pr__nfet_01v8_2BSVCH  XMsd3
timestamp 1725599052
transform 0 1 -890 -1 0 1196
box -216 -540 216 540
<< labels >>
flabel metal3 -1300 5500 -1200 5600 0 FreeSans 480 0 0 0 bias1
port 21 nsew
flabel metal3 -1000 5500 -900 5600 0 FreeSans 480 0 0 0 bias2
port 22 nsew
flabel metal3 -700 5500 -600 5600 0 FreeSans 480 0 0 0 bias3
port 24 nsew
flabel metal2 60 5500 160 5600 0 FreeSans 480 0 0 0 sa1
port 25 nsew
flabel metal2 470 5500 570 5600 0 FreeSans 480 0 0 0 sa2
port 26 nsew
flabel metal2 880 5500 980 5600 0 FreeSans 480 0 0 0 sa3
port 27 nsew
flabel metal2 1420 5500 1520 5600 0 FreeSans 480 0 0 0 sb1
port 30 nsew
flabel metal2 1770 5500 1870 5600 0 FreeSans 480 0 0 0 sb2
port 31 nsew
flabel metal2 2030 5500 2130 5600 0 FreeSans 480 0 0 0 sb3
port 32 nsew
flabel metal2 3210 5500 3310 5600 0 FreeSans 480 0 0 0 sc1
port 33 nsew
flabel metal2 3370 5500 3470 5600 0 FreeSans 480 0 0 0 sc2
port 34 nsew
flabel metal2 3530 5500 3630 5600 0 FreeSans 480 0 0 0 sc3
port 35 nsew
flabel metal2 3690 5500 3790 5600 0 FreeSans 480 0 0 0 sd1
port 36 nsew
flabel metal2 3850 5500 3950 5600 0 FreeSans 480 0 0 0 sd2
port 37 nsew
flabel metal2 4010 5500 4110 5600 0 FreeSans 480 0 0 0 sd3
port 38 nsew
flabel metal4 -1900 3140 -1500 3540 0 FreeSans 1600 0 0 0 vcc
port 19 nsew
flabel metal4 -1900 2620 -1500 3020 0 FreeSans 1600 0 0 0 vss
port 20 nsew
flabel metal1 -1901 2349 -1739 2511 0 FreeSans 480 0 0 0 Vbias
port 28 nsew
flabel metal3 3480 -360 4160 320 0 FreeSans 1600 0 0 0 Vout
port 29 nsew
<< end >>

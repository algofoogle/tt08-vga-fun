magic
tech sky130A
timestamp 1725599052
<< pwell >>
rect -158 -130 158 130
<< nmos >>
rect -60 -25 60 25
<< ndiff >>
rect -89 19 -60 25
rect -89 -19 -83 19
rect -66 -19 -60 19
rect -89 -25 -60 -19
rect 60 19 89 25
rect 60 -19 66 19
rect 83 -19 89 19
rect 60 -25 89 -19
<< ndiffc >>
rect -83 -19 -66 19
rect 66 -19 83 19
<< psubdiff >>
rect -140 95 -92 112
rect 92 95 140 112
rect -140 64 -123 95
rect 123 64 140 95
rect -140 -95 -123 -64
rect 123 -95 140 -64
rect -140 -112 -92 -95
rect 92 -112 140 -95
<< psubdiffcont >>
rect -92 95 92 112
rect -140 -64 -123 64
rect 123 -64 140 64
rect -92 -112 92 -95
<< poly >>
rect -60 61 60 69
rect -60 44 -52 61
rect 52 44 60 61
rect -60 25 60 44
rect -60 -44 60 -25
rect -60 -61 -52 -44
rect 52 -61 60 -44
rect -60 -69 60 -61
<< polycont >>
rect -52 44 52 61
rect -52 -61 52 -44
<< locali >>
rect -140 95 -92 112
rect 92 95 140 112
rect -140 64 -123 95
rect 123 64 140 95
rect -60 44 -52 61
rect 52 44 60 61
rect -83 19 -66 27
rect -83 -27 -66 -19
rect 66 19 83 27
rect 66 -27 83 -19
rect -60 -61 -52 -44
rect 52 -61 60 -44
rect -140 -95 -123 -64
rect 123 -95 140 -64
rect -140 -112 -92 -95
rect 92 -112 140 -95
<< viali >>
rect -52 44 52 61
rect -83 -19 -66 19
rect 66 -19 83 19
rect -52 -61 52 -44
<< metal1 >>
rect -58 61 58 64
rect -58 44 -52 61
rect 52 44 58 61
rect -58 41 58 44
rect -86 19 -63 25
rect -86 -19 -83 19
rect -66 -19 -63 19
rect -86 -25 -63 -19
rect 63 19 86 25
rect 63 -19 66 19
rect 83 -19 86 19
rect 63 -25 86 -19
rect -58 -44 58 -41
rect -58 -61 -52 -44
rect 52 -61 58 -44
rect -58 -64 58 -61
<< properties >>
string FIXED_BBOX -131 -103 131 103
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.5 l 1.2 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

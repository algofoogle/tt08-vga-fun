magic
tech sky130A
timestamp 1723780759
<< pwell >>
rect -123 -130 123 130
<< nmos >>
rect -25 -25 25 25
<< ndiff >>
rect -54 19 -25 25
rect -54 -19 -48 19
rect -31 -19 -25 19
rect -54 -25 -25 -19
rect 25 19 54 25
rect 25 -19 31 19
rect 48 -19 54 19
rect 25 -25 54 -19
<< ndiffc >>
rect -48 -19 -31 19
rect 31 -19 48 19
<< psubdiff >>
rect -105 95 -57 112
rect 57 95 105 112
rect -105 64 -88 95
rect 88 64 105 95
rect -105 -95 -88 -64
rect 88 -95 105 -64
rect -105 -112 -57 -95
rect 57 -112 105 -95
<< psubdiffcont >>
rect -57 95 57 112
rect -105 -64 -88 64
rect 88 -64 105 64
rect -57 -112 57 -95
<< poly >>
rect -25 61 25 69
rect -25 44 -17 61
rect 17 44 25 61
rect -25 25 25 44
rect -25 -44 25 -25
rect -25 -61 -17 -44
rect 17 -61 25 -44
rect -25 -69 25 -61
<< polycont >>
rect -17 44 17 61
rect -17 -61 17 -44
<< locali >>
rect -105 95 -57 112
rect 57 95 105 112
rect -105 64 -88 95
rect 88 64 105 95
rect -25 44 -17 61
rect 17 44 25 61
rect -48 19 -31 27
rect -48 -27 -31 -19
rect 31 19 48 27
rect 31 -27 48 -19
rect -25 -61 -17 -44
rect 17 -61 25 -44
rect -105 -95 -88 -64
rect 88 -95 105 -64
rect -105 -112 -57 -95
rect 57 -112 105 -95
<< viali >>
rect -17 44 17 61
rect -48 -19 -31 19
rect 31 -19 48 19
rect -17 -61 17 -44
<< metal1 >>
rect -23 61 23 64
rect -23 44 -17 61
rect 17 44 23 61
rect -23 41 23 44
rect -51 19 -28 25
rect -51 -19 -48 19
rect -31 -19 -28 19
rect -51 -25 -28 -19
rect 28 19 51 25
rect 28 -19 31 19
rect 48 -19 51 19
rect 28 -25 51 -19
rect -23 -44 23 -41
rect -23 -61 -17 -44
rect 17 -61 23 -44
rect -23 -64 23 -61
<< properties >>
string FIXED_BBOX -96 -103 96 103
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.5 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

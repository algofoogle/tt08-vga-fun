magic
tech sky130A
magscale 1 2
timestamp 1724295482
<< viali >>
rect 8125 23273 8159 23307
rect 10333 23273 10367 23307
rect 10609 23273 10643 23307
rect 11437 23273 11471 23307
rect 11805 23273 11839 23307
rect 13369 23273 13403 23307
rect 20085 23273 20119 23307
rect 16405 23205 16439 23239
rect 18337 23205 18371 23239
rect 18972 23205 19006 23239
rect 22937 23205 22971 23239
rect 2237 23137 2271 23171
rect 2421 23137 2455 23171
rect 3249 23137 3283 23171
rect 3505 23137 3539 23171
rect 4721 23137 4755 23171
rect 5825 23137 5859 23171
rect 6009 23137 6043 23171
rect 6736 23137 6770 23171
rect 7941 23137 7975 23171
rect 9698 23137 9732 23171
rect 10149 23137 10183 23171
rect 10793 23137 10827 23171
rect 10977 23137 11011 23171
rect 11253 23137 11287 23171
rect 11621 23137 11655 23171
rect 11989 23137 12023 23171
rect 12245 23137 12279 23171
rect 13737 23137 13771 23171
rect 15678 23137 15712 23171
rect 16845 23137 16879 23171
rect 20269 23137 20303 23171
rect 22405 23137 22439 23171
rect 4997 23069 5031 23103
rect 6469 23069 6503 23103
rect 9965 23069 9999 23103
rect 13829 23069 13863 23103
rect 15945 23069 15979 23103
rect 16589 23069 16623 23103
rect 18705 23069 18739 23103
rect 20545 23069 20579 23103
rect 22661 23069 22695 23103
rect 4813 23001 4847 23035
rect 11161 23001 11195 23035
rect 14565 23001 14599 23035
rect 16221 23001 16255 23035
rect 17969 23001 18003 23035
rect 2329 22933 2363 22967
rect 4629 22933 4663 22967
rect 4905 22933 4939 22967
rect 5917 22933 5951 22967
rect 7849 22933 7883 22967
rect 8585 22933 8619 22967
rect 13553 22933 13587 22967
rect 14473 22933 14507 22967
rect 18429 22933 18463 22967
rect 21281 22933 21315 22967
rect 22845 22933 22879 22967
rect 5549 22729 5583 22763
rect 5733 22729 5767 22763
rect 6653 22729 6687 22763
rect 9229 22729 9263 22763
rect 9505 22729 9539 22763
rect 9873 22729 9907 22763
rect 12081 22729 12115 22763
rect 8953 22661 8987 22695
rect 14381 22661 14415 22695
rect 18705 22661 18739 22695
rect 21557 22661 21591 22695
rect 1593 22593 1627 22627
rect 1961 22593 1995 22627
rect 2697 22593 2731 22627
rect 2973 22593 3007 22627
rect 3617 22593 3651 22627
rect 4445 22593 4479 22627
rect 7389 22593 7423 22627
rect 8125 22593 8159 22627
rect 8493 22593 8527 22627
rect 12817 22593 12851 22627
rect 14933 22593 14967 22627
rect 17601 22593 17635 22627
rect 19257 22593 19291 22627
rect 20085 22593 20119 22627
rect 1501 22525 1535 22559
rect 1685 22525 1719 22559
rect 1777 22525 1811 22559
rect 2145 22525 2179 22559
rect 2605 22525 2639 22559
rect 3525 22525 3559 22559
rect 3709 22525 3743 22559
rect 3985 22525 4019 22559
rect 4169 22525 4203 22559
rect 4721 22525 4755 22559
rect 5457 22525 5491 22559
rect 5641 22525 5675 22559
rect 5917 22525 5951 22559
rect 6377 22525 6411 22559
rect 6469 22525 6503 22559
rect 8585 22525 8619 22559
rect 9045 22525 9079 22559
rect 9321 22525 9355 22559
rect 9689 22525 9723 22559
rect 10057 22525 10091 22559
rect 11529 22525 11563 22559
rect 11713 22525 11747 22559
rect 11805 22525 11839 22559
rect 11989 22525 12023 22559
rect 12265 22525 12299 22559
rect 12541 22525 12575 22559
rect 12725 22525 12759 22559
rect 13001 22525 13035 22559
rect 13093 22525 13127 22559
rect 13553 22525 13587 22559
rect 13737 22525 13771 22559
rect 15117 22525 15151 22559
rect 15577 22525 15611 22559
rect 18429 22525 18463 22559
rect 19073 22525 19107 22559
rect 19165 22525 19199 22559
rect 20545 22525 20579 22559
rect 20913 22525 20947 22559
rect 21189 22525 21223 22559
rect 22937 22525 22971 22559
rect 1869 22457 1903 22491
rect 6101 22457 6135 22491
rect 7113 22457 7147 22491
rect 7573 22457 7607 22491
rect 10324 22457 10358 22491
rect 11621 22457 11655 22491
rect 13921 22457 13955 22491
rect 14013 22457 14047 22491
rect 15822 22457 15856 22491
rect 17417 22457 17451 22491
rect 17877 22457 17911 22491
rect 20637 22457 20671 22491
rect 20729 22457 20763 22491
rect 22692 22457 22726 22491
rect 3801 22389 3835 22423
rect 5365 22389 5399 22423
rect 6193 22389 6227 22423
rect 6745 22389 6779 22423
rect 7205 22389 7239 22423
rect 11437 22389 11471 22423
rect 11897 22389 11931 22423
rect 14473 22389 14507 22423
rect 15025 22389 15059 22423
rect 15485 22389 15519 22423
rect 16957 22389 16991 22423
rect 17049 22389 17083 22423
rect 17509 22389 17543 22423
rect 19533 22389 19567 22423
rect 19901 22389 19935 22423
rect 19993 22389 20027 22423
rect 20361 22389 20395 22423
rect 21097 22389 21131 22423
rect 1961 22185 1995 22219
rect 2605 22185 2639 22219
rect 2881 22185 2915 22219
rect 4813 22185 4847 22219
rect 7297 22185 7331 22219
rect 8309 22185 8343 22219
rect 9045 22185 9079 22219
rect 9321 22185 9355 22219
rect 10333 22185 10367 22219
rect 11713 22185 11747 22219
rect 15577 22185 15611 22219
rect 16313 22185 16347 22219
rect 17325 22185 17359 22219
rect 19165 22185 19199 22219
rect 20269 22185 20303 22219
rect 2329 22117 2363 22151
rect 3709 22117 3743 22151
rect 9965 22117 9999 22151
rect 10165 22117 10199 22151
rect 11253 22117 11287 22151
rect 13645 22117 13679 22151
rect 14657 22117 14691 22151
rect 14841 22117 14875 22151
rect 15025 22117 15059 22151
rect 20545 22117 20579 22151
rect 22937 22117 22971 22151
rect 1685 22049 1719 22083
rect 1869 22049 1903 22083
rect 2145 22049 2179 22083
rect 2421 22049 2455 22083
rect 2789 22049 2823 22083
rect 2973 22049 3007 22083
rect 3341 22049 3375 22083
rect 3617 22049 3651 22083
rect 3801 22049 3835 22083
rect 3893 22049 3927 22083
rect 4169 22049 4203 22083
rect 4353 22049 4387 22083
rect 4629 22049 4663 22083
rect 5089 22049 5123 22083
rect 5273 22049 5307 22083
rect 5457 22049 5491 22083
rect 5549 22049 5583 22083
rect 6009 22049 6043 22083
rect 7113 22049 7147 22083
rect 7665 22049 7699 22083
rect 7941 22049 7975 22083
rect 8217 22049 8251 22083
rect 8401 22049 8435 22083
rect 10609 22049 10643 22083
rect 10793 22049 10827 22083
rect 11437 22049 11471 22083
rect 11897 22049 11931 22083
rect 11989 22049 12023 22083
rect 12173 22049 12207 22083
rect 12909 22049 12943 22083
rect 13553 22049 13587 22083
rect 13829 22049 13863 22083
rect 13921 22049 13955 22083
rect 14197 22049 14231 22083
rect 15117 22049 15151 22083
rect 15393 22049 15427 22083
rect 15669 22049 15703 22083
rect 16129 22049 16163 22083
rect 16865 22049 16899 22083
rect 18449 22049 18483 22083
rect 18705 22049 18739 22083
rect 19809 22049 19843 22083
rect 19901 22049 19935 22083
rect 19993 22049 20027 22083
rect 20177 22049 20211 22083
rect 20453 22049 20487 22083
rect 20637 22049 20671 22083
rect 20821 22049 20855 22083
rect 21097 22049 21131 22083
rect 21548 22049 21582 22083
rect 3065 21981 3099 22015
rect 4445 21981 4479 22015
rect 6101 21981 6135 22015
rect 6837 21981 6871 22015
rect 9505 21981 9539 22015
rect 9597 21981 9631 22015
rect 9689 21981 9723 22015
rect 9781 21981 9815 22015
rect 14289 21981 14323 22015
rect 16957 21981 16991 22015
rect 17141 21981 17175 22015
rect 18981 21981 19015 22015
rect 19073 21981 19107 22015
rect 21281 21981 21315 22015
rect 3157 21913 3191 21947
rect 4537 21913 4571 21947
rect 5365 21913 5399 21947
rect 6929 21913 6963 21947
rect 7389 21913 7423 21947
rect 8033 21913 8067 21947
rect 8585 21913 8619 21947
rect 8677 21913 8711 21947
rect 9229 21913 9263 21947
rect 11069 21913 11103 21947
rect 13093 21913 13127 21947
rect 13369 21913 13403 21947
rect 15301 21913 15335 21947
rect 19625 21913 19659 21947
rect 22661 21913 22695 21947
rect 1869 21845 1903 21879
rect 3249 21845 3283 21879
rect 4077 21845 4111 21879
rect 4905 21845 4939 21879
rect 6377 21845 6411 21879
rect 7573 21845 7607 21879
rect 9045 21845 9079 21879
rect 10149 21845 10183 21879
rect 10425 21845 10459 21879
rect 12081 21845 12115 21879
rect 12541 21845 12575 21879
rect 13645 21845 13679 21879
rect 14565 21845 14599 21879
rect 15853 21845 15887 21879
rect 16497 21845 16531 21879
rect 19533 21845 19567 21879
rect 20913 21845 20947 21879
rect 22845 21845 22879 21879
rect 2881 21641 2915 21675
rect 3433 21641 3467 21675
rect 5917 21641 5951 21675
rect 6377 21641 6411 21675
rect 7481 21641 7515 21675
rect 9045 21641 9079 21675
rect 10149 21641 10183 21675
rect 14013 21641 14047 21675
rect 14841 21641 14875 21675
rect 18153 21641 18187 21675
rect 19901 21641 19935 21675
rect 20545 21641 20579 21675
rect 4353 21573 4387 21607
rect 7205 21573 7239 21607
rect 8769 21573 8803 21607
rect 9505 21573 9539 21607
rect 10885 21573 10919 21607
rect 13369 21573 13403 21607
rect 21373 21573 21407 21607
rect 2237 21505 2271 21539
rect 2789 21505 2823 21539
rect 2973 21505 3007 21539
rect 3709 21505 3743 21539
rect 4077 21505 4111 21539
rect 6791 21505 6825 21539
rect 12541 21505 12575 21539
rect 16773 21505 16807 21539
rect 19165 21505 19199 21539
rect 22753 21505 22787 21539
rect 1970 21437 2004 21471
rect 2513 21437 2547 21471
rect 3065 21437 3099 21471
rect 3893 21437 3927 21471
rect 4537 21437 4571 21471
rect 4721 21437 4755 21471
rect 5181 21437 5215 21471
rect 5457 21437 5491 21471
rect 5825 21437 5859 21471
rect 6101 21437 6135 21471
rect 6193 21437 6227 21471
rect 6653 21437 6687 21471
rect 6929 21437 6963 21471
rect 7021 21437 7055 21471
rect 7113 21437 7147 21471
rect 7389 21437 7423 21471
rect 7481 21437 7515 21471
rect 7665 21437 7699 21471
rect 8585 21437 8619 21471
rect 8677 21437 8711 21471
rect 9229 21437 9263 21471
rect 9321 21437 9355 21471
rect 9781 21437 9815 21471
rect 10057 21437 10091 21471
rect 10241 21437 10275 21471
rect 10609 21437 10643 21471
rect 11069 21437 11103 21471
rect 11621 21437 11655 21471
rect 11897 21437 11931 21471
rect 12449 21437 12483 21471
rect 13185 21437 13219 21471
rect 13737 21437 13771 21471
rect 14197 21437 14231 21471
rect 14289 21437 14323 21471
rect 14381 21437 14415 21471
rect 14473 21437 14507 21471
rect 14657 21437 14691 21471
rect 14841 21437 14875 21471
rect 16681 21437 16715 21471
rect 17029 21437 17063 21471
rect 18337 21437 18371 21471
rect 20085 21437 20119 21471
rect 20177 21437 20211 21471
rect 20269 21437 20303 21471
rect 20453 21437 20487 21471
rect 20729 21437 20763 21471
rect 20913 21437 20947 21471
rect 21097 21437 21131 21471
rect 23029 21437 23063 21471
rect 3401 21369 3435 21403
rect 3617 21369 3651 21403
rect 14933 21369 14967 21403
rect 18797 21369 18831 21403
rect 19349 21369 19383 21403
rect 20821 21369 20855 21403
rect 22486 21369 22520 21403
rect 857 21301 891 21335
rect 2697 21301 2731 21335
rect 3249 21301 3283 21335
rect 4629 21301 4663 21335
rect 4905 21301 4939 21335
rect 5089 21301 5123 21335
rect 5641 21301 5675 21335
rect 8401 21301 8435 21335
rect 9965 21301 9999 21335
rect 10701 21301 10735 21335
rect 11437 21301 11471 21335
rect 11713 21301 11747 21335
rect 12817 21301 12851 21335
rect 13921 21301 13955 21335
rect 18429 21301 18463 21335
rect 18889 21301 18923 21335
rect 19441 21301 19475 21335
rect 19809 21301 19843 21335
rect 22845 21301 22879 21335
rect 2513 21097 2547 21131
rect 3801 21097 3835 21131
rect 5365 21097 5399 21131
rect 5641 21097 5675 21131
rect 6285 21097 6319 21131
rect 7113 21097 7147 21131
rect 7849 21097 7883 21131
rect 8585 21097 8619 21131
rect 12173 21097 12207 21131
rect 15209 21097 15243 21131
rect 15945 21097 15979 21131
rect 20545 21097 20579 21131
rect 21649 21097 21683 21131
rect 1685 21029 1719 21063
rect 2145 21029 2179 21063
rect 2345 21029 2379 21063
rect 2973 21029 3007 21063
rect 8468 21029 8502 21063
rect 9137 21029 9171 21063
rect 15485 21029 15519 21063
rect 15669 21029 15703 21063
rect 20821 21029 20855 21063
rect 20913 21029 20947 21063
rect 21465 21029 21499 21063
rect 1593 20961 1627 20995
rect 1777 20961 1811 20995
rect 1869 20961 1903 20995
rect 2789 20961 2823 20995
rect 3341 20961 3375 20995
rect 3985 20961 4019 20995
rect 4261 20961 4295 20995
rect 4445 20961 4479 20995
rect 4537 20961 4571 20995
rect 4629 20961 4663 20995
rect 4721 20961 4755 20995
rect 4997 20961 5031 20995
rect 5273 20961 5307 20995
rect 5457 20961 5491 20995
rect 5825 20961 5859 20995
rect 6101 20961 6135 20995
rect 6469 20961 6503 20995
rect 6561 20961 6595 20995
rect 7205 20961 7239 20995
rect 7665 20961 7699 20995
rect 7941 20961 7975 20995
rect 8125 20961 8159 20995
rect 9045 20961 9079 20995
rect 9873 20961 9907 20995
rect 10977 20961 11011 20995
rect 11161 20961 11195 20995
rect 11253 20961 11287 20995
rect 11345 20961 11379 20995
rect 11989 20961 12023 20995
rect 12081 20961 12115 20995
rect 13286 20961 13320 20995
rect 13553 20961 13587 20995
rect 13829 20961 13863 20995
rect 14473 20961 14507 20995
rect 14841 20961 14875 20995
rect 15761 20961 15795 20995
rect 16396 20961 16430 20995
rect 18705 20961 18739 20995
rect 20729 20961 20763 20995
rect 21097 20961 21131 20995
rect 22762 20961 22796 20995
rect 23029 20961 23063 20995
rect 6837 20893 6871 20927
rect 7389 20893 7423 20927
rect 7481 20893 7515 20927
rect 8033 20893 8067 20927
rect 8677 20893 8711 20927
rect 8953 20893 8987 20927
rect 9689 20893 9723 20927
rect 9781 20893 9815 20927
rect 9965 20893 9999 20927
rect 13921 20893 13955 20927
rect 14197 20893 14231 20927
rect 14749 20893 14783 20927
rect 16129 20893 16163 20927
rect 17601 20893 17635 20927
rect 17877 20893 17911 20927
rect 20453 20893 20487 20927
rect 2053 20825 2087 20859
rect 3157 20825 3191 20859
rect 5089 20825 5123 20859
rect 7573 20825 7607 20859
rect 8309 20825 8343 20859
rect 11621 20825 11655 20859
rect 17509 20825 17543 20859
rect 2329 20757 2363 20791
rect 2605 20757 2639 20791
rect 4077 20757 4111 20791
rect 6101 20757 6135 20791
rect 6837 20757 6871 20791
rect 9505 20757 9539 20791
rect 11713 20757 11747 20791
rect 11989 20757 12023 20791
rect 14289 20757 14323 20791
rect 15301 20757 15335 20791
rect 21373 20757 21407 20791
rect 6377 20553 6411 20587
rect 6837 20553 6871 20587
rect 7205 20553 7239 20587
rect 7941 20553 7975 20587
rect 10609 20553 10643 20587
rect 10793 20553 10827 20587
rect 11437 20553 11471 20587
rect 13185 20553 13219 20587
rect 13553 20553 13587 20587
rect 14289 20553 14323 20587
rect 14565 20553 14599 20587
rect 14749 20553 14783 20587
rect 15761 20553 15795 20587
rect 16589 20553 16623 20587
rect 20177 20553 20211 20587
rect 21741 20553 21775 20587
rect 22661 20553 22695 20587
rect 7573 20485 7607 20519
rect 8953 20485 8987 20519
rect 17141 20485 17175 20519
rect 20821 20485 20855 20519
rect 21465 20485 21499 20519
rect 3249 20417 3283 20451
rect 7665 20417 7699 20451
rect 9413 20417 9447 20451
rect 11805 20417 11839 20451
rect 13921 20417 13955 20451
rect 15117 20417 15151 20451
rect 16221 20417 16255 20451
rect 16405 20417 16439 20451
rect 16957 20417 16991 20451
rect 19349 20417 19383 20451
rect 1593 20349 1627 20383
rect 1869 20349 1903 20383
rect 2053 20349 2087 20383
rect 2513 20349 2547 20383
rect 2697 20349 2731 20383
rect 6929 20349 6963 20383
rect 7389 20349 7423 20383
rect 7941 20349 7975 20383
rect 8033 20349 8067 20383
rect 8217 20349 8251 20383
rect 8585 20349 8619 20383
rect 8769 20349 8803 20383
rect 9597 20349 9631 20383
rect 9689 20349 9723 20383
rect 9965 20349 9999 20383
rect 10077 20349 10111 20383
rect 10241 20349 10275 20383
rect 10333 20349 10367 20383
rect 10425 20349 10459 20383
rect 10977 20349 11011 20383
rect 11069 20349 11103 20383
rect 13737 20349 13771 20383
rect 14105 20349 14139 20383
rect 14381 20349 14415 20383
rect 14657 20349 14691 20383
rect 14841 20349 14875 20383
rect 15301 20349 15335 20383
rect 15485 20349 15519 20383
rect 16129 20349 16163 20383
rect 16773 20349 16807 20383
rect 16865 20349 16899 20383
rect 18521 20349 18555 20383
rect 20361 20349 20395 20383
rect 20729 20349 20763 20383
rect 21005 20349 21039 20383
rect 21097 20349 21131 20383
rect 21373 20349 21407 20383
rect 21741 20349 21775 20383
rect 21925 20349 21959 20383
rect 22201 20349 22235 20383
rect 22385 20349 22419 20383
rect 1777 20281 1811 20315
rect 3494 20281 3528 20315
rect 4905 20281 4939 20315
rect 9137 20281 9171 20315
rect 9321 20281 9355 20315
rect 12072 20281 12106 20315
rect 18276 20281 18310 20315
rect 18705 20281 18739 20315
rect 18889 20281 18923 20315
rect 20453 20281 20487 20315
rect 20545 20281 20579 20315
rect 21189 20281 21223 20315
rect 22477 20281 22511 20315
rect 22693 20281 22727 20315
rect 1409 20213 1443 20247
rect 1961 20213 1995 20247
rect 2697 20213 2731 20247
rect 4629 20213 4663 20247
rect 7757 20213 7791 20247
rect 8585 20213 8619 20247
rect 9781 20213 9815 20247
rect 11437 20213 11471 20247
rect 11621 20213 11655 20247
rect 19073 20213 19107 20247
rect 19441 20213 19475 20247
rect 19533 20213 19567 20247
rect 19901 20213 19935 20247
rect 22017 20213 22051 20247
rect 22845 20213 22879 20247
rect 1777 20009 1811 20043
rect 2805 20009 2839 20043
rect 4629 20009 4663 20043
rect 5089 20009 5123 20043
rect 5825 20009 5859 20043
rect 6193 20009 6227 20043
rect 6285 20009 6319 20043
rect 6653 20009 6687 20043
rect 10333 20009 10367 20043
rect 11437 20009 11471 20043
rect 11529 20009 11563 20043
rect 13645 20009 13679 20043
rect 15209 20009 15243 20043
rect 15945 20009 15979 20043
rect 16615 20009 16649 20043
rect 19257 20009 19291 20043
rect 23029 20009 23063 20043
rect 1133 19941 1167 19975
rect 2513 19941 2547 19975
rect 2605 19941 2639 19975
rect 5181 19941 5215 19975
rect 9045 19941 9079 19975
rect 16405 19941 16439 19975
rect 1593 19873 1627 19907
rect 1869 19873 1903 19907
rect 2053 19873 2087 19907
rect 2329 19873 2363 19907
rect 3157 19873 3191 19907
rect 3424 19873 3458 19907
rect 4813 19873 4847 19907
rect 5457 19873 5491 19907
rect 5641 19873 5675 19907
rect 6837 19873 6871 19907
rect 7113 19873 7147 19907
rect 7389 19873 7423 19907
rect 7757 19873 7791 19907
rect 7941 19873 7975 19907
rect 8401 19873 8435 19907
rect 8585 19873 8619 19907
rect 8769 19873 8803 19907
rect 8953 19873 8987 19907
rect 10977 19873 11011 19907
rect 11069 19873 11103 19907
rect 11253 19873 11287 19907
rect 11713 19873 11747 19907
rect 11805 19873 11839 19907
rect 11989 19873 12023 19907
rect 12173 19873 12207 19907
rect 12532 19873 12566 19907
rect 13737 19873 13771 19907
rect 13993 19873 14027 19907
rect 15393 19873 15427 19907
rect 15669 19873 15703 19907
rect 15761 19873 15795 19907
rect 16129 19873 16163 19907
rect 16313 19873 16347 19907
rect 16865 19873 16899 19907
rect 19533 19873 19567 19907
rect 20361 19873 20395 19907
rect 20637 19873 20671 19907
rect 21097 19873 21131 19907
rect 21465 19873 21499 19907
rect 21649 19873 21683 19907
rect 21905 19873 21939 19907
rect 1501 19805 1535 19839
rect 4905 19805 4939 19839
rect 5273 19805 5307 19839
rect 6377 19805 6411 19839
rect 6929 19805 6963 19839
rect 12265 19805 12299 19839
rect 18797 19805 18831 19839
rect 18889 19805 18923 19839
rect 18981 19805 19015 19839
rect 19073 19805 19107 19839
rect 19625 19805 19659 19839
rect 20545 19805 20579 19839
rect 5549 19737 5583 19771
rect 7849 19737 7883 19771
rect 15485 19737 15519 19771
rect 19901 19737 19935 19771
rect 20821 19737 20855 19771
rect 21281 19737 21315 19771
rect 1961 19669 1995 19703
rect 2145 19669 2179 19703
rect 2789 19669 2823 19703
rect 2973 19669 3007 19703
rect 4537 19669 4571 19703
rect 7113 19669 7147 19703
rect 7205 19669 7239 19703
rect 8493 19669 8527 19703
rect 8769 19669 8803 19703
rect 12081 19669 12115 19703
rect 15117 19669 15151 19703
rect 16313 19669 16347 19703
rect 16589 19669 16623 19703
rect 16773 19669 16807 19703
rect 18153 19669 18187 19703
rect 20177 19669 20211 19703
rect 20913 19669 20947 19703
rect 2881 19465 2915 19499
rect 3525 19465 3559 19499
rect 4905 19465 4939 19499
rect 5365 19465 5399 19499
rect 8769 19465 8803 19499
rect 10149 19465 10183 19499
rect 10425 19465 10459 19499
rect 11437 19465 11471 19499
rect 12081 19465 12115 19499
rect 12909 19465 12943 19499
rect 13737 19465 13771 19499
rect 14381 19465 14415 19499
rect 14565 19465 14599 19499
rect 20729 19465 20763 19499
rect 20821 19465 20855 19499
rect 21649 19465 21683 19499
rect 22753 19465 22787 19499
rect 2513 19397 2547 19431
rect 3801 19397 3835 19431
rect 4629 19397 4663 19431
rect 8953 19397 8987 19431
rect 16037 19397 16071 19431
rect 857 19329 891 19363
rect 9413 19329 9447 19363
rect 12541 19329 12575 19363
rect 20453 19329 20487 19363
rect 22017 19329 22051 19363
rect 22201 19329 22235 19363
rect 1685 19261 1719 19295
rect 1869 19261 1903 19295
rect 2237 19261 2271 19295
rect 2421 19261 2455 19295
rect 3433 19261 3467 19295
rect 3709 19261 3743 19295
rect 3801 19261 3835 19295
rect 3985 19261 4019 19295
rect 4169 19261 4203 19295
rect 4353 19261 4387 19295
rect 4445 19261 4479 19295
rect 4721 19261 4755 19295
rect 5181 19261 5215 19295
rect 6745 19261 6779 19295
rect 6837 19261 6871 19295
rect 9505 19261 9539 19295
rect 9965 19261 9999 19295
rect 10057 19261 10091 19295
rect 10333 19261 10367 19295
rect 10609 19261 10643 19295
rect 13553 19261 13587 19295
rect 14013 19261 14047 19295
rect 14657 19261 14691 19295
rect 16129 19261 16163 19295
rect 17601 19261 17635 19295
rect 17877 19261 17911 19295
rect 18705 19261 18739 19295
rect 20361 19261 20395 19295
rect 20821 19261 20855 19295
rect 21005 19261 21039 19295
rect 21465 19261 21499 19295
rect 21833 19261 21867 19295
rect 22109 19261 22143 19295
rect 22385 19261 22419 19295
rect 22845 19261 22879 19295
rect 6500 19193 6534 19227
rect 7104 19193 7138 19227
rect 8585 19193 8619 19227
rect 11621 19193 11655 19227
rect 11805 19193 11839 19227
rect 11897 19193 11931 19227
rect 12097 19193 12131 19227
rect 14924 19193 14958 19227
rect 16374 19193 16408 19227
rect 18972 19193 19006 19227
rect 2421 19125 2455 19159
rect 2881 19125 2915 19159
rect 3065 19125 3099 19159
rect 3249 19125 3283 19159
rect 4261 19125 4295 19159
rect 4997 19125 5031 19159
rect 8217 19125 8251 19159
rect 8785 19125 8819 19159
rect 9045 19125 9079 19159
rect 9689 19125 9723 19159
rect 12265 19125 12299 19159
rect 12909 19125 12943 19159
rect 13093 19125 13127 19159
rect 14381 19125 14415 19159
rect 17509 19125 17543 19159
rect 20085 19125 20119 19159
rect 21189 19125 21223 19159
rect 21281 19125 21315 19159
rect 22569 19125 22603 19159
rect 6193 18921 6227 18955
rect 7665 18921 7699 18955
rect 8769 18921 8803 18955
rect 12633 18921 12667 18955
rect 12909 18921 12943 18955
rect 13921 18921 13955 18955
rect 14381 18921 14415 18955
rect 15761 18921 15795 18955
rect 17049 18921 17083 18955
rect 17509 18921 17543 18955
rect 17969 18921 18003 18955
rect 18153 18921 18187 18955
rect 18429 18921 18463 18955
rect 21649 18921 21683 18955
rect 8493 18853 8527 18887
rect 11161 18853 11195 18887
rect 11621 18853 11655 18887
rect 15301 18853 15335 18887
rect 1869 18785 1903 18819
rect 2697 18785 2731 18819
rect 2973 18785 3007 18819
rect 3229 18785 3263 18819
rect 4629 18785 4663 18819
rect 5089 18785 5123 18819
rect 5365 18785 5399 18819
rect 5831 18785 5865 18819
rect 6009 18785 6043 18819
rect 6285 18785 6319 18819
rect 7297 18785 7331 18819
rect 7757 18785 7791 18819
rect 8309 18785 8343 18819
rect 8769 18785 8803 18819
rect 8861 18785 8895 18819
rect 9321 18785 9355 18819
rect 10526 18785 10560 18819
rect 10793 18785 10827 18819
rect 11805 18785 11839 18819
rect 11989 18785 12023 18819
rect 12081 18785 12115 18819
rect 12357 18785 12391 18819
rect 12449 18785 12483 18819
rect 13093 18785 13127 18819
rect 13277 18785 13311 18819
rect 13553 18785 13587 18819
rect 14105 18785 14139 18819
rect 14289 18785 14323 18819
rect 14565 18785 14599 18819
rect 14749 18785 14783 18819
rect 15577 18785 15611 18819
rect 16773 18785 16807 18819
rect 16865 18785 16899 18819
rect 17325 18785 17359 18819
rect 17601 18785 17635 18819
rect 18245 18785 18279 18819
rect 19441 18785 19475 18819
rect 19901 18785 19935 18819
rect 20545 18785 20579 18819
rect 21465 18785 21499 18819
rect 22773 18785 22807 18819
rect 1961 18717 1995 18751
rect 2513 18717 2547 18751
rect 4537 18717 4571 18751
rect 7021 18717 7055 18751
rect 7205 18717 7239 18751
rect 19165 18717 19199 18751
rect 19625 18717 19659 18751
rect 19809 18717 19843 18751
rect 20453 18717 20487 18751
rect 20913 18717 20947 18751
rect 23029 18717 23063 18751
rect 2881 18649 2915 18683
rect 4353 18649 4387 18683
rect 5273 18649 5307 18683
rect 8677 18649 8711 18683
rect 9137 18649 9171 18683
rect 11529 18649 11563 18683
rect 12173 18649 12207 18683
rect 14933 18649 14967 18683
rect 15485 18649 15519 18683
rect 20269 18649 20303 18683
rect 4905 18581 4939 18615
rect 5549 18581 5583 18615
rect 6009 18581 6043 18615
rect 9045 18581 9079 18615
rect 9413 18581 9447 18615
rect 10977 18581 11011 18615
rect 11161 18581 11195 18615
rect 13369 18581 13403 18615
rect 15301 18581 15335 18615
rect 17969 18581 18003 18615
rect 21281 18581 21315 18615
rect 4261 18377 4295 18411
rect 6469 18377 6503 18411
rect 6929 18377 6963 18411
rect 7757 18377 7791 18411
rect 8125 18377 8159 18411
rect 10425 18377 10459 18411
rect 11161 18377 11195 18411
rect 13553 18377 13587 18411
rect 13737 18377 13771 18411
rect 16773 18377 16807 18411
rect 18061 18377 18095 18411
rect 21097 18377 21131 18411
rect 1961 18309 1995 18343
rect 5917 18309 5951 18343
rect 8493 18309 8527 18343
rect 9597 18309 9631 18343
rect 13369 18309 13403 18343
rect 14933 18309 14967 18343
rect 18245 18309 18279 18343
rect 18337 18309 18371 18343
rect 22293 18309 22327 18343
rect 22845 18309 22879 18343
rect 1777 18241 1811 18275
rect 4353 18241 4387 18275
rect 7113 18241 7147 18275
rect 16221 18241 16255 18275
rect 16681 18241 16715 18275
rect 17233 18241 17267 18275
rect 17693 18241 17727 18275
rect 19441 18241 19475 18275
rect 21281 18241 21315 18275
rect 22477 18241 22511 18275
rect 2053 18173 2087 18207
rect 2881 18173 2915 18207
rect 3065 18173 3099 18207
rect 3985 18173 4019 18207
rect 4537 18173 4571 18207
rect 5089 18173 5123 18207
rect 5365 18173 5399 18207
rect 5641 18173 5675 18207
rect 6193 18173 6227 18207
rect 6653 18173 6687 18207
rect 6745 18173 6779 18207
rect 7021 18173 7055 18207
rect 7297 18173 7331 18207
rect 7389 18173 7423 18207
rect 7481 18173 7515 18207
rect 7573 18173 7607 18207
rect 7757 18173 7791 18207
rect 7941 18173 7975 18207
rect 8033 18173 8067 18207
rect 8861 18173 8895 18207
rect 8953 18173 8987 18207
rect 9137 18173 9171 18207
rect 9321 18173 9355 18207
rect 9689 18173 9723 18207
rect 9873 18173 9907 18207
rect 10241 18173 10275 18207
rect 11713 18173 11747 18207
rect 11989 18173 12023 18207
rect 14197 18173 14231 18207
rect 14841 18173 14875 18207
rect 15117 18173 15151 18207
rect 16313 18173 16347 18207
rect 17141 18173 17175 18207
rect 17417 18173 17451 18207
rect 17601 18173 17635 18207
rect 18521 18173 18555 18207
rect 19349 18173 19383 18207
rect 19708 18173 19742 18207
rect 20913 18173 20947 18207
rect 22017 18173 22051 18207
rect 22753 18173 22787 18207
rect 23029 18173 23063 18207
rect 4261 18105 4295 18139
rect 5273 18105 5307 18139
rect 5917 18105 5951 18139
rect 9597 18105 9631 18139
rect 10977 18105 11011 18139
rect 11193 18105 11227 18139
rect 12234 18105 12268 18139
rect 13721 18105 13755 18139
rect 13921 18105 13955 18139
rect 16957 18105 16991 18139
rect 18061 18105 18095 18139
rect 18705 18105 18739 18139
rect 18889 18105 18923 18139
rect 1777 18037 1811 18071
rect 2973 18037 3007 18071
rect 4169 18037 4203 18071
rect 4721 18037 4755 18071
rect 4905 18037 4939 18071
rect 5733 18037 5767 18071
rect 6009 18037 6043 18071
rect 8401 18037 8435 18071
rect 9045 18037 9079 18071
rect 9413 18037 9447 18071
rect 9781 18037 9815 18071
rect 11345 18037 11379 18071
rect 11897 18037 11931 18071
rect 14381 18037 14415 18071
rect 14657 18037 14691 18071
rect 19073 18037 19107 18071
rect 19165 18037 19199 18071
rect 20821 18037 20855 18071
rect 21465 18037 21499 18071
rect 21557 18037 21591 18071
rect 21925 18037 21959 18071
rect 22569 18037 22603 18071
rect 2329 17833 2363 17867
rect 2697 17833 2731 17867
rect 4169 17833 4203 17867
rect 4905 17833 4939 17867
rect 6193 17833 6227 17867
rect 6377 17833 6411 17867
rect 7757 17833 7791 17867
rect 8125 17833 8159 17867
rect 8769 17833 8803 17867
rect 10793 17833 10827 17867
rect 13737 17833 13771 17867
rect 17785 17833 17819 17867
rect 17953 17833 17987 17867
rect 21097 17833 21131 17867
rect 21465 17833 21499 17867
rect 5273 17765 5307 17799
rect 7297 17765 7331 17799
rect 7389 17765 7423 17799
rect 13277 17765 13311 17799
rect 15117 17765 15151 17799
rect 18153 17765 18187 17799
rect 19064 17765 19098 17799
rect 21905 17765 21939 17799
rect 1216 17697 1250 17731
rect 2421 17697 2455 17731
rect 3056 17697 3090 17731
rect 4629 17697 4663 17731
rect 4721 17697 4755 17731
rect 6009 17697 6043 17731
rect 6285 17697 6319 17731
rect 6561 17697 6595 17731
rect 6653 17697 6687 17731
rect 6929 17697 6963 17731
rect 7021 17697 7055 17731
rect 7113 17697 7147 17731
rect 8309 17697 8343 17731
rect 8401 17697 8435 17731
rect 8493 17697 8527 17731
rect 8953 17697 8987 17731
rect 9137 17697 9171 17731
rect 9229 17697 9263 17731
rect 9413 17697 9447 17731
rect 9680 17697 9714 17731
rect 10977 17697 11011 17731
rect 11233 17697 11267 17731
rect 12633 17697 12667 17731
rect 12909 17697 12943 17731
rect 13093 17697 13127 17731
rect 13829 17697 13863 17731
rect 14105 17697 14139 17731
rect 14565 17697 14599 17731
rect 14749 17697 14783 17731
rect 15025 17697 15059 17731
rect 15209 17697 15243 17731
rect 15577 17697 15611 17731
rect 15669 17697 15703 17731
rect 15853 17697 15887 17731
rect 16313 17697 16347 17731
rect 16773 17697 16807 17731
rect 16957 17697 16991 17731
rect 18797 17697 18831 17731
rect 20729 17697 20763 17731
rect 21281 17697 21315 17731
rect 21649 17697 21683 17731
rect 949 17629 983 17663
rect 2697 17629 2731 17663
rect 2789 17629 2823 17663
rect 4261 17629 4295 17663
rect 5825 17629 5859 17663
rect 6377 17629 6411 17663
rect 7573 17629 7607 17663
rect 7665 17629 7699 17663
rect 7941 17629 7975 17663
rect 8033 17629 8067 17663
rect 9045 17629 9079 17663
rect 12817 17629 12851 17663
rect 13369 17629 13403 17663
rect 14013 17629 14047 17663
rect 14657 17629 14691 17663
rect 15301 17629 15335 17663
rect 15485 17629 15519 17663
rect 16405 17629 16439 17663
rect 16865 17629 16899 17663
rect 20453 17629 20487 17663
rect 20637 17629 20671 17663
rect 5641 17561 5675 17595
rect 6745 17561 6779 17595
rect 8677 17561 8711 17595
rect 13553 17561 13587 17595
rect 15761 17561 15795 17595
rect 16681 17561 16715 17595
rect 2513 17493 2547 17527
rect 5089 17493 5123 17527
rect 5273 17493 5307 17527
rect 12357 17493 12391 17527
rect 12449 17493 12483 17527
rect 14381 17493 14415 17527
rect 15393 17493 15427 17527
rect 17969 17493 18003 17527
rect 20177 17493 20211 17527
rect 23029 17493 23063 17527
rect 1593 17289 1627 17323
rect 2237 17289 2271 17323
rect 2697 17289 2731 17323
rect 2881 17289 2915 17323
rect 6193 17289 6227 17323
rect 6653 17289 6687 17323
rect 7481 17289 7515 17323
rect 8769 17289 8803 17323
rect 9597 17289 9631 17323
rect 10793 17289 10827 17323
rect 11345 17289 11379 17323
rect 11529 17289 11563 17323
rect 13645 17289 13679 17323
rect 14197 17289 14231 17323
rect 15853 17289 15887 17323
rect 16865 17289 16899 17323
rect 5273 17221 5307 17255
rect 6101 17221 6135 17255
rect 7297 17221 7331 17255
rect 7573 17221 7607 17255
rect 8401 17221 8435 17255
rect 10241 17221 10275 17255
rect 9505 17153 9539 17187
rect 10425 17153 10459 17187
rect 11621 17153 11655 17187
rect 21281 17153 21315 17187
rect 1317 17085 1351 17119
rect 1593 17085 1627 17119
rect 1777 17085 1811 17119
rect 1961 17085 1995 17119
rect 2053 17085 2087 17119
rect 4997 17085 5031 17119
rect 5089 17085 5123 17119
rect 5917 17085 5951 17119
rect 6377 17085 6411 17119
rect 7757 17085 7791 17119
rect 9045 17085 9079 17119
rect 9689 17085 9723 17119
rect 9781 17085 9815 17119
rect 10609 17085 10643 17119
rect 13369 17085 13403 17119
rect 14105 17085 14139 17119
rect 14289 17085 14323 17119
rect 14565 17085 14599 17119
rect 14657 17085 14691 17119
rect 15117 17085 15151 17119
rect 15393 17085 15427 17119
rect 15577 17085 15611 17119
rect 15669 17085 15703 17119
rect 15853 17085 15887 17119
rect 15945 17085 15979 17119
rect 17509 17085 17543 17119
rect 18153 17085 18187 17119
rect 18245 17085 18279 17119
rect 18429 17085 18463 17119
rect 18705 17085 18739 17119
rect 18889 17085 18923 17119
rect 19441 17085 19475 17119
rect 21189 17085 21223 17119
rect 21649 17085 21683 17119
rect 21916 17085 21950 17119
rect 6607 17051 6641 17085
rect 3065 17017 3099 17051
rect 5457 17017 5491 17051
rect 5641 17017 5675 17051
rect 6837 17017 6871 17051
rect 7021 17017 7055 17051
rect 9965 17017 9999 17051
rect 11161 17017 11195 17051
rect 11361 17017 11395 17051
rect 13829 17017 13863 17051
rect 14013 17017 14047 17051
rect 14841 17017 14875 17051
rect 15025 17017 15059 17051
rect 17049 17017 17083 17051
rect 17693 17017 17727 17051
rect 17877 17017 17911 17051
rect 19165 17017 19199 17051
rect 19349 17017 19383 17051
rect 21465 17017 21499 17051
rect 1133 16949 1167 16983
rect 2865 16949 2899 16983
rect 3709 16949 3743 16983
rect 6469 16949 6503 16983
rect 8769 16949 8803 16983
rect 8953 16949 8987 16983
rect 9229 16949 9263 16983
rect 14381 16949 14415 16983
rect 15301 16949 15335 16983
rect 15577 16949 15611 16983
rect 16129 16949 16163 16983
rect 16681 16949 16715 16983
rect 16849 16949 16883 16983
rect 17969 16949 18003 16983
rect 18429 16949 18463 16983
rect 18889 16949 18923 16983
rect 23029 16949 23063 16983
rect 3893 16745 3927 16779
rect 4261 16745 4295 16779
rect 4445 16745 4479 16779
rect 5411 16745 5445 16779
rect 7665 16745 7699 16779
rect 7849 16745 7883 16779
rect 8125 16745 8159 16779
rect 10701 16745 10735 16779
rect 14749 16745 14783 16779
rect 16306 16745 16340 16779
rect 17969 16745 18003 16779
rect 20729 16745 20763 16779
rect 21465 16745 21499 16779
rect 23029 16745 23063 16779
rect 1216 16677 1250 16711
rect 3157 16677 3191 16711
rect 8309 16677 8343 16711
rect 8861 16677 8895 16711
rect 16405 16677 16439 16711
rect 19901 16677 19935 16711
rect 20085 16677 20119 16711
rect 949 16609 983 16643
rect 2421 16609 2455 16643
rect 2605 16609 2639 16643
rect 2697 16609 2731 16643
rect 2789 16609 2823 16643
rect 3433 16609 3467 16643
rect 3525 16609 3559 16643
rect 3617 16609 3651 16643
rect 3801 16609 3835 16643
rect 4077 16609 4111 16643
rect 4169 16609 4203 16643
rect 4537 16609 4571 16643
rect 5641 16609 5675 16643
rect 5825 16609 5859 16643
rect 6081 16609 6115 16643
rect 7297 16609 7331 16643
rect 7481 16609 7515 16643
rect 7757 16609 7791 16643
rect 7941 16609 7975 16643
rect 9045 16609 9079 16643
rect 9312 16609 9346 16643
rect 10609 16609 10643 16643
rect 10793 16609 10827 16643
rect 11161 16609 11195 16643
rect 11805 16609 11839 16643
rect 11989 16609 12023 16643
rect 12081 16609 12115 16643
rect 12173 16609 12207 16643
rect 12357 16609 12391 16643
rect 12541 16609 12575 16643
rect 12633 16609 12667 16643
rect 12817 16609 12851 16643
rect 13093 16609 13127 16643
rect 13369 16609 13403 16643
rect 13645 16609 13679 16643
rect 14565 16609 14599 16643
rect 14749 16609 14783 16643
rect 15025 16609 15059 16643
rect 15209 16609 15243 16643
rect 15301 16609 15335 16643
rect 15577 16609 15611 16643
rect 16129 16609 16163 16643
rect 16221 16609 16255 16643
rect 17049 16609 17083 16643
rect 17233 16609 17267 16643
rect 17417 16609 17451 16643
rect 17509 16609 17543 16643
rect 17693 16609 17727 16643
rect 17785 16609 17819 16643
rect 18705 16609 18739 16643
rect 18981 16609 19015 16643
rect 19165 16609 19199 16643
rect 19349 16609 19383 16643
rect 20361 16609 20395 16643
rect 20545 16609 20579 16643
rect 20637 16609 20671 16643
rect 20821 16609 20855 16643
rect 20913 16609 20947 16643
rect 21281 16609 21315 16643
rect 21649 16609 21683 16643
rect 21916 16609 21950 16643
rect 8401 16541 8435 16575
rect 11069 16541 11103 16575
rect 15669 16541 15703 16575
rect 18613 16541 18647 16575
rect 3065 16473 3099 16507
rect 8861 16473 8895 16507
rect 12909 16473 12943 16507
rect 14841 16473 14875 16507
rect 18337 16473 18371 16507
rect 2329 16405 2363 16439
rect 7205 16405 7239 16439
rect 10425 16405 10459 16439
rect 11529 16405 11563 16439
rect 11621 16405 11655 16439
rect 12725 16405 12759 16439
rect 13185 16405 13219 16439
rect 13461 16405 13495 16439
rect 15945 16405 15979 16439
rect 17509 16405 17543 16439
rect 19073 16405 19107 16439
rect 20269 16405 20303 16439
rect 20453 16405 20487 16439
rect 21097 16405 21131 16439
rect 6193 16201 6227 16235
rect 7757 16201 7791 16235
rect 8401 16201 8435 16235
rect 8769 16201 8803 16235
rect 9873 16201 9907 16235
rect 10701 16201 10735 16235
rect 10885 16201 10919 16235
rect 11897 16201 11931 16235
rect 16497 16201 16531 16235
rect 22109 16201 22143 16235
rect 22845 16201 22879 16235
rect 2237 16133 2271 16167
rect 6469 16133 6503 16167
rect 14105 16133 14139 16167
rect 21833 16133 21867 16167
rect 22477 16133 22511 16167
rect 857 16065 891 16099
rect 3065 16065 3099 16099
rect 4905 16065 4939 16099
rect 5733 16065 5767 16099
rect 5825 16065 5859 16099
rect 6101 16065 6135 16099
rect 7113 16065 7147 16099
rect 7389 16065 7423 16099
rect 9137 16065 9171 16099
rect 9505 16065 9539 16099
rect 10149 16065 10183 16099
rect 12633 16065 12667 16099
rect 13001 16065 13035 16099
rect 13277 16065 13311 16099
rect 14473 16065 14507 16099
rect 14933 16065 14967 16099
rect 22661 16065 22695 16099
rect 1124 15997 1158 16031
rect 2421 15997 2455 16031
rect 2881 15997 2915 16031
rect 3249 15997 3283 16031
rect 3505 15997 3539 16031
rect 5641 15997 5675 16031
rect 5917 15997 5951 16031
rect 6377 15997 6411 16031
rect 6561 15997 6595 16031
rect 6653 15997 6687 16031
rect 6837 15997 6871 16031
rect 7021 15997 7055 16031
rect 8033 15997 8067 16031
rect 8217 15997 8251 16031
rect 8585 15997 8619 16031
rect 8953 15997 8987 16031
rect 9045 15997 9079 16031
rect 9229 15997 9263 16031
rect 9597 15997 9631 16031
rect 10057 15997 10091 16031
rect 10241 15997 10275 16031
rect 10333 15997 10367 16031
rect 10609 15997 10643 16031
rect 10786 15997 10820 16031
rect 11069 15997 11103 16031
rect 11253 15997 11287 16031
rect 11529 15997 11563 16031
rect 11805 15997 11839 16031
rect 11989 15997 12023 16031
rect 12449 15997 12483 16031
rect 12909 15997 12943 16031
rect 13553 15997 13587 16031
rect 13737 15997 13771 16031
rect 14381 15997 14415 16031
rect 14841 15997 14875 16031
rect 16405 15997 16439 16031
rect 16681 15997 16715 16031
rect 17049 15997 17083 16031
rect 19809 15997 19843 16031
rect 20085 15997 20119 16031
rect 20269 15997 20303 16031
rect 21373 15997 21407 16031
rect 21557 15997 21591 16031
rect 21649 15997 21683 16031
rect 21925 15997 21959 16031
rect 22293 15997 22327 16031
rect 22569 15997 22603 16031
rect 22753 15997 22787 16031
rect 23029 15997 23063 16031
rect 7481 15929 7515 15963
rect 7598 15929 7632 15963
rect 12081 15929 12115 15963
rect 12173 15929 12207 15963
rect 13829 15929 13863 15963
rect 2605 15861 2639 15895
rect 2697 15861 2731 15895
rect 4629 15861 4663 15895
rect 4997 15861 5031 15895
rect 5089 15861 5123 15895
rect 5457 15861 5491 15895
rect 6929 15861 6963 15895
rect 8033 15861 8067 15895
rect 10517 15861 10551 15895
rect 11345 15861 11379 15895
rect 13737 15861 13771 15895
rect 15209 15861 15243 15895
rect 16221 15861 16255 15895
rect 17233 15861 17267 15895
rect 19993 15861 20027 15895
rect 20269 15861 20303 15895
rect 21465 15861 21499 15895
rect 2973 15657 3007 15691
rect 3801 15657 3835 15691
rect 6469 15657 6503 15691
rect 6929 15657 6963 15691
rect 11161 15657 11195 15691
rect 13737 15657 13771 15691
rect 13921 15657 13955 15691
rect 15393 15657 15427 15691
rect 19533 15657 19567 15691
rect 22845 15657 22879 15691
rect 1225 15589 1259 15623
rect 1441 15589 1475 15623
rect 1777 15589 1811 15623
rect 2421 15589 2455 15623
rect 3893 15589 3927 15623
rect 5641 15589 5675 15623
rect 8401 15589 8435 15623
rect 8617 15589 8651 15623
rect 10517 15589 10551 15623
rect 10701 15589 10735 15623
rect 12265 15589 12299 15623
rect 20637 15589 20671 15623
rect 21005 15589 21039 15623
rect 22385 15589 22419 15623
rect 1685 15521 1719 15555
rect 1869 15521 1903 15555
rect 2605 15521 2639 15555
rect 2881 15521 2915 15555
rect 6009 15521 6043 15555
rect 7113 15521 7147 15555
rect 7205 15521 7239 15555
rect 7389 15521 7423 15555
rect 7665 15521 7699 15555
rect 8309 15505 8343 15539
rect 9689 15521 9723 15555
rect 9873 15521 9907 15555
rect 10241 15521 10275 15555
rect 10977 15521 11011 15555
rect 12449 15521 12483 15555
rect 12725 15521 12759 15555
rect 12909 15521 12943 15555
rect 13369 15521 13403 15555
rect 13553 15521 13587 15555
rect 13829 15521 13863 15555
rect 14013 15521 14047 15555
rect 14657 15521 14691 15555
rect 15025 15521 15059 15555
rect 15117 15521 15151 15555
rect 15577 15521 15611 15555
rect 15669 15521 15703 15555
rect 16589 15521 16623 15555
rect 17877 15521 17911 15555
rect 18337 15521 18371 15555
rect 18613 15521 18647 15555
rect 18797 15521 18831 15555
rect 18889 15521 18923 15555
rect 19073 15521 19107 15555
rect 19441 15521 19475 15555
rect 19901 15521 19935 15555
rect 20361 15521 20395 15555
rect 20913 15521 20947 15555
rect 21097 15521 21131 15555
rect 21649 15521 21683 15555
rect 21833 15521 21867 15555
rect 21925 15521 21959 15555
rect 22017 15521 22051 15555
rect 22201 15521 22235 15555
rect 22293 15521 22327 15555
rect 22569 15521 22603 15555
rect 22753 15521 22787 15555
rect 23029 15521 23063 15555
rect 2789 15453 2823 15487
rect 3341 15453 3375 15487
rect 6285 15453 6319 15487
rect 6377 15453 6411 15487
rect 7297 15453 7331 15487
rect 9229 15453 9263 15487
rect 9321 15453 9355 15487
rect 9413 15453 9447 15487
rect 9505 15453 9539 15487
rect 16681 15453 16715 15487
rect 16957 15453 16991 15487
rect 17233 15453 17267 15487
rect 17325 15453 17359 15487
rect 17417 15453 17451 15487
rect 17509 15453 17543 15487
rect 17693 15453 17727 15487
rect 18061 15453 18095 15487
rect 18153 15453 18187 15487
rect 18705 15453 18739 15487
rect 18981 15453 19015 15487
rect 19993 15453 20027 15487
rect 20637 15453 20671 15487
rect 3617 15385 3651 15419
rect 5825 15385 5859 15419
rect 7481 15385 7515 15419
rect 9873 15385 9907 15419
rect 10333 15385 10367 15419
rect 14473 15385 14507 15419
rect 15301 15385 15335 15419
rect 15853 15385 15887 15419
rect 18521 15385 18555 15419
rect 22109 15385 22143 15419
rect 1409 15317 1443 15351
rect 1593 15317 1627 15351
rect 6837 15317 6871 15351
rect 8125 15317 8159 15351
rect 8585 15317 8619 15351
rect 8769 15317 8803 15351
rect 9045 15317 9079 15351
rect 12633 15317 12667 15351
rect 12817 15317 12851 15351
rect 14841 15317 14875 15351
rect 17049 15317 17083 15351
rect 20269 15317 20303 15351
rect 20453 15317 20487 15351
rect 21465 15317 21499 15351
rect 22569 15317 22603 15351
rect 4445 15113 4479 15147
rect 6377 15113 6411 15147
rect 6837 15113 6871 15147
rect 9137 15113 9171 15147
rect 10333 15113 10367 15147
rect 14657 15113 14691 15147
rect 16405 15113 16439 15147
rect 6469 15045 6503 15079
rect 11529 15045 11563 15079
rect 15485 15045 15519 15079
rect 19349 15045 19383 15079
rect 19901 15045 19935 15079
rect 20453 15045 20487 15079
rect 2513 14977 2547 15011
rect 2973 14977 3007 15011
rect 8585 14977 8619 15011
rect 9321 14977 9355 15011
rect 11805 14977 11839 15011
rect 11943 14977 11977 15011
rect 15025 14977 15059 15011
rect 15945 14977 15979 15011
rect 16589 14977 16623 15011
rect 16773 14977 16807 15011
rect 17233 14977 17267 15011
rect 18889 14977 18923 15011
rect 18981 14977 19015 15011
rect 19165 14977 19199 15011
rect 22569 14977 22603 15011
rect 2329 14909 2363 14943
rect 2605 14909 2639 14943
rect 3341 14909 3375 14943
rect 3801 14909 3835 14943
rect 3985 14909 4019 14943
rect 4261 14909 4295 14943
rect 4997 14909 5031 14943
rect 5089 14909 5123 14943
rect 5849 14909 5883 14943
rect 6193 14909 6227 14943
rect 6653 14909 6687 14943
rect 6929 14909 6963 14943
rect 7021 14909 7055 14943
rect 7297 14909 7331 14943
rect 8217 14909 8251 14943
rect 9597 14909 9631 14943
rect 10241 14909 10275 14943
rect 10425 14909 10459 14943
rect 10609 14909 10643 14943
rect 10885 14909 10919 14943
rect 11069 14909 11103 14943
rect 12081 14909 12115 14943
rect 12817 14909 12851 14943
rect 13001 14909 13035 14943
rect 13093 14909 13127 14943
rect 13553 14909 13587 14943
rect 14013 14909 14047 14943
rect 14197 14909 14231 14943
rect 14749 14909 14783 14943
rect 15117 14909 15151 14943
rect 15853 14909 15887 14943
rect 16313 14909 16347 14943
rect 16681 14909 16715 14943
rect 16865 14909 16899 14943
rect 17141 14909 17175 14943
rect 19073 14909 19107 14943
rect 19533 14909 19567 14943
rect 21005 14909 21039 14943
rect 22477 14909 22511 14943
rect 2084 14841 2118 14875
rect 4721 14841 4755 14875
rect 5457 14841 5491 14875
rect 13737 14841 13771 14875
rect 13921 14841 13955 14875
rect 19625 14841 19659 14875
rect 20177 14841 20211 14875
rect 949 14773 983 14807
rect 3525 14773 3559 14807
rect 3709 14773 3743 14807
rect 4077 14773 4111 14807
rect 6009 14773 6043 14807
rect 8033 14773 8067 14807
rect 8677 14773 8711 14807
rect 8769 14773 8803 14807
rect 10793 14773 10827 14807
rect 12725 14773 12759 14807
rect 12909 14773 12943 14807
rect 13277 14773 13311 14807
rect 14197 14773 14231 14807
rect 16221 14773 16255 14807
rect 16589 14773 16623 14807
rect 17509 14773 17543 14807
rect 18705 14773 18739 14807
rect 20085 14773 20119 14807
rect 20637 14773 20671 14807
rect 21189 14773 21223 14807
rect 22109 14773 22143 14807
rect 1409 14569 1443 14603
rect 3433 14569 3467 14603
rect 3985 14569 4019 14603
rect 4261 14569 4295 14603
rect 7573 14569 7607 14603
rect 8493 14569 8527 14603
rect 9045 14569 9079 14603
rect 11345 14569 11379 14603
rect 12265 14569 12299 14603
rect 17417 14569 17451 14603
rect 17693 14569 17727 14603
rect 1317 14501 1351 14535
rect 1777 14501 1811 14535
rect 4997 14501 5031 14535
rect 5365 14501 5399 14535
rect 7941 14501 7975 14535
rect 12173 14501 12207 14535
rect 13737 14501 13771 14535
rect 21373 14501 21407 14535
rect 1041 14433 1075 14467
rect 1133 14433 1167 14467
rect 1593 14433 1627 14467
rect 2053 14433 2087 14467
rect 2329 14433 2363 14467
rect 2973 14433 3007 14467
rect 3617 14433 3651 14467
rect 3801 14433 3835 14467
rect 4537 14433 4571 14467
rect 4629 14433 4663 14467
rect 6101 14433 6135 14467
rect 7021 14433 7055 14467
rect 7481 14433 7515 14467
rect 7757 14433 7791 14467
rect 8401 14433 8435 14467
rect 8585 14433 8619 14467
rect 8677 14433 8711 14467
rect 8861 14433 8895 14467
rect 9229 14433 9263 14467
rect 9413 14433 9447 14467
rect 9597 14433 9631 14467
rect 9689 14433 9723 14467
rect 9781 14433 9815 14467
rect 10149 14433 10183 14467
rect 10333 14433 10367 14467
rect 11529 14433 11563 14467
rect 11805 14433 11839 14467
rect 12817 14433 12851 14467
rect 14013 14433 14047 14467
rect 14657 14433 14691 14467
rect 15301 14433 15335 14467
rect 17601 14433 17635 14467
rect 17693 14433 17727 14467
rect 17877 14433 17911 14467
rect 20177 14433 20211 14467
rect 20361 14433 20395 14467
rect 20453 14433 20487 14467
rect 21557 14433 21591 14467
rect 22017 14433 22051 14467
rect 22109 14433 22143 14467
rect 22293 14433 22327 14467
rect 2421 14365 2455 14399
rect 2881 14365 2915 14399
rect 5825 14365 5859 14399
rect 7205 14365 7239 14399
rect 12081 14365 12115 14399
rect 13093 14365 13127 14399
rect 13921 14365 13955 14399
rect 14381 14365 14415 14399
rect 14749 14365 14783 14399
rect 15117 14365 15151 14399
rect 19073 14365 19107 14399
rect 19349 14365 19383 14399
rect 21741 14365 21775 14399
rect 2697 14297 2731 14331
rect 1869 14229 1903 14263
rect 3249 14229 3283 14263
rect 5549 14229 5583 14263
rect 6837 14229 6871 14263
rect 10057 14229 10091 14263
rect 10241 14229 10275 14263
rect 11621 14229 11655 14263
rect 12633 14229 12667 14263
rect 15025 14229 15059 14263
rect 15485 14229 15519 14263
rect 19993 14229 20027 14263
rect 21833 14229 21867 14263
rect 22201 14229 22235 14263
rect 2973 14025 3007 14059
rect 6009 14025 6043 14059
rect 10793 14025 10827 14059
rect 12541 14025 12575 14059
rect 13921 14025 13955 14059
rect 2881 13957 2915 13991
rect 8125 13957 8159 13991
rect 9873 13957 9907 13991
rect 10977 13957 11011 13991
rect 13093 13957 13127 13991
rect 13737 13957 13771 13991
rect 16773 13957 16807 13991
rect 20729 13957 20763 13991
rect 22109 13957 22143 13991
rect 3065 13889 3099 13923
rect 12173 13889 12207 13923
rect 15393 13889 15427 13923
rect 17325 13889 17359 13923
rect 19165 13889 19199 13923
rect 19441 13889 19475 13923
rect 20269 13889 20303 13923
rect 21557 13889 21591 13923
rect 22017 13889 22051 13923
rect 22385 13889 22419 13923
rect 857 13821 891 13855
rect 1317 13821 1351 13855
rect 1584 13821 1618 13855
rect 2789 13821 2823 13855
rect 3709 13821 3743 13855
rect 3893 13821 3927 13855
rect 5825 13821 5859 13855
rect 7205 13821 7239 13855
rect 8953 13821 8987 13855
rect 10149 13821 10183 13855
rect 10425 13821 10459 13855
rect 10793 13821 10827 13855
rect 11621 13821 11655 13855
rect 11897 13821 11931 13855
rect 12357 13821 12391 13855
rect 12633 13821 12667 13855
rect 12909 13821 12943 13855
rect 13369 13821 13403 13855
rect 13553 13821 13587 13855
rect 13829 13821 13863 13855
rect 14013 13821 14047 13855
rect 14657 13821 14691 13855
rect 14933 13821 14967 13855
rect 15025 13821 15059 13855
rect 15209 13821 15243 13855
rect 15301 13821 15335 13855
rect 15485 13821 15519 13855
rect 16037 13821 16071 13855
rect 16221 13821 16255 13855
rect 16497 13821 16531 13855
rect 16773 13821 16807 13855
rect 16957 13821 16991 13855
rect 17049 13821 17083 13855
rect 18245 13821 18279 13855
rect 19073 13821 19107 13855
rect 19349 13821 19383 13855
rect 19533 13821 19567 13855
rect 19625 13821 19659 13855
rect 19809 13821 19843 13855
rect 19901 13821 19935 13855
rect 20361 13821 20395 13855
rect 21097 13821 21131 13855
rect 21649 13821 21683 13855
rect 22477 13821 22511 13855
rect 1041 13753 1075 13787
rect 7113 13753 7147 13787
rect 7573 13753 7607 13787
rect 8861 13753 8895 13787
rect 9321 13753 9355 13787
rect 9689 13753 9723 13787
rect 12725 13753 12759 13787
rect 14473 13753 14507 13787
rect 16313 13753 16347 13787
rect 18429 13753 18463 13787
rect 1225 13685 1259 13719
rect 2697 13685 2731 13719
rect 4077 13685 4111 13719
rect 6837 13685 6871 13719
rect 7941 13685 7975 13719
rect 8585 13685 8619 13719
rect 10333 13685 10367 13719
rect 13185 13685 13219 13719
rect 14841 13685 14875 13719
rect 15117 13685 15151 13719
rect 16221 13685 16255 13719
rect 16681 13685 16715 13719
rect 17555 13685 17589 13719
rect 18705 13685 18739 13719
rect 19901 13685 19935 13719
rect 19993 13685 20027 13719
rect 20637 13685 20671 13719
rect 1869 13481 1903 13515
rect 2053 13481 2087 13515
rect 6285 13481 6319 13515
rect 8677 13481 8711 13515
rect 9873 13481 9907 13515
rect 10609 13481 10643 13515
rect 10977 13481 11011 13515
rect 16681 13481 16715 13515
rect 19441 13481 19475 13515
rect 1225 13413 1259 13447
rect 2881 13413 2915 13447
rect 6561 13413 6595 13447
rect 7021 13413 7055 13447
rect 7389 13413 7423 13447
rect 11805 13413 11839 13447
rect 11989 13413 12023 13447
rect 857 13345 891 13379
rect 1501 13345 1535 13379
rect 2605 13345 2639 13379
rect 3157 13345 3191 13379
rect 3617 13345 3651 13379
rect 4261 13345 4295 13379
rect 5825 13345 5859 13379
rect 6653 13345 6687 13379
rect 8493 13345 8527 13379
rect 9229 13345 9263 13379
rect 9413 13345 9447 13379
rect 9505 13345 9539 13379
rect 9597 13345 9631 13379
rect 10241 13345 10275 13379
rect 10517 13345 10551 13379
rect 10793 13345 10827 13379
rect 11253 13345 11287 13379
rect 11345 13345 11379 13379
rect 11621 13345 11655 13379
rect 12449 13345 12483 13379
rect 12541 13345 12575 13379
rect 13093 13345 13127 13379
rect 13921 13345 13955 13379
rect 15117 13345 15151 13379
rect 16313 13345 16347 13379
rect 16773 13345 16807 13379
rect 16957 13345 16991 13379
rect 17233 13345 17267 13379
rect 17509 13345 17543 13379
rect 17693 13345 17727 13379
rect 17969 13345 18003 13379
rect 19625 13345 19659 13379
rect 2237 13277 2271 13311
rect 2697 13277 2731 13311
rect 3709 13277 3743 13311
rect 3985 13277 4019 13311
rect 4169 13277 4203 13311
rect 11161 13277 11195 13311
rect 11437 13277 11471 13311
rect 12817 13277 12851 13311
rect 13829 13277 13863 13311
rect 15025 13277 15059 13311
rect 16221 13277 16255 13311
rect 16865 13277 16899 13311
rect 17877 13277 17911 13311
rect 2973 13209 3007 13243
rect 4629 13209 4663 13243
rect 6009 13209 6043 13243
rect 7573 13209 7607 13243
rect 9965 13209 9999 13243
rect 1225 13141 1259 13175
rect 1409 13141 1443 13175
rect 1869 13141 1903 13175
rect 10149 13141 10183 13175
rect 12725 13141 12759 13175
rect 14197 13141 14231 13175
rect 14841 13141 14875 13175
rect 17049 13141 17083 13175
rect 18245 13141 18279 13175
rect 949 12937 983 12971
rect 1133 12937 1167 12971
rect 6745 12937 6779 12971
rect 9505 12937 9539 12971
rect 10977 12937 11011 12971
rect 11897 12937 11931 12971
rect 14657 12937 14691 12971
rect 19441 12937 19475 12971
rect 1685 12869 1719 12903
rect 7481 12869 7515 12903
rect 9965 12869 9999 12903
rect 11621 12869 11655 12903
rect 13093 12869 13127 12903
rect 14565 12869 14599 12903
rect 15209 12869 15243 12903
rect 16865 12869 16899 12903
rect 17417 12869 17451 12903
rect 20085 12869 20119 12903
rect 7021 12801 7055 12835
rect 11437 12801 11471 12835
rect 14105 12801 14139 12835
rect 17601 12801 17635 12835
rect 18797 12801 18831 12835
rect 19257 12801 19291 12835
rect 20545 12801 20579 12835
rect 20729 12801 20763 12835
rect 2605 12733 2639 12767
rect 3433 12733 3467 12767
rect 3617 12733 3651 12767
rect 3893 12733 3927 12767
rect 4169 12733 4203 12767
rect 4629 12733 4663 12767
rect 6561 12733 6595 12767
rect 7113 12733 7147 12767
rect 7573 12733 7607 12767
rect 8585 12733 8619 12767
rect 8769 12733 8803 12767
rect 9689 12733 9723 12767
rect 9781 12733 9815 12767
rect 10057 12733 10091 12767
rect 10149 12733 10183 12767
rect 10333 12733 10367 12767
rect 11161 12733 11195 12767
rect 11253 12733 11287 12767
rect 11529 12733 11563 12767
rect 12081 12733 12115 12767
rect 12357 12733 12391 12767
rect 12909 12733 12943 12767
rect 14197 12733 14231 12767
rect 14841 12733 14875 12767
rect 15117 12733 15151 12767
rect 15393 12733 15427 12767
rect 16773 12733 16807 12767
rect 16957 12733 16991 12767
rect 17049 12733 17083 12767
rect 17325 12733 17359 12767
rect 18889 12733 18923 12767
rect 19349 12733 19383 12767
rect 19526 12733 19560 12767
rect 19901 12733 19935 12767
rect 20085 12733 20119 12767
rect 20821 12733 20855 12767
rect 21373 12733 21407 12767
rect 1087 12699 1121 12733
rect 1317 12665 1351 12699
rect 2145 12665 2179 12699
rect 2329 12665 2363 12699
rect 3709 12665 3743 12699
rect 4077 12665 4111 12699
rect 5365 12665 5399 12699
rect 5457 12665 5491 12699
rect 5825 12665 5859 12699
rect 6193 12665 6227 12699
rect 15025 12665 15059 12699
rect 15301 12665 15335 12699
rect 21618 12665 21652 12699
rect 1961 12597 1995 12631
rect 2421 12597 2455 12631
rect 3525 12597 3559 12631
rect 4813 12597 4847 12631
rect 5089 12597 5123 12631
rect 6377 12597 6411 12631
rect 7757 12597 7791 12631
rect 8677 12597 8711 12631
rect 10333 12597 10367 12631
rect 12173 12597 12207 12631
rect 17233 12597 17267 12631
rect 17601 12597 17635 12631
rect 21189 12597 21223 12631
rect 22753 12597 22787 12631
rect 949 12393 983 12427
rect 1777 12393 1811 12427
rect 15301 12393 15335 12427
rect 17049 12393 17083 12427
rect 18245 12393 18279 12427
rect 18429 12393 18463 12427
rect 19901 12393 19935 12427
rect 21465 12393 21499 12427
rect 2320 12325 2354 12359
rect 4445 12325 4479 12359
rect 4721 12325 4755 12359
rect 7757 12325 7791 12359
rect 15485 12325 15519 12359
rect 16497 12325 16531 12359
rect 1133 12257 1167 12291
rect 2053 12257 2087 12291
rect 3525 12257 3559 12291
rect 3709 12257 3743 12291
rect 3801 12257 3835 12291
rect 4261 12257 4295 12291
rect 4353 12257 4387 12291
rect 4537 12257 4571 12291
rect 4629 12257 4663 12291
rect 4813 12257 4847 12291
rect 5457 12257 5491 12291
rect 6009 12257 6043 12291
rect 6561 12257 6595 12291
rect 6745 12257 6779 12291
rect 7021 12257 7055 12291
rect 7297 12257 7331 12291
rect 7481 12257 7515 12291
rect 7573 12257 7607 12291
rect 8309 12257 8343 12291
rect 8401 12257 8435 12291
rect 8677 12257 8711 12291
rect 8769 12257 8803 12291
rect 8861 12257 8895 12291
rect 9137 12257 9171 12291
rect 11713 12257 11747 12291
rect 11805 12257 11839 12291
rect 12633 12257 12667 12291
rect 13369 12257 13403 12291
rect 15117 12257 15151 12291
rect 15393 12257 15427 12291
rect 15669 12257 15703 12291
rect 16313 12257 16347 12291
rect 16405 12257 16439 12291
rect 16681 12257 16715 12291
rect 16773 12257 16807 12291
rect 16865 12257 16899 12291
rect 17141 12257 17175 12291
rect 17785 12257 17819 12291
rect 17969 12257 18003 12291
rect 18061 12257 18095 12291
rect 18337 12257 18371 12291
rect 18613 12257 18647 12291
rect 19257 12257 19291 12291
rect 19349 12257 19383 12291
rect 19441 12257 19475 12291
rect 19533 12257 19567 12291
rect 20085 12257 20119 12291
rect 20729 12257 20763 12291
rect 21281 12257 21315 12291
rect 22762 12257 22796 12291
rect 23029 12257 23063 12291
rect 1317 12189 1351 12223
rect 4905 12189 4939 12223
rect 5549 12189 5583 12223
rect 5917 12189 5951 12223
rect 6653 12189 6687 12223
rect 12265 12189 12299 12223
rect 12541 12189 12575 12223
rect 13001 12189 13035 12223
rect 13277 12189 13311 12223
rect 20269 12189 20303 12223
rect 20545 12189 20579 12223
rect 20637 12189 20671 12223
rect 1409 12121 1443 12155
rect 1961 12121 1995 12155
rect 3433 12121 3467 12155
rect 5181 12121 5215 12155
rect 6377 12121 6411 12155
rect 16865 12121 16899 12155
rect 1777 12053 1811 12087
rect 3709 12053 3743 12087
rect 3985 12053 4019 12087
rect 4077 12053 4111 12087
rect 6837 12053 6871 12087
rect 7941 12053 7975 12087
rect 8585 12053 8619 12087
rect 8953 12053 8987 12087
rect 13645 12053 13679 12087
rect 14933 12053 14967 12087
rect 15853 12053 15887 12087
rect 16129 12053 16163 12087
rect 17969 12053 18003 12087
rect 18797 12053 18831 12087
rect 19073 12053 19107 12087
rect 21097 12053 21131 12087
rect 21649 12053 21683 12087
rect 1133 11849 1167 11883
rect 2421 11849 2455 11883
rect 5089 11849 5123 11883
rect 10057 11849 10091 11883
rect 16865 11849 16899 11883
rect 16957 11849 16991 11883
rect 17601 11849 17635 11883
rect 18797 11849 18831 11883
rect 19533 11849 19567 11883
rect 20085 11849 20119 11883
rect 21649 11849 21683 11883
rect 17969 11781 18003 11815
rect 19165 11781 19199 11815
rect 20177 11781 20211 11815
rect 1409 11713 1443 11747
rect 1593 11713 1627 11747
rect 1685 11713 1719 11747
rect 1777 11713 1811 11747
rect 4261 11713 4295 11747
rect 8953 11713 8987 11747
rect 9413 11713 9447 11747
rect 9965 11713 9999 11747
rect 11437 11713 11471 11747
rect 11529 11713 11563 11747
rect 11897 11713 11931 11747
rect 12173 11713 12207 11747
rect 15393 11713 15427 11747
rect 15485 11713 15519 11747
rect 15577 11713 15611 11747
rect 17693 11713 17727 11747
rect 18705 11713 18739 11747
rect 19349 11713 19383 11747
rect 19993 11713 20027 11747
rect 1869 11645 1903 11679
rect 2237 11645 2271 11679
rect 2789 11645 2823 11679
rect 2881 11645 2915 11679
rect 3065 11645 3099 11679
rect 3433 11645 3467 11679
rect 3709 11645 3743 11679
rect 3893 11645 3927 11679
rect 4169 11645 4203 11679
rect 4813 11645 4847 11679
rect 5457 11645 5491 11679
rect 8585 11645 8619 11679
rect 9045 11645 9079 11679
rect 9689 11645 9723 11679
rect 9873 11645 9907 11679
rect 10241 11645 10275 11679
rect 10425 11645 10459 11679
rect 10517 11645 10551 11679
rect 10793 11645 10827 11679
rect 11253 11645 11287 11679
rect 11805 11645 11839 11679
rect 13001 11645 13035 11679
rect 13277 11645 13311 11679
rect 13737 11645 13771 11679
rect 13829 11645 13863 11679
rect 14013 11645 14047 11679
rect 14289 11645 14323 11679
rect 14473 11645 14507 11679
rect 14933 11645 14967 11679
rect 15117 11645 15151 11679
rect 15301 11645 15335 11679
rect 16589 11645 16623 11679
rect 16681 11645 16715 11679
rect 16865 11645 16899 11679
rect 17141 11645 17175 11679
rect 17417 11645 17451 11679
rect 17877 11645 17911 11679
rect 18245 11645 18279 11679
rect 18981 11645 19015 11679
rect 19625 11645 19659 11679
rect 20269 11645 20303 11679
rect 20913 11645 20947 11679
rect 21373 11645 21407 11679
rect 21465 11645 21499 11679
rect 21925 11645 21959 11679
rect 22201 11645 22235 11679
rect 22477 11645 22511 11679
rect 1117 11577 1151 11611
rect 1317 11577 1351 11611
rect 2053 11577 2087 11611
rect 3249 11577 3283 11611
rect 5273 11577 5307 11611
rect 15025 11577 15059 11611
rect 17785 11577 17819 11611
rect 18153 11577 18187 11611
rect 19349 11577 19383 11611
rect 21281 11577 21315 11611
rect 949 11509 983 11543
rect 4537 11509 4571 11543
rect 4629 11509 4663 11543
rect 8401 11509 8435 11543
rect 9781 11509 9815 11543
rect 10609 11509 10643 11543
rect 10977 11509 11011 11543
rect 11069 11509 11103 11543
rect 12817 11509 12851 11543
rect 13185 11509 13219 11543
rect 14197 11509 14231 11543
rect 14381 11509 14415 11543
rect 15761 11509 15795 11543
rect 17233 11509 17267 11543
rect 20729 11509 20763 11543
rect 21741 11509 21775 11543
rect 22017 11509 22051 11543
rect 22293 11509 22327 11543
rect 2789 11305 2823 11339
rect 4537 11305 4571 11339
rect 8401 11305 8435 11339
rect 8769 11305 8803 11339
rect 11161 11305 11195 11339
rect 11621 11305 11655 11339
rect 14013 11305 14047 11339
rect 14933 11305 14967 11339
rect 15669 11305 15703 11339
rect 18521 11305 18555 11339
rect 3893 11237 3927 11271
rect 5089 11237 5123 11271
rect 6653 11237 6687 11271
rect 12449 11237 12483 11271
rect 13461 11237 13495 11271
rect 15853 11237 15887 11271
rect 20269 11237 20303 11271
rect 21916 11237 21950 11271
rect 1308 11169 1342 11203
rect 2605 11169 2639 11203
rect 3065 11169 3099 11203
rect 3249 11169 3283 11203
rect 3341 11169 3375 11203
rect 3617 11169 3651 11203
rect 3801 11169 3835 11203
rect 4077 11169 4111 11203
rect 4353 11169 4387 11203
rect 4721 11169 4755 11203
rect 4905 11169 4939 11203
rect 5457 11169 5491 11203
rect 5641 11169 5675 11203
rect 6009 11169 6043 11203
rect 6561 11169 6595 11203
rect 6745 11169 6779 11203
rect 7021 11169 7055 11203
rect 7757 11169 7791 11203
rect 7849 11169 7883 11203
rect 8585 11169 8619 11203
rect 8861 11169 8895 11203
rect 10149 11169 10183 11203
rect 11069 11169 11103 11203
rect 11345 11169 11379 11203
rect 11621 11169 11655 11203
rect 11805 11169 11839 11203
rect 12173 11169 12207 11203
rect 12633 11169 12667 11203
rect 12725 11169 12759 11203
rect 13001 11169 13035 11203
rect 13277 11169 13311 11203
rect 13369 11169 13403 11203
rect 13645 11169 13679 11203
rect 13737 11169 13771 11203
rect 14010 11169 14044 11203
rect 14381 11169 14415 11203
rect 14473 11169 14507 11203
rect 14749 11169 14783 11203
rect 14933 11169 14967 11203
rect 15025 11169 15059 11203
rect 15301 11169 15335 11203
rect 15485 11169 15519 11203
rect 15577 11169 15611 11203
rect 16313 11169 16347 11203
rect 18429 11169 18463 11203
rect 18613 11169 18647 11203
rect 18705 11169 18739 11203
rect 18889 11169 18923 11203
rect 19165 11169 19199 11203
rect 19257 11169 19291 11203
rect 19901 11169 19935 11203
rect 20085 11169 20119 11203
rect 20177 11169 20211 11203
rect 20361 11169 20395 11203
rect 20545 11169 20579 11203
rect 20729 11169 20763 11203
rect 21097 11169 21131 11203
rect 21465 11169 21499 11203
rect 21649 11169 21683 11203
rect 1041 11101 1075 11135
rect 2881 11101 2915 11135
rect 4261 11101 4295 11135
rect 5549 11101 5583 11135
rect 6101 11101 6135 11135
rect 6377 11101 6411 11135
rect 7113 11101 7147 11135
rect 7573 11101 7607 11135
rect 7665 11101 7699 11135
rect 8033 11101 8067 11135
rect 15117 11101 15151 11135
rect 17141 11101 17175 11135
rect 17417 11101 17451 11135
rect 17509 11101 17543 11135
rect 17785 11101 17819 11135
rect 18797 11101 18831 11135
rect 19717 11101 19751 11135
rect 7389 11033 7423 11067
rect 11529 11033 11563 11067
rect 11989 11033 12023 11067
rect 12909 11033 12943 11067
rect 13093 11033 13127 11067
rect 13829 11033 13863 11067
rect 16129 11033 16163 11067
rect 21281 11033 21315 11067
rect 2421 10965 2455 10999
rect 3433 10965 3467 10999
rect 10333 10965 10367 10999
rect 12449 10965 12483 10999
rect 15853 10965 15887 10999
rect 18981 10965 19015 10999
rect 19441 10965 19475 10999
rect 21005 10965 21039 10999
rect 23029 10965 23063 10999
rect 1225 10761 1259 10795
rect 1869 10761 1903 10795
rect 5365 10761 5399 10795
rect 6377 10761 6411 10795
rect 6929 10761 6963 10795
rect 7389 10761 7423 10795
rect 11161 10761 11195 10795
rect 14197 10761 14231 10795
rect 14841 10761 14875 10795
rect 16589 10761 16623 10795
rect 17785 10761 17819 10795
rect 20085 10761 20119 10795
rect 21373 10761 21407 10795
rect 22477 10761 22511 10795
rect 1409 10693 1443 10727
rect 3893 10693 3927 10727
rect 9045 10693 9079 10727
rect 10517 10693 10551 10727
rect 12173 10693 12207 10727
rect 20729 10693 20763 10727
rect 2053 10625 2087 10659
rect 3433 10625 3467 10659
rect 4261 10625 4295 10659
rect 5549 10625 5583 10659
rect 5917 10625 5951 10659
rect 6009 10625 6043 10659
rect 8769 10625 8803 10659
rect 10057 10625 10091 10659
rect 11621 10625 11655 10659
rect 11713 10625 11747 10659
rect 12817 10625 12851 10659
rect 12909 10625 12943 10659
rect 15025 10625 15059 10659
rect 15117 10625 15151 10659
rect 15301 10625 15335 10659
rect 17049 10625 17083 10659
rect 18705 10625 18739 10659
rect 21005 10625 21039 10659
rect 21833 10625 21867 10659
rect 1041 10557 1075 10591
rect 1317 10557 1351 10591
rect 1501 10557 1535 10591
rect 1685 10557 1719 10591
rect 2329 10557 2363 10591
rect 3525 10557 3559 10591
rect 4353 10557 4387 10591
rect 5273 10557 5307 10591
rect 5457 10557 5491 10591
rect 6561 10557 6595 10591
rect 6745 10557 6779 10591
rect 7205 10557 7239 10591
rect 8677 10557 8711 10591
rect 9137 10557 9171 10591
rect 9321 10557 9355 10591
rect 10149 10557 10183 10591
rect 10241 10557 10275 10591
rect 10333 10557 10367 10591
rect 10517 10557 10551 10591
rect 10701 10557 10735 10591
rect 10793 10557 10827 10591
rect 10885 10557 10919 10591
rect 10977 10557 11011 10591
rect 11437 10557 11471 10591
rect 11989 10557 12023 10591
rect 12173 10557 12207 10591
rect 12633 10557 12667 10591
rect 12725 10557 12759 10591
rect 13093 10557 13127 10591
rect 13645 10557 13679 10591
rect 14105 10557 14139 10591
rect 14289 10557 14323 10591
rect 14657 10557 14691 10591
rect 15209 10557 15243 10591
rect 15853 10557 15887 10591
rect 16129 10557 16163 10591
rect 16313 10557 16347 10591
rect 16773 10557 16807 10591
rect 16957 10557 16991 10591
rect 17325 10557 17359 10591
rect 17417 10557 17451 10591
rect 17601 10557 17635 10591
rect 17877 10557 17911 10591
rect 18337 10557 18371 10591
rect 18521 10557 18555 10591
rect 18981 10557 19015 10591
rect 20269 10557 20303 10591
rect 20545 10557 20579 10591
rect 20637 10557 20671 10591
rect 20821 10557 20855 10591
rect 21465 10557 21499 10591
rect 22109 10557 22143 10591
rect 22753 10557 22787 10591
rect 23029 10557 23063 10591
rect 7021 10489 7055 10523
rect 11161 10489 11195 10523
rect 11253 10489 11287 10523
rect 11805 10489 11839 10523
rect 15991 10489 16025 10523
rect 16221 10489 16255 10523
rect 19809 10489 19843 10523
rect 19993 10489 20027 10523
rect 22017 10489 22051 10523
rect 4721 10421 4755 10455
rect 6193 10421 6227 10455
rect 9229 10421 9263 10455
rect 9873 10421 9907 10455
rect 12449 10421 12483 10455
rect 13277 10421 13311 10455
rect 13829 10421 13863 10455
rect 14473 10421 14507 10455
rect 16497 10421 16531 10455
rect 18061 10421 18095 10455
rect 18429 10421 18463 10455
rect 19625 10421 19659 10455
rect 20361 10421 20395 10455
rect 22569 10421 22603 10455
rect 22937 10421 22971 10455
rect 3617 10217 3651 10251
rect 4629 10217 4663 10251
rect 6745 10217 6779 10251
rect 11989 10217 12023 10251
rect 12817 10217 12851 10251
rect 16221 10217 16255 10251
rect 20269 10217 20303 10251
rect 21465 10217 21499 10251
rect 4169 10149 4203 10183
rect 6009 10149 6043 10183
rect 6193 10149 6227 10183
rect 15761 10149 15795 10183
rect 17785 10149 17819 10183
rect 857 10081 891 10115
rect 1124 10081 1158 10115
rect 2329 10081 2363 10115
rect 2605 10081 2639 10115
rect 2789 10081 2823 10115
rect 3157 10081 3191 10115
rect 3985 10081 4019 10115
rect 4445 10081 4479 10115
rect 6469 10081 6503 10115
rect 6929 10081 6963 10115
rect 7205 10081 7239 10115
rect 7389 10081 7423 10115
rect 7941 10081 7975 10115
rect 8033 10081 8067 10115
rect 8217 10081 8251 10115
rect 8493 10081 8527 10115
rect 8677 10081 8711 10115
rect 8769 10081 8803 10115
rect 8861 10081 8895 10115
rect 9229 10081 9263 10115
rect 9689 10081 9723 10115
rect 9873 10081 9907 10115
rect 9965 10081 9999 10115
rect 10057 10081 10091 10115
rect 10517 10081 10551 10115
rect 11805 10081 11839 10115
rect 12265 10081 12299 10115
rect 13001 10081 13035 10115
rect 13093 10081 13127 10115
rect 13277 10081 13311 10115
rect 13369 10081 13403 10115
rect 13645 10081 13679 10115
rect 14657 10081 14691 10115
rect 15669 10081 15703 10115
rect 15945 10081 15979 10115
rect 16129 10081 16163 10115
rect 16313 10081 16347 10115
rect 17693 10081 17727 10115
rect 17877 10081 17911 10115
rect 18061 10081 18095 10115
rect 18153 10081 18187 10115
rect 18337 10081 18371 10115
rect 19165 10081 19199 10115
rect 19349 10081 19383 10115
rect 19625 10081 19659 10115
rect 20637 10081 20671 10115
rect 20913 10081 20947 10115
rect 21649 10081 21683 10115
rect 22477 10081 22511 10115
rect 22753 10081 22787 10115
rect 23029 10081 23063 10115
rect 6653 10013 6687 10047
rect 7665 10013 7699 10047
rect 13185 10013 13219 10047
rect 14749 10013 14783 10047
rect 19073 10013 19107 10047
rect 19257 10013 19291 10047
rect 19533 10013 19567 10047
rect 21281 10013 21315 10047
rect 2513 9945 2547 9979
rect 6285 9945 6319 9979
rect 7849 9945 7883 9979
rect 10333 9945 10367 9979
rect 15025 9945 15059 9979
rect 15853 9945 15887 9979
rect 18337 9945 18371 9979
rect 19809 9945 19843 9979
rect 22845 9945 22879 9979
rect 2237 9877 2271 9911
rect 2973 9877 3007 9911
rect 3433 9877 3467 9911
rect 4353 9877 4387 9911
rect 5825 9877 5859 9911
rect 7205 9877 7239 9911
rect 7757 9877 7791 9911
rect 8217 9877 8251 9911
rect 8401 9877 8435 9911
rect 9137 9877 9171 9911
rect 9413 9877 9447 9911
rect 10701 9877 10735 9911
rect 12081 9877 12115 9911
rect 20085 9877 20119 9911
rect 20269 9877 20303 9911
rect 20729 9877 20763 9911
rect 21649 9877 21683 9911
rect 22293 9877 22327 9911
rect 22661 9877 22695 9911
rect 2375 9673 2409 9707
rect 8493 9673 8527 9707
rect 21741 9673 21775 9707
rect 6377 9605 6411 9639
rect 7021 9605 7055 9639
rect 8125 9605 8159 9639
rect 9873 9605 9907 9639
rect 12449 9605 12483 9639
rect 16497 9605 16531 9639
rect 20913 9605 20947 9639
rect 22201 9605 22235 9639
rect 4353 9537 4387 9571
rect 4997 9537 5031 9571
rect 6101 9537 6135 9571
rect 6929 9537 6963 9571
rect 8861 9537 8895 9571
rect 8953 9537 8987 9571
rect 9045 9537 9079 9571
rect 11621 9537 11655 9571
rect 11989 9537 12023 9571
rect 12817 9537 12851 9571
rect 12909 9537 12943 9571
rect 13645 9537 13679 9571
rect 16405 9537 16439 9571
rect 17509 9537 17543 9571
rect 19533 9537 19567 9571
rect 22845 9537 22879 9571
rect 1041 9469 1075 9503
rect 1409 9469 1443 9503
rect 2145 9469 2179 9503
rect 3525 9469 3559 9503
rect 3617 9469 3651 9503
rect 3709 9469 3743 9503
rect 3893 9469 3927 9503
rect 3985 9469 4019 9503
rect 4169 9469 4203 9503
rect 4445 9469 4479 9503
rect 4905 9469 4939 9503
rect 5089 9469 5123 9503
rect 5457 9469 5491 9503
rect 5641 9469 5675 9503
rect 5733 9469 5767 9503
rect 6009 9469 6043 9503
rect 6653 9469 6687 9503
rect 6837 9469 6871 9503
rect 7448 9469 7482 9503
rect 7665 9469 7699 9503
rect 7941 9469 7975 9503
rect 8401 9469 8435 9503
rect 8585 9469 8619 9503
rect 9137 9469 9171 9503
rect 9597 9469 9631 9503
rect 9689 9469 9723 9503
rect 9965 9469 9999 9503
rect 10425 9469 10459 9503
rect 10609 9469 10643 9503
rect 10701 9469 10735 9503
rect 10793 9469 10827 9503
rect 10977 9469 11011 9503
rect 11161 9469 11195 9503
rect 11253 9469 11287 9503
rect 11437 9469 11471 9503
rect 11529 9469 11563 9503
rect 11816 9469 11850 9503
rect 12541 9469 12575 9503
rect 12725 9469 12759 9503
rect 13093 9469 13127 9503
rect 13829 9469 13863 9503
rect 14105 9469 14139 9503
rect 14289 9469 14323 9503
rect 16681 9469 16715 9503
rect 17233 9469 17267 9503
rect 17325 9469 17359 9503
rect 17601 9469 17635 9503
rect 17693 9469 17727 9503
rect 17877 9469 17911 9503
rect 19257 9469 19291 9503
rect 19441 9469 19475 9503
rect 19809 9469 19843 9503
rect 20637 9469 20671 9503
rect 20821 9469 20855 9503
rect 21097 9469 21131 9503
rect 21557 9469 21591 9503
rect 21649 9469 21683 9503
rect 21833 9469 21867 9503
rect 22109 9469 22143 9503
rect 22385 9469 22419 9503
rect 22477 9469 22511 9503
rect 22661 9469 22695 9503
rect 22753 9469 22787 9503
rect 22937 9469 22971 9503
rect 4077 9401 4111 9435
rect 7757 9401 7791 9435
rect 10149 9401 10183 9435
rect 10333 9401 10367 9435
rect 12081 9401 12115 9435
rect 12265 9401 12299 9435
rect 16865 9401 16899 9435
rect 22569 9401 22603 9435
rect 2053 9333 2087 9367
rect 3249 9333 3283 9367
rect 4813 9333 4847 9367
rect 5273 9333 5307 9367
rect 6837 9333 6871 9367
rect 7389 9333 7423 9367
rect 7573 9333 7607 9367
rect 9321 9333 9355 9367
rect 9413 9333 9447 9367
rect 13277 9333 13311 9367
rect 14013 9333 14047 9367
rect 14197 9333 14231 9367
rect 17049 9333 17083 9367
rect 17785 9333 17819 9367
rect 19349 9333 19383 9367
rect 20453 9333 20487 9367
rect 21373 9333 21407 9367
rect 21925 9333 21959 9367
rect 1133 9129 1167 9163
rect 1593 9129 1627 9163
rect 4353 9129 4387 9163
rect 6285 9129 6319 9163
rect 11345 9129 11379 9163
rect 22017 9129 22051 9163
rect 2145 9061 2179 9095
rect 2697 9061 2731 9095
rect 8769 9061 8803 9095
rect 8953 9061 8987 9095
rect 11161 9061 11195 9095
rect 16129 9061 16163 9095
rect 16313 9061 16347 9095
rect 17969 9061 18003 9095
rect 19165 9061 19199 9095
rect 22477 9061 22511 9095
rect 1317 8993 1351 9027
rect 1777 8993 1811 9027
rect 1961 8993 1995 9027
rect 2329 8993 2363 9027
rect 2605 8993 2639 9027
rect 2789 8993 2823 9027
rect 2973 8993 3007 9027
rect 3065 8993 3099 9027
rect 3341 8993 3375 9027
rect 3985 8993 4019 9027
rect 4445 8993 4479 9027
rect 5825 8993 5859 9027
rect 7205 8993 7239 9027
rect 7477 8993 7511 9027
rect 10977 8993 11011 9027
rect 14105 8993 14139 9027
rect 14197 8993 14231 9027
rect 14473 8993 14507 9027
rect 14749 8993 14783 9027
rect 14841 8993 14875 9027
rect 15117 8993 15151 9027
rect 15209 8993 15243 9027
rect 15485 8993 15519 9027
rect 15669 8993 15703 9027
rect 17785 8993 17819 9027
rect 18265 8993 18299 9027
rect 18429 8993 18463 9027
rect 18521 8993 18555 9027
rect 18613 8993 18647 9027
rect 18909 8993 18943 9027
rect 19073 8993 19107 9027
rect 19257 8993 19291 9027
rect 19809 8993 19843 9027
rect 20085 8993 20119 9027
rect 21465 8993 21499 9027
rect 22201 8993 22235 9027
rect 22661 8993 22695 9027
rect 22753 8993 22787 9027
rect 22937 8993 22971 9027
rect 3249 8925 3283 8959
rect 7849 8925 7883 8959
rect 8125 8925 8159 8959
rect 22845 8925 22879 8959
rect 2421 8857 2455 8891
rect 7389 8857 7423 8891
rect 14381 8857 14415 8891
rect 15393 8857 15427 8891
rect 19901 8857 19935 8891
rect 19993 8857 20027 8891
rect 22293 8857 22327 8891
rect 3617 8789 3651 8823
rect 4169 8789 4203 8823
rect 5917 8789 5951 8823
rect 7021 8789 7055 8823
rect 9137 8789 9171 8823
rect 13921 8789 13955 8823
rect 14565 8789 14599 8823
rect 15025 8789 15059 8823
rect 15853 8789 15887 8823
rect 16497 8789 16531 8823
rect 18153 8789 18187 8823
rect 18797 8789 18831 8823
rect 19441 8789 19475 8823
rect 20269 8789 20303 8823
rect 21281 8789 21315 8823
rect 3525 8585 3559 8619
rect 5273 8585 5307 8619
rect 5733 8585 5767 8619
rect 19809 8585 19843 8619
rect 21189 8585 21223 8619
rect 1869 8517 1903 8551
rect 2605 8517 2639 8551
rect 4077 8517 4111 8551
rect 11989 8517 12023 8551
rect 13645 8517 13679 8551
rect 13921 8517 13955 8551
rect 18153 8517 18187 8551
rect 1593 8449 1627 8483
rect 2145 8449 2179 8483
rect 3709 8449 3743 8483
rect 4537 8449 4571 8483
rect 4813 8449 4847 8483
rect 6561 8449 6595 8483
rect 8401 8449 8435 8483
rect 8677 8449 8711 8483
rect 10609 8449 10643 8483
rect 13829 8449 13863 8483
rect 16405 8449 16439 8483
rect 17233 8449 17267 8483
rect 22477 8449 22511 8483
rect 1501 8381 1535 8415
rect 2237 8381 2271 8415
rect 3433 8381 3467 8415
rect 3801 8381 3835 8415
rect 4445 8381 4479 8415
rect 5181 8381 5215 8415
rect 5457 8381 5491 8415
rect 5549 8381 5583 8415
rect 6009 8381 6043 8415
rect 6193 8381 6227 8415
rect 6285 8381 6319 8415
rect 7941 8381 7975 8415
rect 8217 8381 8251 8415
rect 9321 8381 9355 8415
rect 9505 8381 9539 8415
rect 9597 8381 9631 8415
rect 9689 8381 9723 8415
rect 9873 8381 9907 8415
rect 10333 8381 10367 8415
rect 10425 8381 10459 8415
rect 10701 8381 10735 8415
rect 11713 8381 11747 8415
rect 11805 8381 11839 8415
rect 12081 8381 12115 8415
rect 12449 8381 12483 8415
rect 12633 8381 12667 8415
rect 12725 8381 12759 8415
rect 12817 8381 12851 8415
rect 13001 8381 13035 8415
rect 13553 8381 13587 8415
rect 14105 8381 14139 8415
rect 16037 8381 16071 8415
rect 16221 8381 16255 8415
rect 16313 8381 16347 8415
rect 16589 8381 16623 8415
rect 16865 8381 16899 8415
rect 17049 8381 17083 8415
rect 17141 8381 17175 8415
rect 17417 8381 17451 8415
rect 17877 8381 17911 8415
rect 17969 8381 18003 8415
rect 18245 8381 18279 8415
rect 19993 8381 20027 8415
rect 20269 8381 20303 8415
rect 21005 8381 21039 8415
rect 21373 8381 21407 8415
rect 21465 8381 21499 8415
rect 21925 8381 21959 8415
rect 22109 8381 22143 8415
rect 22201 8381 22235 8415
rect 4077 8313 4111 8347
rect 10149 8313 10183 8347
rect 16773 8313 16807 8347
rect 17601 8313 17635 8347
rect 3709 8245 3743 8279
rect 3893 8245 3927 8279
rect 4997 8245 5031 8279
rect 6101 8245 6135 8279
rect 10057 8245 10091 8279
rect 11529 8245 11563 8279
rect 13185 8245 13219 8279
rect 13829 8245 13863 8279
rect 17693 8245 17727 8279
rect 20085 8245 20119 8279
rect 20821 8245 20855 8279
rect 21649 8245 21683 8279
rect 22017 8245 22051 8279
rect 1961 8041 1995 8075
rect 2329 8041 2363 8075
rect 12357 8041 12391 8075
rect 15485 8041 15519 8075
rect 21481 8041 21515 8075
rect 1685 7973 1719 8007
rect 11989 7973 12023 8007
rect 12173 7973 12207 8007
rect 19165 7973 19199 8007
rect 21281 7973 21315 8007
rect 1225 7905 1259 7939
rect 1869 7905 1903 7939
rect 2145 7905 2179 7939
rect 2513 7905 2547 7939
rect 2697 7905 2731 7939
rect 2789 7905 2823 7939
rect 2881 7905 2915 7939
rect 3065 7905 3099 7939
rect 3157 7905 3191 7939
rect 3617 7905 3651 7939
rect 4629 7905 4663 7939
rect 6193 7905 6227 7939
rect 6377 7905 6411 7939
rect 6469 7905 6503 7939
rect 6653 7905 6687 7939
rect 6745 7905 6779 7939
rect 6929 7905 6963 7939
rect 7297 7905 7331 7939
rect 7573 7905 7607 7939
rect 7849 7905 7883 7939
rect 7941 7905 7975 7939
rect 9137 7905 9171 7939
rect 9229 7905 9263 7939
rect 9873 7905 9907 7939
rect 9965 7905 9999 7939
rect 10241 7905 10275 7939
rect 10333 7905 10367 7939
rect 10517 7905 10551 7939
rect 10701 7905 10735 7939
rect 10977 7905 11011 7939
rect 11161 7905 11195 7939
rect 11253 7905 11287 7939
rect 11529 7905 11563 7939
rect 14289 7905 14323 7939
rect 14657 7905 14691 7939
rect 15669 7905 15703 7939
rect 15761 7905 15795 7939
rect 18153 7905 18187 7939
rect 18521 7905 18555 7939
rect 18705 7905 18739 7939
rect 18981 7905 19015 7939
rect 19257 7905 19291 7939
rect 19533 7905 19567 7939
rect 19717 7905 19751 7939
rect 19809 7905 19843 7939
rect 1317 7837 1351 7871
rect 3525 7837 3559 7871
rect 4721 7837 4755 7871
rect 6561 7837 6595 7871
rect 7021 7837 7055 7871
rect 7113 7837 7147 7871
rect 8861 7837 8895 7871
rect 9505 7837 9539 7871
rect 11345 7837 11379 7871
rect 14565 7837 14599 7871
rect 14933 7837 14967 7871
rect 18337 7837 18371 7871
rect 18429 7837 18463 7871
rect 1501 7769 1535 7803
rect 2881 7769 2915 7803
rect 4997 7769 5031 7803
rect 7665 7769 7699 7803
rect 9321 7769 9355 7803
rect 10149 7769 10183 7803
rect 14473 7769 14507 7803
rect 857 7701 891 7735
rect 3341 7701 3375 7735
rect 3893 7701 3927 7735
rect 6285 7701 6319 7735
rect 7481 7701 7515 7735
rect 8125 7701 8159 7735
rect 9413 7701 9447 7735
rect 9689 7701 9723 7735
rect 11713 7701 11747 7735
rect 14381 7701 14415 7735
rect 14749 7701 14783 7735
rect 14841 7701 14875 7735
rect 15945 7701 15979 7735
rect 17969 7701 18003 7735
rect 18797 7701 18831 7735
rect 19349 7701 19383 7735
rect 21465 7701 21499 7735
rect 21649 7701 21683 7735
rect 1317 7497 1351 7531
rect 2145 7497 2179 7531
rect 7113 7497 7147 7531
rect 7205 7497 7239 7531
rect 21649 7497 21683 7531
rect 6929 7429 6963 7463
rect 9229 7429 9263 7463
rect 11345 7429 11379 7463
rect 16865 7429 16899 7463
rect 18245 7429 18279 7463
rect 21833 7429 21867 7463
rect 22201 7429 22235 7463
rect 1777 7361 1811 7395
rect 2789 7361 2823 7395
rect 3065 7361 3099 7395
rect 3617 7361 3651 7395
rect 5917 7361 5951 7395
rect 7021 7361 7055 7395
rect 7757 7361 7791 7395
rect 9413 7361 9447 7395
rect 11529 7361 11563 7395
rect 13829 7361 13863 7395
rect 17049 7361 17083 7395
rect 19441 7361 19475 7395
rect 19993 7361 20027 7395
rect 20269 7361 20303 7395
rect 22293 7361 22327 7395
rect 1041 7293 1075 7327
rect 1501 7293 1535 7327
rect 1961 7293 1995 7327
rect 3341 7293 3375 7327
rect 4445 7293 4479 7327
rect 4629 7293 4663 7327
rect 5273 7293 5307 7327
rect 5549 7293 5583 7327
rect 6009 7293 6043 7327
rect 6380 7293 6414 7327
rect 6745 7293 6779 7327
rect 6929 7293 6963 7327
rect 7297 7293 7331 7327
rect 7573 7293 7607 7327
rect 7849 7293 7883 7327
rect 8401 7293 8435 7327
rect 8585 7293 8619 7327
rect 8677 7293 8711 7327
rect 8769 7293 8803 7327
rect 9137 7293 9171 7327
rect 10241 7293 10275 7327
rect 11253 7293 11287 7327
rect 13645 7293 13679 7327
rect 13737 7293 13771 7327
rect 13921 7293 13955 7327
rect 14381 7293 14415 7327
rect 14565 7293 14599 7327
rect 14749 7293 14783 7327
rect 15485 7293 15519 7327
rect 16773 7293 16807 7327
rect 18429 7293 18463 7327
rect 19349 7293 19383 7327
rect 19625 7293 19659 7327
rect 19717 7293 19751 7327
rect 21925 7293 21959 7327
rect 14473 7225 14507 7259
rect 21465 7225 21499 7259
rect 21665 7225 21699 7259
rect 22385 7225 22419 7259
rect 1133 7157 1167 7191
rect 4537 7157 4571 7191
rect 5365 7157 5399 7191
rect 5733 7157 5767 7191
rect 6377 7157 6411 7191
rect 6561 7157 6595 7191
rect 7389 7157 7423 7191
rect 9045 7157 9079 7191
rect 9413 7157 9447 7191
rect 10425 7157 10459 7191
rect 11529 7157 11563 7191
rect 14105 7157 14139 7191
rect 14197 7157 14231 7191
rect 15669 7157 15703 7191
rect 17049 7157 17083 7191
rect 19901 7157 19935 7191
rect 22017 7157 22051 7191
rect 1685 6953 1719 6987
rect 6285 6953 6319 6987
rect 9137 6953 9171 6987
rect 13461 6953 13495 6987
rect 16589 6953 16623 6987
rect 5089 6885 5123 6919
rect 1225 6817 1259 6851
rect 1685 6817 1719 6851
rect 1869 6817 1903 6851
rect 1961 6817 1995 6851
rect 2145 6817 2179 6851
rect 2329 6817 2363 6851
rect 2513 6817 2547 6851
rect 2789 6817 2823 6851
rect 3525 6817 3559 6851
rect 3709 6817 3743 6851
rect 4169 6817 4203 6851
rect 4261 6817 4295 6851
rect 4445 6817 4479 6851
rect 4813 6817 4847 6851
rect 5365 6817 5399 6851
rect 5549 6817 5583 6851
rect 5641 6817 5675 6851
rect 6344 6817 6378 6851
rect 8309 6817 8343 6851
rect 8401 6817 8435 6851
rect 9196 6817 9230 6851
rect 9597 6817 9631 6851
rect 9781 6817 9815 6851
rect 9873 6817 9907 6851
rect 10149 6817 10183 6851
rect 10425 6817 10459 6851
rect 10609 6817 10643 6851
rect 10793 6817 10827 6851
rect 10977 6817 11011 6851
rect 11161 6817 11195 6851
rect 11253 6817 11287 6851
rect 11529 6817 11563 6851
rect 11805 6817 11839 6851
rect 11989 6817 12023 6851
rect 12173 6817 12207 6851
rect 12449 6817 12483 6851
rect 12633 6817 12667 6851
rect 13001 6817 13035 6851
rect 13402 6817 13436 6851
rect 13829 6817 13863 6851
rect 14197 6817 14231 6851
rect 14381 6817 14415 6851
rect 14657 6817 14691 6851
rect 15209 6817 15243 6851
rect 15301 6817 15335 6851
rect 15393 6817 15427 6851
rect 16497 6817 16531 6851
rect 17049 6817 17083 6851
rect 17325 6817 17359 6851
rect 17417 6817 17451 6851
rect 17509 6817 17543 6851
rect 18245 6817 18279 6851
rect 18337 6817 18371 6851
rect 20039 6817 20073 6851
rect 20453 6817 20487 6851
rect 20545 6817 20579 6851
rect 20637 6817 20671 6851
rect 21465 6817 21499 6851
rect 21557 6817 21591 6851
rect 21833 6817 21867 6851
rect 1133 6749 1167 6783
rect 2053 6749 2087 6783
rect 2881 6749 2915 6783
rect 5089 6749 5123 6783
rect 5825 6749 5859 6783
rect 7113 6749 7147 6783
rect 7389 6749 7423 6783
rect 8677 6749 8711 6783
rect 8769 6749 8803 6783
rect 9965 6749 9999 6783
rect 11345 6749 11379 6783
rect 12725 6749 12759 6783
rect 12817 6749 12851 6783
rect 13921 6749 13955 6783
rect 14749 6749 14783 6783
rect 14933 6749 14967 6783
rect 15025 6749 15059 6783
rect 16773 6749 16807 6783
rect 17233 6749 17267 6783
rect 17693 6749 17727 6783
rect 18521 6749 18555 6783
rect 19809 6749 19843 6783
rect 20177 6749 20211 6783
rect 20361 6749 20395 6783
rect 20821 6749 20855 6783
rect 21281 6749 21315 6783
rect 1593 6681 1627 6715
rect 2513 6681 2547 6715
rect 3157 6681 3191 6715
rect 6469 6681 6503 6715
rect 13277 6681 13311 6715
rect 14841 6681 14875 6715
rect 15117 6681 15151 6715
rect 3893 6613 3927 6647
rect 4629 6613 4663 6647
rect 4905 6613 4939 6647
rect 5181 6613 5215 6647
rect 5917 6613 5951 6647
rect 8079 6613 8113 6647
rect 8585 6613 8619 6647
rect 9321 6613 9355 6647
rect 10333 6613 10367 6647
rect 11713 6613 11747 6647
rect 13185 6613 13219 6647
rect 14381 6613 14415 6647
rect 14565 6613 14599 6647
rect 15577 6613 15611 6647
rect 16129 6613 16163 6647
rect 18429 6613 18463 6647
rect 20269 6613 20303 6647
rect 20729 6613 20763 6647
rect 21741 6613 21775 6647
rect 5641 6409 5675 6443
rect 5825 6409 5859 6443
rect 6469 6409 6503 6443
rect 9597 6409 9631 6443
rect 10885 6409 10919 6443
rect 12173 6409 12207 6443
rect 14105 6409 14139 6443
rect 14933 6409 14967 6443
rect 19809 6409 19843 6443
rect 20085 6409 20119 6443
rect 21005 6409 21039 6443
rect 5273 6341 5307 6375
rect 7573 6341 7607 6375
rect 14473 6341 14507 6375
rect 16773 6341 16807 6375
rect 21833 6341 21867 6375
rect 2973 6273 3007 6307
rect 3801 6273 3835 6307
rect 4077 6273 4111 6307
rect 5733 6273 5767 6307
rect 6193 6273 6227 6307
rect 7297 6273 7331 6307
rect 12265 6273 12299 6307
rect 14289 6273 14323 6307
rect 16129 6273 16163 6307
rect 16221 6273 16255 6307
rect 16405 6273 16439 6307
rect 17417 6273 17451 6307
rect 17877 6273 17911 6307
rect 19165 6273 19199 6307
rect 19257 6273 19291 6307
rect 22385 6273 22419 6307
rect 1869 6205 1903 6239
rect 2053 6205 2087 6239
rect 2329 6205 2363 6239
rect 2881 6205 2915 6239
rect 3065 6205 3099 6239
rect 3617 6205 3651 6239
rect 3893 6205 3927 6239
rect 4169 6205 4203 6239
rect 4629 6205 4663 6239
rect 4813 6205 4847 6239
rect 5457 6205 5491 6239
rect 6009 6205 6043 6239
rect 6101 6205 6135 6239
rect 6285 6205 6319 6239
rect 6653 6205 6687 6239
rect 6929 6205 6963 6239
rect 7205 6205 7239 6239
rect 8585 6205 8619 6239
rect 8677 6205 8711 6239
rect 8769 6205 8803 6239
rect 8953 6205 8987 6239
rect 9045 6205 9079 6239
rect 9229 6205 9263 6239
rect 9413 6205 9447 6239
rect 11069 6205 11103 6239
rect 11746 6205 11780 6239
rect 13921 6205 13955 6239
rect 14197 6205 14231 6239
rect 14381 6205 14415 6239
rect 14657 6205 14691 6239
rect 15209 6205 15243 6239
rect 15301 6205 15335 6239
rect 15393 6205 15427 6239
rect 15577 6205 15611 6239
rect 15669 6205 15703 6239
rect 15853 6205 15887 6239
rect 16313 6205 16347 6239
rect 19809 6205 19843 6239
rect 19993 6205 20027 6239
rect 20269 6205 20303 6239
rect 20913 6205 20947 6239
rect 21189 6205 21223 6239
rect 21281 6205 21315 6239
rect 3433 6137 3467 6171
rect 4721 6137 4755 6171
rect 15761 6137 15795 6171
rect 17233 6137 17267 6171
rect 18153 6137 18187 6171
rect 1961 6069 1995 6103
rect 2145 6069 2179 6103
rect 4537 6069 4571 6103
rect 6837 6069 6871 6103
rect 8401 6069 8435 6103
rect 11621 6069 11655 6103
rect 11805 6069 11839 6103
rect 15945 6069 15979 6103
rect 17141 6069 17175 6103
rect 18061 6069 18095 6103
rect 18521 6069 18555 6103
rect 18705 6069 18739 6103
rect 19073 6069 19107 6103
rect 21465 6069 21499 6103
rect 22201 6069 22235 6103
rect 22293 6069 22327 6103
rect 2697 5865 2731 5899
rect 3479 5865 3513 5899
rect 4445 5865 4479 5899
rect 8401 5865 8435 5899
rect 13369 5865 13403 5899
rect 13921 5865 13955 5899
rect 15577 5865 15611 5899
rect 22385 5865 22419 5899
rect 9045 5797 9079 5831
rect 14933 5797 14967 5831
rect 16865 5797 16899 5831
rect 22477 5797 22511 5831
rect 1041 5729 1075 5763
rect 1501 5729 1535 5763
rect 1685 5729 1719 5763
rect 1961 5729 1995 5763
rect 2329 5729 2363 5763
rect 3709 5729 3743 5763
rect 3801 5729 3835 5763
rect 4169 5729 4203 5763
rect 4353 5729 4387 5763
rect 4445 5729 4479 5763
rect 4629 5729 4663 5763
rect 5181 5729 5215 5763
rect 5825 5729 5859 5763
rect 6285 5729 6319 5763
rect 6837 5729 6871 5763
rect 8033 5729 8067 5763
rect 8217 5729 8251 5763
rect 8493 5729 8527 5763
rect 8953 5729 8987 5763
rect 9137 5729 9171 5763
rect 9413 5729 9447 5763
rect 9505 5729 9539 5763
rect 9689 5729 9723 5763
rect 9781 5729 9815 5763
rect 9965 5729 9999 5763
rect 10425 5729 10459 5763
rect 11161 5729 11195 5763
rect 11437 5729 11471 5763
rect 11529 5729 11563 5763
rect 11989 5729 12023 5763
rect 12081 5729 12115 5763
rect 12265 5729 12299 5763
rect 12909 5729 12943 5763
rect 13001 5729 13035 5763
rect 13553 5729 13587 5763
rect 14105 5729 14139 5763
rect 14381 5729 14415 5763
rect 14473 5729 14507 5763
rect 15117 5729 15151 5763
rect 15393 5729 15427 5763
rect 17049 5729 17083 5763
rect 17785 5729 17819 5763
rect 17969 5729 18003 5763
rect 18061 5729 18095 5763
rect 18521 5729 18555 5763
rect 18613 5729 18647 5763
rect 19165 5729 19199 5763
rect 19349 5729 19383 5763
rect 19441 5729 19475 5763
rect 19533 5729 19567 5763
rect 20637 5729 20671 5763
rect 20729 5729 20763 5763
rect 20913 5729 20947 5763
rect 949 5661 983 5695
rect 1869 5661 1903 5695
rect 2421 5661 2455 5695
rect 5089 5661 5123 5695
rect 6561 5661 6595 5695
rect 6745 5661 6779 5695
rect 7205 5661 7239 5695
rect 7941 5661 7975 5695
rect 8125 5661 8159 5695
rect 8585 5661 8619 5695
rect 10057 5661 10091 5695
rect 10517 5661 10551 5695
rect 13185 5661 13219 5695
rect 19717 5661 19751 5695
rect 20361 5661 20395 5695
rect 22569 5661 22603 5695
rect 1409 5593 1443 5627
rect 5549 5593 5583 5627
rect 6009 5593 6043 5627
rect 9229 5593 9263 5627
rect 10333 5593 10367 5627
rect 11253 5593 11287 5627
rect 11805 5593 11839 5627
rect 12173 5593 12207 5627
rect 12541 5593 12575 5627
rect 19257 5593 19291 5627
rect 3985 5525 4019 5559
rect 4261 5525 4295 5559
rect 6377 5525 6411 5559
rect 6469 5525 6503 5559
rect 8585 5525 8619 5559
rect 8861 5525 8895 5559
rect 9965 5525 9999 5559
rect 10425 5525 10459 5559
rect 10793 5525 10827 5559
rect 11713 5525 11747 5559
rect 14197 5525 14231 5559
rect 14657 5525 14691 5559
rect 15301 5525 15335 5559
rect 17233 5525 17267 5559
rect 17601 5525 17635 5559
rect 18521 5525 18555 5559
rect 18889 5525 18923 5559
rect 19625 5525 19659 5559
rect 20821 5525 20855 5559
rect 22017 5525 22051 5559
rect 1593 5321 1627 5355
rect 1961 5321 1995 5355
rect 3801 5321 3835 5355
rect 8585 5321 8619 5355
rect 10333 5321 10367 5355
rect 10425 5321 10459 5355
rect 11805 5321 11839 5355
rect 11897 5321 11931 5355
rect 12449 5321 12483 5355
rect 12817 5321 12851 5355
rect 17049 5321 17083 5355
rect 19625 5321 19659 5355
rect 20453 5321 20487 5355
rect 20545 5321 20579 5355
rect 21833 5321 21867 5355
rect 5917 5253 5951 5287
rect 6285 5253 6319 5287
rect 8217 5253 8251 5287
rect 4169 5185 4203 5219
rect 7389 5185 7423 5219
rect 9137 5185 9171 5219
rect 9781 5185 9815 5219
rect 10977 5185 11011 5219
rect 14105 5185 14139 5219
rect 15577 5185 15611 5219
rect 16681 5185 16715 5219
rect 16773 5185 16807 5219
rect 17509 5185 17543 5219
rect 19073 5185 19107 5219
rect 21925 5185 21959 5219
rect 1225 5117 1259 5151
rect 1409 5117 1443 5151
rect 1501 5117 1535 5151
rect 1685 5117 1719 5151
rect 2145 5117 2179 5151
rect 2881 5117 2915 5151
rect 3893 5117 3927 5151
rect 4997 5117 5031 5151
rect 5273 5117 5307 5151
rect 5457 5117 5491 5151
rect 5917 5117 5951 5151
rect 6193 5117 6227 5151
rect 6653 5117 6687 5151
rect 6745 5117 6779 5151
rect 6929 5117 6963 5151
rect 7021 5117 7055 5151
rect 7113 5117 7147 5151
rect 7573 5117 7607 5151
rect 7757 5117 7791 5151
rect 7849 5117 7883 5151
rect 7941 5117 7975 5151
rect 9045 5117 9079 5151
rect 10793 5117 10827 5151
rect 11253 5117 11287 5151
rect 11345 5117 11379 5151
rect 11529 5117 11563 5151
rect 11621 5117 11655 5151
rect 12081 5117 12115 5151
rect 12357 5117 12391 5151
rect 12633 5117 12667 5151
rect 12725 5117 12759 5151
rect 12909 5117 12943 5151
rect 14013 5117 14047 5151
rect 14565 5117 14599 5151
rect 14841 5117 14875 5151
rect 15761 5117 15795 5151
rect 16497 5117 16531 5151
rect 17233 5117 17267 5151
rect 17417 5117 17451 5151
rect 17601 5117 17635 5151
rect 17785 5117 17819 5151
rect 18797 5117 18831 5151
rect 18889 5117 18923 5151
rect 18981 5117 19015 5151
rect 19533 5117 19567 5151
rect 19809 5117 19843 5151
rect 20269 5117 20303 5151
rect 20729 5117 20763 5151
rect 21189 5117 21223 5151
rect 21557 5117 21591 5151
rect 2329 5049 2363 5083
rect 3433 5049 3467 5083
rect 3617 5049 3651 5083
rect 4813 5049 4847 5083
rect 6469 5049 6503 5083
rect 8953 5049 8987 5083
rect 9873 5049 9907 5083
rect 10885 5049 10919 5083
rect 16313 5049 16347 5083
rect 20085 5049 20119 5083
rect 20913 5049 20947 5083
rect 21649 5049 21683 5083
rect 22017 5049 22051 5083
rect 1317 4981 1351 5015
rect 2697 4981 2731 5015
rect 5181 4981 5215 5015
rect 5365 4981 5399 5015
rect 6101 4981 6135 5015
rect 9965 4981 9999 5015
rect 12173 4981 12207 5015
rect 13553 4981 13587 5015
rect 13921 4981 13955 5015
rect 14381 4981 14415 5015
rect 14657 4981 14691 5015
rect 15669 4981 15703 5015
rect 16129 4981 16163 5015
rect 19257 4981 19291 5015
rect 19349 4981 19383 5015
rect 19993 4981 20027 5015
rect 21005 4981 21039 5015
rect 1133 4777 1167 4811
rect 2421 4777 2455 4811
rect 2789 4777 2823 4811
rect 3433 4777 3467 4811
rect 3893 4777 3927 4811
rect 4353 4777 4387 4811
rect 4997 4777 5031 4811
rect 5641 4777 5675 4811
rect 6745 4777 6779 4811
rect 9229 4777 9263 4811
rect 9321 4777 9355 4811
rect 10149 4777 10183 4811
rect 14473 4777 14507 4811
rect 14565 4777 14599 4811
rect 18337 4777 18371 4811
rect 20361 4777 20395 4811
rect 21005 4777 21039 4811
rect 3157 4709 3191 4743
rect 4629 4709 4663 4743
rect 7541 4709 7575 4743
rect 7757 4709 7791 4743
rect 10057 4709 10091 4743
rect 12541 4709 12575 4743
rect 857 4641 891 4675
rect 1041 4641 1075 4675
rect 1317 4641 1351 4675
rect 1409 4641 1443 4675
rect 1869 4641 1903 4675
rect 2053 4641 2087 4675
rect 2145 4641 2179 4675
rect 2329 4641 2363 4675
rect 2605 4641 2639 4675
rect 2881 4641 2915 4675
rect 3341 4641 3375 4675
rect 3617 4641 3651 4675
rect 3709 4641 3743 4675
rect 4077 4641 4111 4675
rect 4169 4641 4203 4675
rect 4813 4641 4847 4675
rect 5273 4641 5307 4675
rect 5825 4641 5859 4675
rect 7113 4641 7147 4675
rect 8217 4641 8251 4675
rect 8585 4641 8619 4675
rect 11805 4641 11839 4675
rect 12081 4641 12115 4675
rect 12265 4641 12299 4675
rect 12357 4641 12391 4675
rect 13001 4641 13035 4675
rect 13461 4641 13495 4675
rect 15117 4641 15151 4675
rect 16129 4641 16163 4675
rect 17233 4641 17267 4675
rect 17877 4641 17911 4675
rect 18153 4641 18187 4675
rect 18337 4641 18371 4675
rect 18429 4641 18463 4675
rect 18521 4641 18555 4675
rect 18705 4641 18739 4675
rect 19165 4641 19199 4675
rect 19717 4641 19751 4675
rect 19901 4641 19935 4675
rect 20545 4641 20579 4675
rect 20821 4641 20855 4675
rect 20913 4641 20947 4675
rect 21097 4641 21131 4675
rect 21281 4641 21315 4675
rect 21373 4641 21407 4675
rect 21557 4641 21591 4675
rect 21649 4641 21683 4675
rect 21925 4641 21959 4675
rect 22109 4641 22143 4675
rect 22293 4641 22327 4675
rect 22477 4641 22511 4675
rect 949 4573 983 4607
rect 1133 4573 1167 4607
rect 4353 4573 4387 4607
rect 5365 4573 5399 4607
rect 6101 4573 6135 4607
rect 6929 4573 6963 4607
rect 7021 4573 7055 4607
rect 7205 4573 7239 4607
rect 9505 4573 9539 4607
rect 10241 4573 10275 4607
rect 12725 4573 12759 4607
rect 13093 4573 13127 4607
rect 13737 4573 13771 4607
rect 14749 4573 14783 4607
rect 16405 4573 16439 4607
rect 17325 4573 17359 4607
rect 17417 4573 17451 4607
rect 17509 4573 17543 4607
rect 18797 4573 18831 4607
rect 19073 4573 19107 4607
rect 22017 4573 22051 4607
rect 1685 4505 1719 4539
rect 7389 4505 7423 4539
rect 8861 4505 8895 4539
rect 14105 4505 14139 4539
rect 16681 4505 16715 4539
rect 19717 4505 19751 4539
rect 20637 4505 20671 4539
rect 2973 4437 3007 4471
rect 7573 4437 7607 4471
rect 8585 4437 8619 4471
rect 8769 4437 8803 4471
rect 9689 4437 9723 4471
rect 11621 4437 11655 4471
rect 13001 4437 13035 4471
rect 13369 4437 13403 4471
rect 13829 4437 13863 4471
rect 14013 4437 14047 4471
rect 14933 4437 14967 4471
rect 16221 4437 16255 4471
rect 17049 4437 17083 4471
rect 17693 4437 17727 4471
rect 18797 4437 18831 4471
rect 21833 4437 21867 4471
rect 22477 4437 22511 4471
rect 2329 4233 2363 4267
rect 4997 4233 5031 4267
rect 5365 4233 5399 4267
rect 6653 4233 6687 4267
rect 7573 4233 7607 4267
rect 7757 4233 7791 4267
rect 8033 4233 8067 4267
rect 8401 4233 8435 4267
rect 10425 4233 10459 4267
rect 12541 4233 12575 4267
rect 13185 4233 13219 4267
rect 1777 4165 1811 4199
rect 4261 4165 4295 4199
rect 6377 4165 6411 4199
rect 10977 4165 11011 4199
rect 22569 4165 22603 4199
rect 1501 4097 1535 4131
rect 1961 4097 1995 4131
rect 2605 4097 2639 4131
rect 3985 4097 4019 4131
rect 4813 4097 4847 4131
rect 5733 4097 5767 4131
rect 5917 4097 5951 4131
rect 7481 4097 7515 4131
rect 11621 4097 11655 4131
rect 11989 4097 12023 4131
rect 12265 4097 12299 4131
rect 14657 4097 14691 4131
rect 14749 4097 14783 4131
rect 15209 4097 15243 4131
rect 15301 4097 15335 4131
rect 15393 4097 15427 4131
rect 16221 4097 16255 4131
rect 16313 4097 16347 4131
rect 16405 4097 16439 4131
rect 16589 4097 16623 4131
rect 21097 4097 21131 4131
rect 1409 4029 1443 4063
rect 2421 4029 2455 4063
rect 2697 4029 2731 4063
rect 3893 4029 3927 4063
rect 4353 4029 4387 4063
rect 4537 4029 4571 4063
rect 4721 4029 4755 4063
rect 4905 4029 4939 4063
rect 5181 4029 5215 4063
rect 5273 4029 5307 4063
rect 5549 4029 5583 4063
rect 6009 4029 6043 4063
rect 6837 4029 6871 4063
rect 7113 4029 7147 4063
rect 7205 4029 7239 4063
rect 8401 4029 8435 4063
rect 8585 4029 8619 4063
rect 9321 4029 9355 4063
rect 10057 4029 10091 4063
rect 10701 4029 10735 4063
rect 11161 4029 11195 4063
rect 11529 4029 11563 4063
rect 11713 4029 11747 4063
rect 12081 4029 12115 4063
rect 12173 4029 12207 4063
rect 12449 4029 12483 4063
rect 12725 4029 12759 4063
rect 12817 4029 12851 4063
rect 13001 4029 13035 4063
rect 13369 4029 13403 4063
rect 13829 4029 13863 4063
rect 13921 4029 13955 4063
rect 14105 4029 14139 4063
rect 14473 4029 14507 4063
rect 14565 4029 14599 4063
rect 15485 4029 15519 4063
rect 15853 4029 15887 4063
rect 16129 4029 16163 4063
rect 19165 4029 19199 4063
rect 19349 4029 19383 4063
rect 19809 4029 19843 4063
rect 19993 4029 20027 4063
rect 20361 4029 20395 4063
rect 20453 4029 20487 4063
rect 20637 4029 20671 4063
rect 20729 4029 20763 4063
rect 21189 4029 21223 4063
rect 21343 4029 21377 4063
rect 21833 4029 21867 4063
rect 22017 4029 22051 4063
rect 22109 4029 22143 4063
rect 22293 4029 22327 4063
rect 22385 4029 22419 4063
rect 22753 4029 22787 4063
rect 8001 3961 8035 3995
rect 8217 3961 8251 3995
rect 9597 3961 9631 3995
rect 9781 3961 9815 3995
rect 10241 3961 10275 3995
rect 19901 3961 19935 3995
rect 21557 3961 21591 3995
rect 3065 3893 3099 3927
rect 4353 3893 4387 3927
rect 7021 3893 7055 3927
rect 7849 3893 7883 3927
rect 8769 3893 8803 3927
rect 9413 3893 9447 3927
rect 9965 3893 9999 3927
rect 10517 3893 10551 3927
rect 11805 3893 11839 3927
rect 13001 3893 13035 3927
rect 13645 3893 13679 3927
rect 14013 3893 14047 3927
rect 14933 3893 14967 3927
rect 15025 3893 15059 3927
rect 15669 3893 15703 3927
rect 19257 3893 19291 3927
rect 20177 3893 20211 3927
rect 20545 3893 20579 3927
rect 20913 3893 20947 3927
rect 21649 3893 21683 3927
rect 22845 3893 22879 3927
rect 1685 3689 1719 3723
rect 3525 3689 3559 3723
rect 7573 3689 7607 3723
rect 12817 3689 12851 3723
rect 14657 3689 14691 3723
rect 1225 3621 1259 3655
rect 6101 3621 6135 3655
rect 6469 3621 6503 3655
rect 7205 3621 7239 3655
rect 12265 3621 12299 3655
rect 15025 3621 15059 3655
rect 3157 3553 3191 3587
rect 4537 3553 4571 3587
rect 4721 3553 4755 3587
rect 6285 3553 6319 3587
rect 7113 3553 7147 3587
rect 7389 3553 7423 3587
rect 8217 3553 8251 3587
rect 8401 3553 8435 3587
rect 8493 3553 8527 3587
rect 8677 3553 8711 3587
rect 8953 3553 8987 3587
rect 9045 3553 9079 3587
rect 9137 3553 9171 3587
rect 9229 3553 9263 3587
rect 9413 3553 9447 3587
rect 9597 3553 9631 3587
rect 9965 3553 9999 3587
rect 10425 3553 10459 3587
rect 10517 3553 10551 3587
rect 11253 3553 11287 3587
rect 11345 3553 11379 3587
rect 11989 3553 12023 3587
rect 12081 3553 12115 3587
rect 12357 3553 12391 3587
rect 12909 3553 12943 3587
rect 13829 3553 13863 3587
rect 14105 3553 14139 3587
rect 14841 3553 14875 3587
rect 16313 3553 16347 3587
rect 16405 3553 16439 3587
rect 16589 3553 16623 3587
rect 16681 3553 16715 3587
rect 17233 3553 17267 3587
rect 17417 3553 17451 3587
rect 17693 3553 17727 3587
rect 17877 3553 17911 3587
rect 18613 3553 18647 3587
rect 19165 3553 19199 3587
rect 19533 3553 19567 3587
rect 19717 3553 19751 3587
rect 19901 3553 19935 3587
rect 20269 3553 20303 3587
rect 20821 3553 20855 3587
rect 21373 3553 21407 3587
rect 21649 3553 21683 3587
rect 22109 3553 22143 3587
rect 22201 3553 22235 3587
rect 22661 3553 22695 3587
rect 3065 3485 3099 3519
rect 9689 3485 9723 3519
rect 9781 3485 9815 3519
rect 10609 3485 10643 3519
rect 10701 3485 10735 3519
rect 11161 3485 11195 3519
rect 11437 3485 11471 3519
rect 12633 3485 12667 3519
rect 13921 3485 13955 3519
rect 14013 3485 14047 3519
rect 17325 3485 17359 3519
rect 18889 3485 18923 3519
rect 19349 3485 19383 3519
rect 19441 3485 19475 3519
rect 20545 3485 20579 3519
rect 21097 3485 21131 3519
rect 1501 3417 1535 3451
rect 8585 3417 8619 3451
rect 10241 3417 10275 3451
rect 12541 3417 12575 3451
rect 18981 3417 19015 3451
rect 20637 3417 20671 3451
rect 21005 3417 21039 3451
rect 21925 3417 21959 3451
rect 4629 3349 4663 3383
rect 8309 3349 8343 3383
rect 8769 3349 8803 3383
rect 10149 3349 10183 3383
rect 10977 3349 11011 3383
rect 12265 3349 12299 3383
rect 12449 3349 12483 3383
rect 13645 3349 13679 3383
rect 16129 3349 16163 3383
rect 17877 3349 17911 3383
rect 18429 3349 18463 3383
rect 18797 3349 18831 3383
rect 20085 3349 20119 3383
rect 20453 3349 20487 3383
rect 21465 3349 21499 3383
rect 21833 3349 21867 3383
rect 22293 3349 22327 3383
rect 22753 3349 22787 3383
rect 5273 3145 5307 3179
rect 7021 3145 7055 3179
rect 10149 3145 10183 3179
rect 10793 3145 10827 3179
rect 19809 3145 19843 3179
rect 20545 3145 20579 3179
rect 21097 3145 21131 3179
rect 2329 3077 2363 3111
rect 3801 3077 3835 3111
rect 4537 3077 4571 3111
rect 5549 3077 5583 3111
rect 12817 3077 12851 3111
rect 13553 3077 13587 3111
rect 17325 3077 17359 3111
rect 17417 3077 17451 3111
rect 17785 3077 17819 3111
rect 22201 3077 22235 3111
rect 22477 3077 22511 3111
rect 1225 3009 1259 3043
rect 1869 3009 1903 3043
rect 3341 3009 3375 3043
rect 4629 3009 4663 3043
rect 4997 3009 5031 3043
rect 6193 3009 6227 3043
rect 8677 3009 8711 3043
rect 8769 3009 8803 3043
rect 8861 3009 8895 3043
rect 9321 3009 9355 3043
rect 9413 3009 9447 3043
rect 9505 3009 9539 3043
rect 20637 3009 20671 3043
rect 21189 3009 21223 3043
rect 1317 2941 1351 2975
rect 1961 2941 1995 2975
rect 3433 2941 3467 2975
rect 4353 2941 4387 2975
rect 4905 2941 4939 2975
rect 5365 2941 5399 2975
rect 6009 2941 6043 2975
rect 7205 2941 7239 2975
rect 7481 2941 7515 2975
rect 8953 2941 8987 2975
rect 9597 2941 9631 2975
rect 9965 2941 9999 2975
rect 10149 2941 10183 2975
rect 10609 2941 10643 2975
rect 10701 2941 10735 2975
rect 10885 2941 10919 2975
rect 11161 2941 11195 2975
rect 11345 2941 11379 2975
rect 11529 2941 11563 2975
rect 11621 2941 11655 2975
rect 12081 2941 12115 2975
rect 12541 2941 12575 2975
rect 13737 2941 13771 2975
rect 13829 2941 13863 2975
rect 14013 2941 14047 2975
rect 14105 2941 14139 2975
rect 15117 2941 15151 2975
rect 16497 2941 16531 2975
rect 17233 2941 17267 2975
rect 17509 2941 17543 2975
rect 17969 2941 18003 2975
rect 18061 2941 18095 2975
rect 19165 2941 19199 2975
rect 19349 2941 19383 2975
rect 19993 2941 20027 2975
rect 20361 2941 20395 2975
rect 20913 2941 20947 2975
rect 21281 2941 21315 2975
rect 21373 2941 21407 2975
rect 21557 2941 21591 2975
rect 21833 2941 21867 2975
rect 22109 2941 22143 2975
rect 22661 2941 22695 2975
rect 22753 2941 22787 2975
rect 12817 2873 12851 2907
rect 13553 2873 13587 2907
rect 17785 2873 17819 2907
rect 19257 2873 19291 2907
rect 1685 2805 1719 2839
rect 4169 2805 4203 2839
rect 5825 2805 5859 2839
rect 7389 2805 7423 2839
rect 8493 2805 8527 2839
rect 9137 2805 9171 2839
rect 10517 2805 10551 2839
rect 11897 2805 11931 2839
rect 12633 2805 12667 2839
rect 15025 2805 15059 2839
rect 16405 2805 16439 2839
rect 17049 2805 17083 2839
rect 20177 2805 20211 2839
rect 20729 2805 20763 2839
rect 21741 2805 21775 2839
rect 22017 2805 22051 2839
rect 22937 2805 22971 2839
rect 2973 2601 3007 2635
rect 4813 2601 4847 2635
rect 5549 2601 5583 2635
rect 6561 2601 6595 2635
rect 7573 2601 7607 2635
rect 8033 2601 8067 2635
rect 8401 2601 8435 2635
rect 8861 2601 8895 2635
rect 11161 2601 11195 2635
rect 11529 2601 11563 2635
rect 12265 2601 12299 2635
rect 13277 2601 13311 2635
rect 16589 2601 16623 2635
rect 19073 2601 19107 2635
rect 6653 2533 6687 2567
rect 6837 2533 6871 2567
rect 9413 2533 9447 2567
rect 10609 2533 10643 2567
rect 11989 2533 12023 2567
rect 12449 2533 12483 2567
rect 14749 2533 14783 2567
rect 15301 2533 15335 2567
rect 16129 2533 16163 2567
rect 17325 2533 17359 2567
rect 18521 2533 18555 2567
rect 18889 2533 18923 2567
rect 21557 2533 21591 2567
rect 21925 2533 21959 2567
rect 22753 2533 22787 2567
rect 2881 2465 2915 2499
rect 3157 2465 3191 2499
rect 3433 2465 3467 2499
rect 3709 2465 3743 2499
rect 4445 2465 4479 2499
rect 5181 2465 5215 2499
rect 5365 2465 5399 2499
rect 5641 2465 5675 2499
rect 6193 2465 6227 2499
rect 7205 2465 7239 2499
rect 7389 2465 7423 2499
rect 7849 2465 7883 2499
rect 8125 2465 8159 2499
rect 8217 2465 8251 2499
rect 8493 2465 8527 2499
rect 8769 2465 8803 2499
rect 9045 2465 9079 2499
rect 9229 2465 9263 2499
rect 9505 2465 9539 2499
rect 9781 2465 9815 2499
rect 10057 2465 10091 2499
rect 10241 2465 10275 2499
rect 10333 2465 10367 2499
rect 10425 2465 10459 2499
rect 10977 2465 11011 2499
rect 11345 2465 11379 2499
rect 11621 2465 11655 2499
rect 11713 2465 11747 2499
rect 11805 2465 11839 2499
rect 12081 2465 12115 2499
rect 12357 2465 12391 2499
rect 12633 2465 12667 2499
rect 12909 2465 12943 2499
rect 13001 2465 13035 2499
rect 13461 2465 13495 2499
rect 13553 2465 13587 2499
rect 13737 2465 13771 2499
rect 13829 2465 13863 2499
rect 13921 2465 13955 2499
rect 14657 2465 14691 2499
rect 14933 2465 14967 2499
rect 15025 2465 15059 2499
rect 15117 2465 15151 2499
rect 15393 2465 15427 2499
rect 15577 2465 15611 2499
rect 16313 2465 16347 2499
rect 16405 2465 16439 2499
rect 16497 2465 16531 2499
rect 16773 2465 16807 2499
rect 17049 2465 17083 2499
rect 17141 2465 17175 2499
rect 18705 2465 18739 2499
rect 18797 2465 18831 2499
rect 19165 2465 19199 2499
rect 20269 2465 20303 2499
rect 20637 2465 20671 2499
rect 20729 2465 20763 2499
rect 21281 2465 21315 2499
rect 21373 2465 21407 2499
rect 21649 2465 21683 2499
rect 21741 2465 21775 2499
rect 22201 2465 22235 2499
rect 22293 2465 22327 2499
rect 22477 2465 22511 2499
rect 22569 2465 22603 2499
rect 22845 2465 22879 2499
rect 3617 2397 3651 2431
rect 4169 2397 4203 2431
rect 4353 2397 4387 2431
rect 6101 2397 6135 2431
rect 7021 2397 7055 2431
rect 7113 2397 7147 2431
rect 3157 2329 3191 2363
rect 9229 2329 9263 2363
rect 11989 2329 12023 2363
rect 13185 2329 13219 2363
rect 14933 2329 14967 2363
rect 15301 2329 15335 2363
rect 15577 2329 15611 2363
rect 20085 2329 20119 2363
rect 22477 2329 22511 2363
rect 3249 2261 3283 2295
rect 3801 2261 3835 2295
rect 7849 2261 7883 2295
rect 8217 2261 8251 2295
rect 9045 2261 9079 2295
rect 9597 2261 9631 2295
rect 10609 2261 10643 2295
rect 11345 2261 11379 2295
rect 12633 2261 12667 2295
rect 12817 2261 12851 2295
rect 13553 2261 13587 2295
rect 14105 2261 14139 2295
rect 16129 2261 16163 2295
rect 16773 2261 16807 2295
rect 17325 2261 17359 2295
rect 18521 2261 18555 2295
rect 18889 2261 18923 2295
rect 20453 2261 20487 2295
rect 20913 2261 20947 2295
rect 21557 2261 21591 2295
rect 21925 2261 21959 2295
rect 22569 2261 22603 2295
rect 3433 2057 3467 2091
rect 6285 2057 6319 2091
rect 7389 2057 7423 2091
rect 8769 2057 8803 2091
rect 10425 2057 10459 2091
rect 11897 2057 11931 2091
rect 19717 2057 19751 2091
rect 20085 2057 20119 2091
rect 20913 2057 20947 2091
rect 22385 2057 22419 2091
rect 22477 2057 22511 2091
rect 3893 1989 3927 2023
rect 10149 1989 10183 2023
rect 17877 1989 17911 2023
rect 20361 1989 20395 2023
rect 22845 1989 22879 2023
rect 2421 1921 2455 1955
rect 5549 1921 5583 1955
rect 6101 1921 6135 1955
rect 8585 1921 8619 1955
rect 8953 1921 8987 1955
rect 15853 1921 15887 1955
rect 18061 1921 18095 1955
rect 19901 1921 19935 1955
rect 20269 1921 20303 1955
rect 22293 1921 22327 1955
rect 1041 1853 1075 1887
rect 2329 1853 2363 1887
rect 3065 1853 3099 1887
rect 3801 1853 3835 1887
rect 4077 1853 4111 1887
rect 4537 1853 4571 1887
rect 5273 1853 5307 1887
rect 5733 1853 5767 1887
rect 6561 1853 6595 1887
rect 7297 1853 7331 1887
rect 7481 1853 7515 1887
rect 8217 1853 8251 1887
rect 8861 1853 8895 1887
rect 9137 1853 9171 1887
rect 9229 1853 9263 1887
rect 9321 1853 9355 1887
rect 9873 1853 9907 1887
rect 9965 1853 9999 1887
rect 10241 1853 10275 1887
rect 10701 1853 10735 1887
rect 10904 1853 10938 1887
rect 11253 1853 11287 1887
rect 11345 1853 11379 1887
rect 11529 1853 11563 1887
rect 11621 1853 11655 1887
rect 11713 1853 11747 1887
rect 12081 1853 12115 1887
rect 12633 1853 12667 1887
rect 12909 1853 12943 1887
rect 14013 1853 14047 1887
rect 15577 1853 15611 1887
rect 15669 1853 15703 1887
rect 17785 1853 17819 1887
rect 18705 1853 18739 1887
rect 19533 1853 19567 1887
rect 19625 1853 19659 1887
rect 19993 1853 20027 1887
rect 20545 1853 20579 1887
rect 21097 1853 21131 1887
rect 21373 1853 21407 1887
rect 21557 1853 21591 1887
rect 21741 1853 21775 1887
rect 22201 1853 22235 1887
rect 22569 1853 22603 1887
rect 22661 1853 22695 1887
rect 3617 1785 3651 1819
rect 8953 1785 8987 1819
rect 10987 1785 11021 1819
rect 15853 1785 15887 1819
rect 18061 1785 18095 1819
rect 21649 1785 21683 1819
rect 857 1717 891 1751
rect 2697 1717 2731 1751
rect 2973 1717 3007 1751
rect 4445 1717 4479 1751
rect 5181 1717 5215 1751
rect 5917 1717 5951 1751
rect 8033 1717 8067 1751
rect 8585 1717 8619 1751
rect 9505 1717 9539 1751
rect 9689 1717 9723 1751
rect 10793 1717 10827 1751
rect 11069 1717 11103 1751
rect 11437 1717 11471 1751
rect 12541 1717 12575 1751
rect 13093 1717 13127 1751
rect 13921 1717 13955 1751
rect 18889 1717 18923 1751
rect 19349 1717 19383 1751
rect 19901 1717 19935 1751
rect 20269 1717 20303 1751
rect 22017 1717 22051 1751
rect 1041 1513 1075 1547
rect 1317 1513 1351 1547
rect 2513 1513 2547 1547
rect 7205 1513 7239 1547
rect 8309 1513 8343 1547
rect 9229 1513 9263 1547
rect 13093 1513 13127 1547
rect 15294 1513 15328 1547
rect 15675 1513 15709 1547
rect 19165 1513 19199 1547
rect 5457 1445 5491 1479
rect 12275 1445 12309 1479
rect 13277 1445 13311 1479
rect 13369 1445 13403 1479
rect 14657 1445 14691 1479
rect 15025 1445 15059 1479
rect 15393 1445 15427 1479
rect 15577 1445 15611 1479
rect 20913 1445 20947 1479
rect 22569 1445 22603 1479
rect 857 1377 891 1411
rect 1501 1377 1535 1411
rect 1869 1377 1903 1411
rect 2053 1377 2087 1411
rect 2145 1377 2179 1411
rect 2329 1377 2363 1411
rect 2789 1377 2823 1411
rect 3341 1377 3375 1411
rect 3985 1377 4019 1411
rect 4629 1377 4663 1411
rect 5273 1377 5307 1411
rect 6009 1377 6043 1411
rect 6745 1377 6779 1411
rect 7389 1377 7423 1411
rect 7573 1377 7607 1411
rect 7941 1377 7975 1411
rect 8125 1377 8159 1411
rect 8493 1377 8527 1411
rect 8677 1377 8711 1411
rect 8953 1377 8987 1411
rect 9045 1377 9079 1411
rect 9413 1377 9447 1411
rect 9597 1377 9631 1411
rect 9873 1377 9907 1411
rect 10425 1377 10459 1411
rect 11345 1377 11379 1411
rect 11529 1377 11563 1411
rect 11713 1377 11747 1411
rect 11989 1377 12023 1411
rect 12081 1377 12115 1411
rect 12192 1377 12226 1411
rect 12541 1377 12575 1411
rect 12725 1377 12759 1411
rect 12909 1377 12943 1411
rect 13001 1377 13035 1411
rect 13645 1377 13679 1411
rect 13921 1377 13955 1411
rect 14289 1377 14323 1411
rect 14473 1377 14507 1411
rect 14749 1377 14783 1411
rect 14841 1377 14875 1411
rect 15117 1377 15151 1411
rect 15209 1377 15243 1411
rect 15761 1377 15795 1411
rect 15853 1377 15887 1411
rect 16221 1377 16255 1411
rect 16589 1377 16623 1411
rect 17049 1377 17083 1411
rect 17141 1377 17175 1411
rect 17877 1377 17911 1411
rect 18613 1377 18647 1411
rect 18797 1377 18831 1411
rect 18981 1377 19015 1411
rect 19073 1377 19107 1411
rect 19717 1377 19751 1411
rect 19993 1377 20027 1411
rect 20361 1377 20395 1411
rect 21281 1377 21315 1411
rect 21557 1377 21591 1411
rect 22201 1377 22235 1411
rect 22845 1377 22879 1411
rect 3433 1309 3467 1343
rect 3709 1309 3743 1343
rect 3893 1309 3927 1343
rect 4537 1309 4571 1343
rect 5917 1309 5951 1343
rect 6837 1309 6871 1343
rect 7113 1309 7147 1343
rect 7665 1309 7699 1343
rect 8217 1309 8251 1343
rect 8769 1309 8803 1343
rect 9229 1309 9263 1343
rect 9321 1309 9355 1343
rect 10149 1309 10183 1343
rect 13369 1309 13403 1343
rect 16773 1309 16807 1343
rect 17325 1309 17359 1343
rect 17601 1309 17635 1343
rect 19441 1309 19475 1343
rect 20269 1309 20303 1343
rect 20637 1309 20671 1343
rect 22293 1309 22327 1343
rect 22477 1309 22511 1343
rect 22569 1309 22603 1343
rect 4353 1241 4387 1275
rect 4997 1241 5031 1275
rect 6377 1241 6411 1275
rect 7757 1241 7791 1275
rect 9781 1241 9815 1275
rect 10241 1241 10275 1275
rect 11345 1241 11379 1275
rect 12541 1241 12575 1275
rect 13553 1241 13587 1275
rect 14289 1241 14323 1275
rect 17233 1241 17267 1275
rect 18613 1241 18647 1275
rect 19901 1241 19935 1275
rect 22385 1241 22419 1275
rect 22753 1241 22787 1275
rect 1685 1173 1719 1207
rect 2973 1173 3007 1207
rect 5641 1173 5675 1207
rect 9965 1173 9999 1207
rect 10609 1173 10643 1207
rect 13277 1173 13311 1207
rect 13829 1173 13863 1207
rect 15025 1173 15059 1207
rect 16313 1173 16347 1207
rect 17693 1173 17727 1207
rect 17785 1173 17819 1207
rect 19533 1173 19567 1207
rect 20085 1173 20119 1207
rect 20177 1173 20211 1207
rect 20453 1173 20487 1207
rect 20545 1173 20579 1207
rect 20821 1173 20855 1207
rect 2513 969 2547 1003
rect 5917 969 5951 1003
rect 6469 969 6503 1003
rect 6837 969 6871 1003
rect 7941 969 7975 1003
rect 8401 969 8435 1003
rect 9229 969 9263 1003
rect 11345 969 11379 1003
rect 14473 969 14507 1003
rect 16681 969 16715 1003
rect 21833 969 21867 1003
rect 22937 969 22971 1003
rect 2145 901 2179 935
rect 3617 901 3651 935
rect 4721 901 4755 935
rect 7389 901 7423 935
rect 8861 901 8895 935
rect 10333 901 10367 935
rect 11713 901 11747 935
rect 15485 901 15519 935
rect 19625 901 19659 935
rect 19901 901 19935 935
rect 20913 901 20947 935
rect 22201 901 22235 935
rect 7021 833 7055 867
rect 7757 833 7791 867
rect 11529 833 11563 867
rect 14289 833 14323 867
rect 20269 833 20303 867
rect 1225 765 1259 799
rect 1593 765 1627 799
rect 1961 765 1995 799
rect 2329 765 2363 799
rect 2697 765 2731 799
rect 3065 765 3099 799
rect 3341 765 3375 799
rect 3433 765 3467 799
rect 3801 765 3835 799
rect 4169 765 4203 799
rect 4537 765 4571 799
rect 4905 765 4939 799
rect 5273 765 5307 799
rect 5641 765 5675 799
rect 5917 765 5951 799
rect 6193 765 6227 799
rect 6377 765 6411 799
rect 7113 765 7147 799
rect 7205 765 7239 799
rect 7481 765 7515 799
rect 8033 765 8067 799
rect 8585 765 8619 799
rect 8677 765 8711 799
rect 9045 765 9079 799
rect 9413 765 9447 799
rect 9781 765 9815 799
rect 10149 765 10183 799
rect 10793 765 10827 799
rect 11069 765 11103 799
rect 11805 765 11839 799
rect 11897 765 11931 799
rect 12541 765 12575 799
rect 12633 765 12667 799
rect 13277 765 13311 799
rect 13829 765 13863 799
rect 14197 765 14231 799
rect 14565 765 14599 799
rect 14657 765 14691 799
rect 15301 765 15335 799
rect 15669 765 15703 799
rect 15853 765 15887 799
rect 15945 765 15979 799
rect 16497 765 16531 799
rect 16681 765 16715 799
rect 17785 765 17819 799
rect 17877 765 17911 799
rect 18153 765 18187 799
rect 18705 765 18739 799
rect 19073 765 19107 799
rect 19441 765 19475 799
rect 19809 765 19843 799
rect 20085 765 20119 799
rect 20361 765 20395 799
rect 20729 765 20763 799
rect 21281 765 21315 799
rect 21649 765 21683 799
rect 22017 765 22051 799
rect 22385 765 22419 799
rect 22753 765 22787 799
rect 6101 697 6135 731
rect 11345 697 11379 731
rect 11529 697 11563 731
rect 14289 697 14323 731
rect 1041 629 1075 663
rect 1409 629 1443 663
rect 1777 629 1811 663
rect 2881 629 2915 663
rect 3985 629 4019 663
rect 4353 629 4387 663
rect 5089 629 5123 663
rect 5457 629 5491 663
rect 7665 629 7699 663
rect 7757 629 7791 663
rect 9597 629 9631 663
rect 9965 629 9999 663
rect 10609 629 10643 663
rect 11161 629 11195 663
rect 12081 629 12115 663
rect 12357 629 12391 663
rect 12817 629 12851 663
rect 13093 629 13127 663
rect 13645 629 13679 663
rect 14013 629 14047 663
rect 14841 629 14875 663
rect 15117 629 15151 663
rect 17693 629 17727 663
rect 18061 629 18095 663
rect 18337 629 18371 663
rect 18889 629 18923 663
rect 19257 629 19291 663
rect 20545 629 20579 663
rect 21465 629 21499 663
rect 22569 629 22603 663
<< metal1 >>
rect 17954 23712 17960 23724
rect 9646 23684 17960 23712
rect 2222 23604 2228 23656
rect 2280 23644 2286 23656
rect 9646 23644 9674 23684
rect 17954 23672 17960 23684
rect 18012 23672 18018 23724
rect 17218 23644 17224 23656
rect 2280 23616 9674 23644
rect 12406 23616 17224 23644
rect 2280 23604 2286 23616
rect 4154 23536 4160 23588
rect 4212 23576 4218 23588
rect 12406 23576 12434 23616
rect 17218 23604 17224 23616
rect 17276 23604 17282 23656
rect 4212 23548 12434 23576
rect 4212 23536 4218 23548
rect 6086 23468 6092 23520
rect 6144 23508 6150 23520
rect 20070 23508 20076 23520
rect 6144 23480 20076 23508
rect 6144 23468 6150 23480
rect 20070 23468 20076 23480
rect 20128 23468 20134 23520
rect 552 23418 23368 23440
rect 552 23366 4366 23418
rect 4418 23366 4430 23418
rect 4482 23366 4494 23418
rect 4546 23366 4558 23418
rect 4610 23366 4622 23418
rect 4674 23366 4686 23418
rect 4738 23366 10366 23418
rect 10418 23366 10430 23418
rect 10482 23366 10494 23418
rect 10546 23366 10558 23418
rect 10610 23366 10622 23418
rect 10674 23366 10686 23418
rect 10738 23366 16366 23418
rect 16418 23366 16430 23418
rect 16482 23366 16494 23418
rect 16546 23366 16558 23418
rect 16610 23366 16622 23418
rect 16674 23366 16686 23418
rect 16738 23366 22366 23418
rect 22418 23366 22430 23418
rect 22482 23366 22494 23418
rect 22546 23366 22558 23418
rect 22610 23366 22622 23418
rect 22674 23366 22686 23418
rect 22738 23366 23368 23418
rect 552 23344 23368 23366
rect 3050 23264 3056 23316
rect 3108 23304 3114 23316
rect 8113 23307 8171 23313
rect 3108 23276 6500 23304
rect 3108 23264 3114 23276
rect 6472 23236 6500 23276
rect 8113 23273 8125 23307
rect 8159 23304 8171 23307
rect 8294 23304 8300 23316
rect 8159 23276 8300 23304
rect 8159 23273 8171 23276
rect 8113 23267 8171 23273
rect 8294 23264 8300 23276
rect 8352 23264 8358 23316
rect 10226 23264 10232 23316
rect 10284 23304 10290 23316
rect 10321 23307 10379 23313
rect 10321 23304 10333 23307
rect 10284 23276 10333 23304
rect 10284 23264 10290 23276
rect 10321 23273 10333 23276
rect 10367 23273 10379 23307
rect 10321 23267 10379 23273
rect 10597 23307 10655 23313
rect 10597 23273 10609 23307
rect 10643 23304 10655 23307
rect 11054 23304 11060 23316
rect 10643 23276 11060 23304
rect 10643 23273 10655 23276
rect 10597 23267 10655 23273
rect 11054 23264 11060 23276
rect 11112 23264 11118 23316
rect 11425 23307 11483 23313
rect 11425 23273 11437 23307
rect 11471 23304 11483 23307
rect 11606 23304 11612 23316
rect 11471 23276 11612 23304
rect 11471 23273 11483 23276
rect 11425 23267 11483 23273
rect 11606 23264 11612 23276
rect 11664 23264 11670 23316
rect 11790 23264 11796 23316
rect 11848 23264 11854 23316
rect 13357 23307 13415 23313
rect 13357 23273 13369 23307
rect 13403 23273 13415 23307
rect 13357 23267 13415 23273
rect 9398 23236 9404 23248
rect 3252 23208 6408 23236
rect 6472 23208 9404 23236
rect 3252 23180 3280 23208
rect 2222 23128 2228 23180
rect 2280 23128 2286 23180
rect 2406 23128 2412 23180
rect 2464 23128 2470 23180
rect 3234 23128 3240 23180
rect 3292 23128 3298 23180
rect 3326 23128 3332 23180
rect 3384 23168 3390 23180
rect 3493 23171 3551 23177
rect 3493 23168 3505 23171
rect 3384 23140 3505 23168
rect 3384 23128 3390 23140
rect 3493 23137 3505 23140
rect 3539 23137 3551 23171
rect 3493 23131 3551 23137
rect 4709 23171 4767 23177
rect 4709 23137 4721 23171
rect 4755 23168 4767 23171
rect 5442 23168 5448 23180
rect 4755 23140 5448 23168
rect 4755 23137 4767 23140
rect 4709 23131 4767 23137
rect 5442 23128 5448 23140
rect 5500 23128 5506 23180
rect 5718 23128 5724 23180
rect 5776 23168 5782 23180
rect 5813 23171 5871 23177
rect 5813 23168 5825 23171
rect 5776 23140 5825 23168
rect 5776 23128 5782 23140
rect 5813 23137 5825 23140
rect 5859 23137 5871 23171
rect 5813 23131 5871 23137
rect 5997 23171 6055 23177
rect 5997 23137 6009 23171
rect 6043 23137 6055 23171
rect 5997 23131 6055 23137
rect 4985 23103 5043 23109
rect 4985 23069 4997 23103
rect 5031 23100 5043 23103
rect 5534 23100 5540 23112
rect 5031 23072 5540 23100
rect 5031 23069 5043 23072
rect 4985 23063 5043 23069
rect 5534 23060 5540 23072
rect 5592 23100 5598 23112
rect 6012 23100 6040 23131
rect 6380 23112 6408 23208
rect 9398 23196 9404 23208
rect 9456 23196 9462 23248
rect 13372 23236 13400 23267
rect 15838 23264 15844 23316
rect 15896 23304 15902 23316
rect 15896 23276 19012 23304
rect 15896 23264 15902 23276
rect 16393 23239 16451 23245
rect 13372 23208 13768 23236
rect 6730 23177 6736 23180
rect 6724 23131 6736 23177
rect 6730 23128 6736 23131
rect 6788 23128 6794 23180
rect 7929 23171 7987 23177
rect 7929 23137 7941 23171
rect 7975 23168 7987 23171
rect 8202 23168 8208 23180
rect 7975 23140 8208 23168
rect 7975 23137 7987 23140
rect 7929 23131 7987 23137
rect 8202 23128 8208 23140
rect 8260 23128 8266 23180
rect 9214 23128 9220 23180
rect 9272 23168 9278 23180
rect 9686 23171 9744 23177
rect 9686 23168 9698 23171
rect 9272 23140 9698 23168
rect 9272 23128 9278 23140
rect 9686 23137 9698 23140
rect 9732 23137 9744 23171
rect 9686 23131 9744 23137
rect 10042 23128 10048 23180
rect 10100 23168 10106 23180
rect 10137 23171 10195 23177
rect 10137 23168 10149 23171
rect 10100 23140 10149 23168
rect 10100 23128 10106 23140
rect 10137 23137 10149 23140
rect 10183 23137 10195 23171
rect 10137 23131 10195 23137
rect 10778 23128 10784 23180
rect 10836 23128 10842 23180
rect 10962 23128 10968 23180
rect 11020 23128 11026 23180
rect 11238 23128 11244 23180
rect 11296 23128 11302 23180
rect 11330 23128 11336 23180
rect 11388 23168 11394 23180
rect 11609 23171 11667 23177
rect 11609 23168 11621 23171
rect 11388 23140 11621 23168
rect 11388 23128 11394 23140
rect 11609 23137 11621 23140
rect 11655 23137 11667 23171
rect 11609 23131 11667 23137
rect 11790 23128 11796 23180
rect 11848 23168 11854 23180
rect 13740 23177 13768 23208
rect 16393 23205 16405 23239
rect 16439 23236 16451 23239
rect 18230 23236 18236 23248
rect 16439 23208 18236 23236
rect 16439 23205 16451 23208
rect 16393 23199 16451 23205
rect 18230 23196 18236 23208
rect 18288 23196 18294 23248
rect 18325 23239 18383 23245
rect 18325 23205 18337 23239
rect 18371 23236 18383 23239
rect 18782 23236 18788 23248
rect 18371 23208 18788 23236
rect 18371 23205 18383 23208
rect 18325 23199 18383 23205
rect 18782 23196 18788 23208
rect 18840 23196 18846 23248
rect 18984 23245 19012 23276
rect 20070 23264 20076 23316
rect 20128 23264 20134 23316
rect 18960 23239 19018 23245
rect 18960 23205 18972 23239
rect 19006 23205 19018 23239
rect 18960 23199 19018 23205
rect 21542 23196 21548 23248
rect 21600 23236 21606 23248
rect 22925 23239 22983 23245
rect 22925 23236 22937 23239
rect 21600 23208 22937 23236
rect 21600 23196 21606 23208
rect 22925 23205 22937 23208
rect 22971 23205 22983 23239
rect 22925 23199 22983 23205
rect 11977 23171 12035 23177
rect 11977 23168 11989 23171
rect 11848 23140 11989 23168
rect 11848 23128 11854 23140
rect 11977 23137 11989 23140
rect 12023 23137 12035 23171
rect 12233 23171 12291 23177
rect 12233 23168 12245 23171
rect 11977 23131 12035 23137
rect 12084 23140 12245 23168
rect 5592 23072 6040 23100
rect 5592 23060 5598 23072
rect 6362 23060 6368 23112
rect 6420 23100 6426 23112
rect 6457 23103 6515 23109
rect 6457 23100 6469 23103
rect 6420 23072 6469 23100
rect 6420 23060 6426 23072
rect 6457 23069 6469 23072
rect 6503 23069 6515 23103
rect 6457 23063 6515 23069
rect 9953 23103 10011 23109
rect 9953 23069 9965 23103
rect 9999 23100 10011 23103
rect 12084 23100 12112 23140
rect 12233 23137 12245 23140
rect 12279 23137 12291 23171
rect 12233 23131 12291 23137
rect 13725 23171 13783 23177
rect 13725 23137 13737 23171
rect 13771 23168 13783 23171
rect 14826 23168 14832 23180
rect 13771 23140 14832 23168
rect 13771 23137 13783 23140
rect 13725 23131 13783 23137
rect 14826 23128 14832 23140
rect 14884 23128 14890 23180
rect 15654 23128 15660 23180
rect 15712 23177 15718 23180
rect 15712 23131 15724 23177
rect 15712 23128 15718 23131
rect 16206 23128 16212 23180
rect 16264 23168 16270 23180
rect 16833 23171 16891 23177
rect 16833 23168 16845 23171
rect 16264 23140 16845 23168
rect 16264 23128 16270 23140
rect 16833 23137 16845 23140
rect 16879 23137 16891 23171
rect 16833 23131 16891 23137
rect 20254 23128 20260 23180
rect 20312 23128 20318 23180
rect 22393 23171 22451 23177
rect 22393 23137 22405 23171
rect 22439 23168 22451 23171
rect 23382 23168 23388 23180
rect 22439 23140 23388 23168
rect 22439 23137 22451 23140
rect 22393 23131 22451 23137
rect 23382 23128 23388 23140
rect 23440 23128 23446 23180
rect 9999 23072 10180 23100
rect 9999 23069 10011 23072
rect 9953 23063 10011 23069
rect 10152 23044 10180 23072
rect 11164 23072 12112 23100
rect 4801 23035 4859 23041
rect 4801 23001 4813 23035
rect 4847 23032 4859 23035
rect 5074 23032 5080 23044
rect 4847 23004 5080 23032
rect 4847 23001 4859 23004
rect 4801 22995 4859 23001
rect 5074 22992 5080 23004
rect 5132 22992 5138 23044
rect 10134 22992 10140 23044
rect 10192 22992 10198 23044
rect 11164 23041 11192 23072
rect 13814 23060 13820 23112
rect 13872 23100 13878 23112
rect 13872 23072 14596 23100
rect 13872 23060 13878 23072
rect 14568 23041 14596 23072
rect 15930 23060 15936 23112
rect 15988 23100 15994 23112
rect 16577 23103 16635 23109
rect 16577 23100 16589 23103
rect 15988 23072 16589 23100
rect 15988 23060 15994 23072
rect 16577 23069 16589 23072
rect 16623 23069 16635 23103
rect 16577 23063 16635 23069
rect 18690 23060 18696 23112
rect 18748 23060 18754 23112
rect 20533 23103 20591 23109
rect 20533 23069 20545 23103
rect 20579 23100 20591 23103
rect 20806 23100 20812 23112
rect 20579 23072 20812 23100
rect 20579 23069 20591 23072
rect 20533 23063 20591 23069
rect 20806 23060 20812 23072
rect 20864 23060 20870 23112
rect 22649 23103 22707 23109
rect 22649 23069 22661 23103
rect 22695 23100 22707 23103
rect 22830 23100 22836 23112
rect 22695 23072 22836 23100
rect 22695 23069 22707 23072
rect 22649 23063 22707 23069
rect 22830 23060 22836 23072
rect 22888 23060 22894 23112
rect 11149 23035 11207 23041
rect 11149 23001 11161 23035
rect 11195 23001 11207 23035
rect 11149 22995 11207 23001
rect 14553 23035 14611 23041
rect 14553 23001 14565 23035
rect 14599 23001 14611 23035
rect 14553 22995 14611 23001
rect 16022 22992 16028 23044
rect 16080 23032 16086 23044
rect 16209 23035 16267 23041
rect 16209 23032 16221 23035
rect 16080 23004 16221 23032
rect 16080 22992 16086 23004
rect 16209 23001 16221 23004
rect 16255 23001 16267 23035
rect 16209 22995 16267 23001
rect 17954 22992 17960 23044
rect 18012 22992 18018 23044
rect 1762 22924 1768 22976
rect 1820 22964 1826 22976
rect 2317 22967 2375 22973
rect 2317 22964 2329 22967
rect 1820 22936 2329 22964
rect 1820 22924 1826 22936
rect 2317 22933 2329 22936
rect 2363 22933 2375 22967
rect 2317 22927 2375 22933
rect 3970 22924 3976 22976
rect 4028 22964 4034 22976
rect 4617 22967 4675 22973
rect 4617 22964 4629 22967
rect 4028 22936 4629 22964
rect 4028 22924 4034 22936
rect 4617 22933 4629 22936
rect 4663 22933 4675 22967
rect 4617 22927 4675 22933
rect 4890 22924 4896 22976
rect 4948 22924 4954 22976
rect 5442 22924 5448 22976
rect 5500 22964 5506 22976
rect 5905 22967 5963 22973
rect 5905 22964 5917 22967
rect 5500 22936 5917 22964
rect 5500 22924 5506 22936
rect 5905 22933 5917 22936
rect 5951 22933 5963 22967
rect 5905 22927 5963 22933
rect 7837 22967 7895 22973
rect 7837 22933 7849 22967
rect 7883 22964 7895 22967
rect 8110 22964 8116 22976
rect 7883 22936 8116 22964
rect 7883 22933 7895 22936
rect 7837 22927 7895 22933
rect 8110 22924 8116 22936
rect 8168 22924 8174 22976
rect 8570 22924 8576 22976
rect 8628 22924 8634 22976
rect 13170 22924 13176 22976
rect 13228 22964 13234 22976
rect 13541 22967 13599 22973
rect 13541 22964 13553 22967
rect 13228 22936 13553 22964
rect 13228 22924 13234 22936
rect 13541 22933 13553 22936
rect 13587 22933 13599 22967
rect 13541 22927 13599 22933
rect 14458 22924 14464 22976
rect 14516 22924 14522 22976
rect 18417 22967 18475 22973
rect 18417 22933 18429 22967
rect 18463 22964 18475 22967
rect 18874 22964 18880 22976
rect 18463 22936 18880 22964
rect 18463 22933 18475 22936
rect 18417 22927 18475 22933
rect 18874 22924 18880 22936
rect 18932 22924 18938 22976
rect 21269 22967 21327 22973
rect 21269 22933 21281 22967
rect 21315 22964 21327 22967
rect 21358 22964 21364 22976
rect 21315 22936 21364 22964
rect 21315 22933 21327 22936
rect 21269 22927 21327 22933
rect 21358 22924 21364 22936
rect 21416 22924 21422 22976
rect 21634 22924 21640 22976
rect 21692 22964 21698 22976
rect 22833 22967 22891 22973
rect 22833 22964 22845 22967
rect 21692 22936 22845 22964
rect 21692 22924 21698 22936
rect 22833 22933 22845 22936
rect 22879 22933 22891 22967
rect 22833 22927 22891 22933
rect 552 22874 23368 22896
rect 552 22822 1366 22874
rect 1418 22822 1430 22874
rect 1482 22822 1494 22874
rect 1546 22822 1558 22874
rect 1610 22822 1622 22874
rect 1674 22822 1686 22874
rect 1738 22822 7366 22874
rect 7418 22822 7430 22874
rect 7482 22822 7494 22874
rect 7546 22822 7558 22874
rect 7610 22822 7622 22874
rect 7674 22822 7686 22874
rect 7738 22822 13366 22874
rect 13418 22822 13430 22874
rect 13482 22822 13494 22874
rect 13546 22822 13558 22874
rect 13610 22822 13622 22874
rect 13674 22822 13686 22874
rect 13738 22822 19366 22874
rect 19418 22822 19430 22874
rect 19482 22822 19494 22874
rect 19546 22822 19558 22874
rect 19610 22822 19622 22874
rect 19674 22822 19686 22874
rect 19738 22822 23368 22874
rect 552 22800 23368 22822
rect 5534 22720 5540 22772
rect 5592 22720 5598 22772
rect 5718 22720 5724 22772
rect 5776 22720 5782 22772
rect 6641 22763 6699 22769
rect 6641 22729 6653 22763
rect 6687 22760 6699 22763
rect 6730 22760 6736 22772
rect 6687 22732 6736 22760
rect 6687 22729 6699 22732
rect 6641 22723 6699 22729
rect 6730 22720 6736 22732
rect 6788 22720 6794 22772
rect 9214 22720 9220 22772
rect 9272 22720 9278 22772
rect 9490 22720 9496 22772
rect 9548 22720 9554 22772
rect 9861 22763 9919 22769
rect 9861 22729 9873 22763
rect 9907 22760 9919 22763
rect 9950 22760 9956 22772
rect 9907 22732 9956 22760
rect 9907 22729 9919 22732
rect 9861 22723 9919 22729
rect 9950 22720 9956 22732
rect 10008 22720 10014 22772
rect 11238 22760 11244 22772
rect 10060 22732 11244 22760
rect 4798 22692 4804 22704
rect 2700 22664 4804 22692
rect 2700 22633 2728 22664
rect 4798 22652 4804 22664
rect 4856 22652 4862 22704
rect 5626 22652 5632 22704
rect 5684 22652 5690 22704
rect 8570 22692 8576 22704
rect 6380 22664 8576 22692
rect 1581 22627 1639 22633
rect 1581 22593 1593 22627
rect 1627 22624 1639 22627
rect 1949 22627 2007 22633
rect 1949 22624 1961 22627
rect 1627 22596 1961 22624
rect 1627 22593 1639 22596
rect 1581 22587 1639 22593
rect 1949 22593 1961 22596
rect 1995 22624 2007 22627
rect 2685 22627 2743 22633
rect 1995 22596 2636 22624
rect 1995 22593 2007 22596
rect 1949 22587 2007 22593
rect 1486 22516 1492 22568
rect 1544 22516 1550 22568
rect 1673 22559 1731 22565
rect 1673 22525 1685 22559
rect 1719 22556 1731 22559
rect 1762 22556 1768 22568
rect 1719 22528 1768 22556
rect 1719 22525 1731 22528
rect 1673 22519 1731 22525
rect 1762 22516 1768 22528
rect 1820 22516 1826 22568
rect 2608 22565 2636 22596
rect 2685 22593 2697 22627
rect 2731 22593 2743 22627
rect 2685 22587 2743 22593
rect 2133 22559 2191 22565
rect 2133 22525 2145 22559
rect 2179 22525 2191 22559
rect 2133 22519 2191 22525
rect 2593 22559 2651 22565
rect 2593 22525 2605 22559
rect 2639 22525 2651 22559
rect 2593 22519 2651 22525
rect 1857 22491 1915 22497
rect 1857 22457 1869 22491
rect 1903 22457 1915 22491
rect 2148 22488 2176 22519
rect 2700 22488 2728 22587
rect 2958 22584 2964 22636
rect 3016 22584 3022 22636
rect 3605 22627 3663 22633
rect 3605 22593 3617 22627
rect 3651 22624 3663 22627
rect 4246 22624 4252 22636
rect 3651 22596 4252 22624
rect 3651 22593 3663 22596
rect 3605 22587 3663 22593
rect 4246 22584 4252 22596
rect 4304 22624 4310 22636
rect 4433 22627 4491 22633
rect 4433 22624 4445 22627
rect 4304 22596 4445 22624
rect 4304 22584 4310 22596
rect 4433 22593 4445 22596
rect 4479 22593 4491 22627
rect 5644 22624 5672 22652
rect 6086 22624 6092 22636
rect 4433 22587 4491 22593
rect 5460 22596 6092 22624
rect 3513 22559 3571 22565
rect 3513 22525 3525 22559
rect 3559 22525 3571 22559
rect 3513 22519 3571 22525
rect 2148 22460 2728 22488
rect 3528 22488 3556 22519
rect 3694 22516 3700 22568
rect 3752 22516 3758 22568
rect 3970 22516 3976 22568
rect 4028 22516 4034 22568
rect 4154 22516 4160 22568
rect 4212 22516 4218 22568
rect 4709 22559 4767 22565
rect 4709 22525 4721 22559
rect 4755 22556 4767 22559
rect 4890 22556 4896 22568
rect 4755 22528 4896 22556
rect 4755 22525 4767 22528
rect 4709 22519 4767 22525
rect 4890 22516 4896 22528
rect 4948 22516 4954 22568
rect 5460 22565 5488 22596
rect 6086 22584 6092 22596
rect 6144 22584 6150 22636
rect 6380 22565 6408 22664
rect 8570 22652 8576 22664
rect 8628 22652 8634 22704
rect 8941 22695 8999 22701
rect 8941 22661 8953 22695
rect 8987 22692 8999 22695
rect 10060 22692 10088 22732
rect 11238 22720 11244 22732
rect 11296 22720 11302 22772
rect 12069 22763 12127 22769
rect 12069 22760 12081 22763
rect 11348 22732 12081 22760
rect 8987 22664 10088 22692
rect 8987 22661 8999 22664
rect 8941 22655 8999 22661
rect 7377 22627 7435 22633
rect 7377 22593 7389 22627
rect 7423 22624 7435 22627
rect 7834 22624 7840 22636
rect 7423 22596 7840 22624
rect 7423 22593 7435 22596
rect 7377 22587 7435 22593
rect 7834 22584 7840 22596
rect 7892 22584 7898 22636
rect 8110 22584 8116 22636
rect 8168 22624 8174 22636
rect 8481 22627 8539 22633
rect 8481 22624 8493 22627
rect 8168 22596 8493 22624
rect 8168 22584 8174 22596
rect 8481 22593 8493 22596
rect 8527 22593 8539 22627
rect 8481 22587 8539 22593
rect 5445 22559 5503 22565
rect 5445 22525 5457 22559
rect 5491 22525 5503 22559
rect 5445 22519 5503 22525
rect 5629 22559 5687 22565
rect 5629 22525 5641 22559
rect 5675 22556 5687 22559
rect 5905 22559 5963 22565
rect 5905 22556 5917 22559
rect 5675 22528 5917 22556
rect 5675 22525 5687 22528
rect 5629 22519 5687 22525
rect 5905 22525 5917 22528
rect 5951 22556 5963 22559
rect 6365 22559 6423 22565
rect 6365 22556 6377 22559
rect 5951 22528 6377 22556
rect 5951 22525 5963 22528
rect 5905 22519 5963 22525
rect 6365 22525 6377 22528
rect 6411 22525 6423 22559
rect 6365 22519 6423 22525
rect 6457 22559 6515 22565
rect 6457 22525 6469 22559
rect 6503 22556 6515 22559
rect 6503 22528 6776 22556
rect 6503 22525 6515 22528
rect 6457 22519 6515 22525
rect 3528 22460 3832 22488
rect 1857 22451 1915 22457
rect 1762 22380 1768 22432
rect 1820 22420 1826 22432
rect 1872 22420 1900 22451
rect 3804 22429 3832 22460
rect 5074 22448 5080 22500
rect 5132 22488 5138 22500
rect 5534 22488 5540 22500
rect 5132 22460 5540 22488
rect 5132 22448 5138 22460
rect 5534 22448 5540 22460
rect 5592 22448 5598 22500
rect 6086 22448 6092 22500
rect 6144 22448 6150 22500
rect 1820 22392 1900 22420
rect 3789 22423 3847 22429
rect 1820 22380 1826 22392
rect 3789 22389 3801 22423
rect 3835 22420 3847 22423
rect 5258 22420 5264 22432
rect 3835 22392 5264 22420
rect 3835 22389 3847 22392
rect 3789 22383 3847 22389
rect 5258 22380 5264 22392
rect 5316 22380 5322 22432
rect 5350 22380 5356 22432
rect 5408 22380 5414 22432
rect 6178 22380 6184 22432
rect 6236 22380 6242 22432
rect 6748 22429 6776 22528
rect 7282 22516 7288 22568
rect 7340 22556 7346 22568
rect 8573 22559 8631 22565
rect 8573 22556 8585 22559
rect 7340 22528 8585 22556
rect 7340 22516 7346 22528
rect 8573 22525 8585 22528
rect 8619 22525 8631 22559
rect 8573 22519 8631 22525
rect 9033 22559 9091 22565
rect 9033 22525 9045 22559
rect 9079 22556 9091 22559
rect 9214 22556 9220 22568
rect 9079 22528 9220 22556
rect 9079 22525 9091 22528
rect 9033 22519 9091 22525
rect 9214 22516 9220 22528
rect 9272 22516 9278 22568
rect 9306 22516 9312 22568
rect 9364 22516 9370 22568
rect 9674 22516 9680 22568
rect 9732 22516 9738 22568
rect 10045 22559 10103 22565
rect 10045 22525 10057 22559
rect 10091 22556 10103 22559
rect 10134 22556 10140 22568
rect 10091 22528 10140 22556
rect 10091 22525 10103 22528
rect 10045 22519 10103 22525
rect 10134 22516 10140 22528
rect 10192 22516 10198 22568
rect 11348 22556 11376 22732
rect 12069 22729 12081 22732
rect 12115 22729 12127 22763
rect 17126 22760 17132 22772
rect 12069 22723 12127 22729
rect 15580 22732 17132 22760
rect 13814 22692 13820 22704
rect 11716 22664 13820 22692
rect 10244 22528 11376 22556
rect 7101 22491 7159 22497
rect 7101 22457 7113 22491
rect 7147 22488 7159 22491
rect 7561 22491 7619 22497
rect 7561 22488 7573 22491
rect 7147 22460 7573 22488
rect 7147 22457 7159 22460
rect 7101 22451 7159 22457
rect 7561 22457 7573 22460
rect 7607 22457 7619 22491
rect 7561 22451 7619 22457
rect 7742 22448 7748 22500
rect 7800 22488 7806 22500
rect 10244 22488 10272 22528
rect 11514 22516 11520 22568
rect 11572 22516 11578 22568
rect 11716 22565 11744 22664
rect 12805 22627 12863 22633
rect 12805 22624 12817 22627
rect 12406 22596 12817 22624
rect 11701 22559 11759 22565
rect 11701 22525 11713 22559
rect 11747 22525 11759 22559
rect 11701 22519 11759 22525
rect 11793 22559 11851 22565
rect 11793 22525 11805 22559
rect 11839 22525 11851 22559
rect 11793 22519 11851 22525
rect 11977 22559 12035 22565
rect 11977 22525 11989 22559
rect 12023 22556 12035 22559
rect 12253 22559 12311 22565
rect 12253 22556 12265 22559
rect 12023 22528 12265 22556
rect 12023 22525 12035 22528
rect 11977 22519 12035 22525
rect 12253 22525 12265 22528
rect 12299 22556 12311 22559
rect 12406 22556 12434 22596
rect 12805 22593 12817 22596
rect 12851 22593 12863 22627
rect 12805 22587 12863 22593
rect 12299 22528 12434 22556
rect 12529 22559 12587 22565
rect 12299 22525 12311 22528
rect 12253 22519 12311 22525
rect 12529 22525 12541 22559
rect 12575 22556 12587 22559
rect 12618 22556 12624 22568
rect 12575 22528 12624 22556
rect 12575 22525 12587 22528
rect 12529 22519 12587 22525
rect 7800 22460 10272 22488
rect 10312 22491 10370 22497
rect 7800 22448 7806 22460
rect 10312 22457 10324 22491
rect 10358 22457 10370 22491
rect 10312 22451 10370 22457
rect 11609 22491 11667 22497
rect 11609 22457 11621 22491
rect 11655 22488 11667 22491
rect 11808 22488 11836 22519
rect 12618 22516 12624 22528
rect 12676 22516 12682 22568
rect 13004 22565 13032 22664
rect 13814 22652 13820 22664
rect 13872 22652 13878 22704
rect 14366 22652 14372 22704
rect 14424 22652 14430 22704
rect 15010 22692 15016 22704
rect 14476 22664 15016 22692
rect 14476 22624 14504 22664
rect 15010 22652 15016 22664
rect 15068 22692 15074 22704
rect 15470 22692 15476 22704
rect 15068 22664 15476 22692
rect 15068 22652 15074 22664
rect 15470 22652 15476 22664
rect 15528 22652 15534 22704
rect 13740 22596 14504 22624
rect 14921 22627 14979 22633
rect 12713 22559 12771 22565
rect 12713 22525 12725 22559
rect 12759 22525 12771 22559
rect 12713 22519 12771 22525
rect 12989 22559 13047 22565
rect 12989 22525 13001 22559
rect 13035 22525 13047 22559
rect 12989 22519 13047 22525
rect 13081 22559 13139 22565
rect 13081 22525 13093 22559
rect 13127 22525 13139 22559
rect 13081 22519 13139 22525
rect 12728 22488 12756 22519
rect 11655 22460 12756 22488
rect 11655 22457 11667 22460
rect 11609 22451 11667 22457
rect 6733 22423 6791 22429
rect 6733 22389 6745 22423
rect 6779 22389 6791 22423
rect 6733 22383 6791 22389
rect 7190 22380 7196 22432
rect 7248 22380 7254 22432
rect 10226 22380 10232 22432
rect 10284 22420 10290 22432
rect 10336 22420 10364 22451
rect 10284 22392 10364 22420
rect 10284 22380 10290 22392
rect 11238 22380 11244 22432
rect 11296 22420 11302 22432
rect 11425 22423 11483 22429
rect 11425 22420 11437 22423
rect 11296 22392 11437 22420
rect 11296 22380 11302 22392
rect 11425 22389 11437 22392
rect 11471 22389 11483 22423
rect 11425 22383 11483 22389
rect 11885 22423 11943 22429
rect 11885 22389 11897 22423
rect 11931 22420 11943 22423
rect 11974 22420 11980 22432
rect 11931 22392 11980 22420
rect 11931 22389 11943 22392
rect 11885 22383 11943 22389
rect 11974 22380 11980 22392
rect 12032 22380 12038 22432
rect 12250 22380 12256 22432
rect 12308 22420 12314 22432
rect 13096 22420 13124 22519
rect 13170 22516 13176 22568
rect 13228 22556 13234 22568
rect 13446 22556 13452 22568
rect 13228 22528 13452 22556
rect 13228 22516 13234 22528
rect 13446 22516 13452 22528
rect 13504 22556 13510 22568
rect 13740 22565 13768 22596
rect 14921 22593 14933 22627
rect 14967 22624 14979 22627
rect 15580 22624 15608 22732
rect 17126 22720 17132 22732
rect 17184 22720 17190 22772
rect 19702 22720 19708 22772
rect 19760 22760 19766 22772
rect 20070 22760 20076 22772
rect 19760 22732 20076 22760
rect 19760 22720 19766 22732
rect 20070 22720 20076 22732
rect 20128 22720 20134 22772
rect 18693 22695 18751 22701
rect 18693 22692 18705 22695
rect 14967 22596 15608 22624
rect 16592 22664 18705 22692
rect 14967 22593 14979 22596
rect 14921 22587 14979 22593
rect 13541 22559 13599 22565
rect 13541 22556 13553 22559
rect 13504 22528 13553 22556
rect 13504 22516 13510 22528
rect 13541 22525 13553 22528
rect 13587 22525 13599 22559
rect 13541 22519 13599 22525
rect 13725 22559 13783 22565
rect 13725 22525 13737 22559
rect 13771 22525 13783 22559
rect 13725 22519 13783 22525
rect 14458 22516 14464 22568
rect 14516 22556 14522 22568
rect 15105 22559 15163 22565
rect 15105 22556 15117 22559
rect 14516 22528 15117 22556
rect 14516 22516 14522 22528
rect 15105 22525 15117 22528
rect 15151 22525 15163 22559
rect 15105 22519 15163 22525
rect 15194 22516 15200 22568
rect 15252 22556 15258 22568
rect 15565 22559 15623 22565
rect 15565 22556 15577 22559
rect 15252 22528 15577 22556
rect 15252 22516 15258 22528
rect 15565 22525 15577 22528
rect 15611 22556 15623 22559
rect 15611 22528 15976 22556
rect 15611 22525 15623 22528
rect 15565 22519 15623 22525
rect 15948 22500 15976 22528
rect 16114 22516 16120 22568
rect 16172 22556 16178 22568
rect 16592 22556 16620 22664
rect 18693 22661 18705 22664
rect 18739 22661 18751 22695
rect 18693 22655 18751 22661
rect 19058 22652 19064 22704
rect 19116 22692 19122 22704
rect 19116 22664 19288 22692
rect 19116 22652 19122 22664
rect 17310 22584 17316 22636
rect 17368 22624 17374 22636
rect 17589 22627 17647 22633
rect 17589 22624 17601 22627
rect 17368 22596 17601 22624
rect 17368 22584 17374 22596
rect 17589 22593 17601 22596
rect 17635 22593 17647 22627
rect 17589 22587 17647 22593
rect 17954 22584 17960 22636
rect 18012 22624 18018 22636
rect 19260 22633 19288 22664
rect 19794 22652 19800 22704
rect 19852 22692 19858 22704
rect 19852 22664 20852 22692
rect 19852 22652 19858 22664
rect 19245 22627 19303 22633
rect 18012 22596 19104 22624
rect 18012 22584 18018 22596
rect 19076 22565 19104 22596
rect 19245 22593 19257 22627
rect 19291 22624 19303 22627
rect 20073 22627 20131 22633
rect 20073 22624 20085 22627
rect 19291 22596 20085 22624
rect 19291 22593 19303 22596
rect 19245 22587 19303 22593
rect 20073 22593 20085 22596
rect 20119 22593 20131 22627
rect 20824 22624 20852 22664
rect 20898 22652 20904 22704
rect 20956 22692 20962 22704
rect 21545 22695 21603 22701
rect 21545 22692 21557 22695
rect 20956 22664 21557 22692
rect 20956 22652 20962 22664
rect 21545 22661 21557 22664
rect 21591 22661 21603 22695
rect 21545 22655 21603 22661
rect 20824 22596 21220 22624
rect 20073 22587 20131 22593
rect 18417 22559 18475 22565
rect 18417 22556 18429 22559
rect 16172 22528 16620 22556
rect 17052 22528 18429 22556
rect 16172 22516 16178 22528
rect 13630 22448 13636 22500
rect 13688 22488 13694 22500
rect 13909 22491 13967 22497
rect 13909 22488 13921 22491
rect 13688 22460 13921 22488
rect 13688 22448 13694 22460
rect 13909 22457 13921 22460
rect 13955 22488 13967 22491
rect 14001 22491 14059 22497
rect 14001 22488 14013 22491
rect 13955 22460 14013 22488
rect 13955 22457 13967 22460
rect 13909 22451 13967 22457
rect 14001 22457 14013 22460
rect 14047 22457 14059 22491
rect 14001 22451 14059 22457
rect 14550 22448 14556 22500
rect 14608 22488 14614 22500
rect 15810 22491 15868 22497
rect 15810 22488 15822 22491
rect 14608 22460 15822 22488
rect 14608 22448 14614 22460
rect 15810 22457 15822 22460
rect 15856 22457 15868 22491
rect 15810 22451 15868 22457
rect 15930 22448 15936 22500
rect 15988 22448 15994 22500
rect 17052 22488 17080 22528
rect 18417 22525 18429 22528
rect 18463 22525 18475 22559
rect 18417 22519 18475 22525
rect 19061 22559 19119 22565
rect 19061 22525 19073 22559
rect 19107 22525 19119 22559
rect 19061 22519 19119 22525
rect 19153 22559 19211 22565
rect 19153 22525 19165 22559
rect 19199 22556 19211 22559
rect 20438 22556 20444 22568
rect 19199 22528 20444 22556
rect 19199 22525 19211 22528
rect 19153 22519 19211 22525
rect 20438 22516 20444 22528
rect 20496 22516 20502 22568
rect 20533 22559 20591 22565
rect 20533 22525 20545 22559
rect 20579 22556 20591 22559
rect 20901 22559 20959 22565
rect 20579 22528 20852 22556
rect 20579 22525 20591 22528
rect 20533 22519 20591 22525
rect 16960 22460 17080 22488
rect 17405 22491 17463 22497
rect 12308 22392 13124 22420
rect 12308 22380 12314 22392
rect 14274 22380 14280 22432
rect 14332 22420 14338 22432
rect 14461 22423 14519 22429
rect 14461 22420 14473 22423
rect 14332 22392 14473 22420
rect 14332 22380 14338 22392
rect 14461 22389 14473 22392
rect 14507 22389 14519 22423
rect 14461 22383 14519 22389
rect 15013 22423 15071 22429
rect 15013 22389 15025 22423
rect 15059 22420 15071 22423
rect 15102 22420 15108 22432
rect 15059 22392 15108 22420
rect 15059 22389 15071 22392
rect 15013 22383 15071 22389
rect 15102 22380 15108 22392
rect 15160 22380 15166 22432
rect 15378 22380 15384 22432
rect 15436 22420 15442 22432
rect 15473 22423 15531 22429
rect 15473 22420 15485 22423
rect 15436 22392 15485 22420
rect 15436 22380 15442 22392
rect 15473 22389 15485 22392
rect 15519 22389 15531 22423
rect 15473 22383 15531 22389
rect 15562 22380 15568 22432
rect 15620 22420 15626 22432
rect 16960 22429 16988 22460
rect 17405 22457 17417 22491
rect 17451 22488 17463 22491
rect 17865 22491 17923 22497
rect 17865 22488 17877 22491
rect 17451 22460 17877 22488
rect 17451 22457 17463 22460
rect 17405 22451 17463 22457
rect 17865 22457 17877 22460
rect 17911 22457 17923 22491
rect 20254 22488 20260 22500
rect 17865 22451 17923 22457
rect 19076 22460 20260 22488
rect 16945 22423 17003 22429
rect 16945 22420 16957 22423
rect 15620 22392 16957 22420
rect 15620 22380 15626 22392
rect 16945 22389 16957 22392
rect 16991 22389 17003 22423
rect 16945 22383 17003 22389
rect 17034 22380 17040 22432
rect 17092 22380 17098 22432
rect 17497 22423 17555 22429
rect 17497 22389 17509 22423
rect 17543 22420 17555 22423
rect 19076 22420 19104 22460
rect 20254 22448 20260 22460
rect 20312 22448 20318 22500
rect 20622 22448 20628 22500
rect 20680 22448 20686 22500
rect 20714 22448 20720 22500
rect 20772 22448 20778 22500
rect 20824 22488 20852 22528
rect 20901 22525 20913 22559
rect 20947 22556 20959 22559
rect 21082 22556 21088 22568
rect 20947 22528 21088 22556
rect 20947 22525 20959 22528
rect 20901 22519 20959 22525
rect 21082 22516 21088 22528
rect 21140 22516 21146 22568
rect 21192 22565 21220 22596
rect 21177 22559 21235 22565
rect 21177 22525 21189 22559
rect 21223 22525 21235 22559
rect 21177 22519 21235 22525
rect 22186 22516 22192 22568
rect 22244 22556 22250 22568
rect 22830 22556 22836 22568
rect 22244 22528 22836 22556
rect 22244 22516 22250 22528
rect 22830 22516 22836 22528
rect 22888 22556 22894 22568
rect 22925 22559 22983 22565
rect 22925 22556 22937 22559
rect 22888 22528 22937 22556
rect 22888 22516 22894 22528
rect 22925 22525 22937 22528
rect 22971 22525 22983 22559
rect 22925 22519 22983 22525
rect 21634 22488 21640 22500
rect 20824 22460 21640 22488
rect 21634 22448 21640 22460
rect 21692 22448 21698 22500
rect 22680 22491 22738 22497
rect 22680 22457 22692 22491
rect 22726 22488 22738 22491
rect 23014 22488 23020 22500
rect 22726 22460 23020 22488
rect 22726 22457 22738 22460
rect 22680 22451 22738 22457
rect 23014 22448 23020 22460
rect 23072 22448 23078 22500
rect 17543 22392 19104 22420
rect 17543 22389 17555 22392
rect 17497 22383 17555 22389
rect 19334 22380 19340 22432
rect 19392 22420 19398 22432
rect 19521 22423 19579 22429
rect 19521 22420 19533 22423
rect 19392 22392 19533 22420
rect 19392 22380 19398 22392
rect 19521 22389 19533 22392
rect 19567 22389 19579 22423
rect 19521 22383 19579 22389
rect 19702 22380 19708 22432
rect 19760 22420 19766 22432
rect 19889 22423 19947 22429
rect 19889 22420 19901 22423
rect 19760 22392 19901 22420
rect 19760 22380 19766 22392
rect 19889 22389 19901 22392
rect 19935 22389 19947 22423
rect 19889 22383 19947 22389
rect 19981 22423 20039 22429
rect 19981 22389 19993 22423
rect 20027 22420 20039 22423
rect 20349 22423 20407 22429
rect 20349 22420 20361 22423
rect 20027 22392 20361 22420
rect 20027 22389 20039 22392
rect 19981 22383 20039 22389
rect 20349 22389 20361 22392
rect 20395 22389 20407 22423
rect 20349 22383 20407 22389
rect 21082 22380 21088 22432
rect 21140 22380 21146 22432
rect 552 22330 23368 22352
rect 552 22278 4366 22330
rect 4418 22278 4430 22330
rect 4482 22278 4494 22330
rect 4546 22278 4558 22330
rect 4610 22278 4622 22330
rect 4674 22278 4686 22330
rect 4738 22278 10366 22330
rect 10418 22278 10430 22330
rect 10482 22278 10494 22330
rect 10546 22278 10558 22330
rect 10610 22278 10622 22330
rect 10674 22278 10686 22330
rect 10738 22278 16366 22330
rect 16418 22278 16430 22330
rect 16482 22278 16494 22330
rect 16546 22278 16558 22330
rect 16610 22278 16622 22330
rect 16674 22278 16686 22330
rect 16738 22278 22366 22330
rect 22418 22278 22430 22330
rect 22482 22278 22494 22330
rect 22546 22278 22558 22330
rect 22610 22278 22622 22330
rect 22674 22278 22686 22330
rect 22738 22278 23368 22330
rect 552 22256 23368 22278
rect 1486 22176 1492 22228
rect 1544 22216 1550 22228
rect 1949 22219 2007 22225
rect 1949 22216 1961 22219
rect 1544 22188 1961 22216
rect 1544 22176 1550 22188
rect 1949 22185 1961 22188
rect 1995 22185 2007 22219
rect 1949 22179 2007 22185
rect 2406 22176 2412 22228
rect 2464 22216 2470 22228
rect 2593 22219 2651 22225
rect 2593 22216 2605 22219
rect 2464 22188 2605 22216
rect 2464 22176 2470 22188
rect 2593 22185 2605 22188
rect 2639 22185 2651 22219
rect 2593 22179 2651 22185
rect 2869 22219 2927 22225
rect 2869 22185 2881 22219
rect 2915 22216 2927 22219
rect 3326 22216 3332 22228
rect 2915 22188 3332 22216
rect 2915 22185 2927 22188
rect 2869 22179 2927 22185
rect 2222 22108 2228 22160
rect 2280 22148 2286 22160
rect 2317 22151 2375 22157
rect 2317 22148 2329 22151
rect 2280 22120 2329 22148
rect 2280 22108 2286 22120
rect 2317 22117 2329 22120
rect 2363 22117 2375 22151
rect 2608 22148 2636 22179
rect 3326 22176 3332 22188
rect 3384 22176 3390 22228
rect 4798 22176 4804 22228
rect 4856 22176 4862 22228
rect 5442 22216 5448 22228
rect 4908 22188 5448 22216
rect 3510 22148 3516 22160
rect 2608 22120 3516 22148
rect 2317 22111 2375 22117
rect 3510 22108 3516 22120
rect 3568 22108 3574 22160
rect 3694 22108 3700 22160
rect 3752 22148 3758 22160
rect 4908 22148 4936 22188
rect 5442 22176 5448 22188
rect 5500 22176 5506 22228
rect 5534 22176 5540 22228
rect 5592 22216 5598 22228
rect 5592 22188 6500 22216
rect 5592 22176 5598 22188
rect 3752 22120 4016 22148
rect 3752 22108 3758 22120
rect 1673 22083 1731 22089
rect 1673 22049 1685 22083
rect 1719 22049 1731 22083
rect 1673 22043 1731 22049
rect 1688 22012 1716 22043
rect 1854 22040 1860 22092
rect 1912 22040 1918 22092
rect 2038 22040 2044 22092
rect 2096 22080 2102 22092
rect 2133 22083 2191 22089
rect 2133 22080 2145 22083
rect 2096 22052 2145 22080
rect 2096 22040 2102 22052
rect 2133 22049 2145 22052
rect 2179 22080 2191 22083
rect 2409 22083 2467 22089
rect 2409 22080 2421 22083
rect 2179 22052 2421 22080
rect 2179 22049 2191 22052
rect 2133 22043 2191 22049
rect 2409 22049 2421 22052
rect 2455 22049 2467 22083
rect 2409 22043 2467 22049
rect 2777 22083 2835 22089
rect 2777 22049 2789 22083
rect 2823 22049 2835 22083
rect 2777 22043 2835 22049
rect 2222 22012 2228 22024
rect 1688 21984 2228 22012
rect 2222 21972 2228 21984
rect 2280 21972 2286 22024
rect 2792 21944 2820 22043
rect 2958 22040 2964 22092
rect 3016 22040 3022 22092
rect 3329 22083 3387 22089
rect 3329 22049 3341 22083
rect 3375 22080 3387 22083
rect 3418 22080 3424 22092
rect 3375 22052 3424 22080
rect 3375 22049 3387 22052
rect 3329 22043 3387 22049
rect 3418 22040 3424 22052
rect 3476 22040 3482 22092
rect 3605 22083 3663 22089
rect 3605 22049 3617 22083
rect 3651 22049 3663 22083
rect 3605 22043 3663 22049
rect 3789 22083 3847 22089
rect 3789 22049 3801 22083
rect 3835 22080 3847 22083
rect 3878 22080 3884 22092
rect 3835 22052 3884 22080
rect 3835 22049 3847 22052
rect 3789 22043 3847 22049
rect 2866 21972 2872 22024
rect 2924 22012 2930 22024
rect 3050 22012 3056 22024
rect 2924 21984 3056 22012
rect 2924 21972 2930 21984
rect 3050 21972 3056 21984
rect 3108 21972 3114 22024
rect 3620 22012 3648 22043
rect 3878 22040 3884 22052
rect 3936 22040 3942 22092
rect 3988 22080 4016 22120
rect 4632 22120 4936 22148
rect 5460 22148 5488 22176
rect 6472 22160 6500 22188
rect 7190 22176 7196 22228
rect 7248 22216 7254 22228
rect 7285 22219 7343 22225
rect 7285 22216 7297 22219
rect 7248 22188 7297 22216
rect 7248 22176 7254 22188
rect 7285 22185 7297 22188
rect 7331 22185 7343 22219
rect 7285 22179 7343 22185
rect 8297 22219 8355 22225
rect 8297 22185 8309 22219
rect 8343 22216 8355 22219
rect 8662 22216 8668 22228
rect 8343 22188 8668 22216
rect 8343 22185 8355 22188
rect 8297 22179 8355 22185
rect 5460 22120 6040 22148
rect 4632 22089 4660 22120
rect 4157 22083 4215 22089
rect 4157 22080 4169 22083
rect 3988 22052 4169 22080
rect 4157 22049 4169 22052
rect 4203 22049 4215 22083
rect 4157 22043 4215 22049
rect 4341 22083 4399 22089
rect 4341 22049 4353 22083
rect 4387 22080 4399 22083
rect 4617 22083 4675 22089
rect 4387 22052 4568 22080
rect 4387 22049 4399 22052
rect 4341 22043 4399 22049
rect 4062 22012 4068 22024
rect 3620 21984 4068 22012
rect 4062 21972 4068 21984
rect 4120 21972 4126 22024
rect 4246 21972 4252 22024
rect 4304 22012 4310 22024
rect 4433 22015 4491 22021
rect 4433 22012 4445 22015
rect 4304 21984 4445 22012
rect 4304 21972 4310 21984
rect 4433 21981 4445 21984
rect 4479 21981 4491 22015
rect 4540 22012 4568 22052
rect 4617 22049 4629 22083
rect 4663 22049 4675 22083
rect 4617 22043 4675 22049
rect 4706 22040 4712 22092
rect 4764 22080 4770 22092
rect 5077 22083 5135 22089
rect 5077 22080 5089 22083
rect 4764 22052 5089 22080
rect 4764 22040 4770 22052
rect 5077 22049 5089 22052
rect 5123 22080 5135 22083
rect 5166 22080 5172 22092
rect 5123 22052 5172 22080
rect 5123 22049 5135 22052
rect 5077 22043 5135 22049
rect 5166 22040 5172 22052
rect 5224 22040 5230 22092
rect 5258 22040 5264 22092
rect 5316 22040 5322 22092
rect 5442 22040 5448 22092
rect 5500 22040 5506 22092
rect 6012 22089 6040 22120
rect 6454 22108 6460 22160
rect 6512 22148 6518 22160
rect 7742 22148 7748 22160
rect 6512 22120 7748 22148
rect 6512 22108 6518 22120
rect 7742 22108 7748 22120
rect 7800 22108 7806 22160
rect 8312 22148 8340 22179
rect 8662 22176 8668 22188
rect 8720 22176 8726 22228
rect 9033 22219 9091 22225
rect 9033 22185 9045 22219
rect 9079 22216 9091 22219
rect 9309 22219 9367 22225
rect 9309 22216 9321 22219
rect 9079 22188 9321 22216
rect 9079 22185 9091 22188
rect 9033 22179 9091 22185
rect 9309 22185 9321 22188
rect 9355 22185 9367 22219
rect 9309 22179 9367 22185
rect 9674 22176 9680 22228
rect 9732 22216 9738 22228
rect 10321 22219 10379 22225
rect 9732 22188 10272 22216
rect 9732 22176 9738 22188
rect 7852 22120 8340 22148
rect 5537 22083 5595 22089
rect 5537 22049 5549 22083
rect 5583 22049 5595 22083
rect 5997 22083 6055 22089
rect 5997 22080 6009 22083
rect 5975 22052 6009 22080
rect 5537 22043 5595 22049
rect 5997 22049 6009 22052
rect 6043 22049 6055 22083
rect 5997 22043 6055 22049
rect 7101 22083 7159 22089
rect 7101 22049 7113 22083
rect 7147 22080 7159 22083
rect 7190 22080 7196 22092
rect 7147 22052 7196 22080
rect 7147 22049 7159 22052
rect 7101 22043 7159 22049
rect 4540 21984 5396 22012
rect 4433 21975 4491 21981
rect 3145 21947 3203 21953
rect 3145 21944 3157 21947
rect 2792 21916 3157 21944
rect 3145 21913 3157 21916
rect 3191 21913 3203 21947
rect 3145 21907 3203 21913
rect 4525 21947 4583 21953
rect 4525 21913 4537 21947
rect 4571 21944 4583 21947
rect 5074 21944 5080 21956
rect 4571 21916 5080 21944
rect 4571 21913 4583 21916
rect 4525 21907 4583 21913
rect 5074 21904 5080 21916
rect 5132 21904 5138 21956
rect 5368 21953 5396 21984
rect 5353 21947 5411 21953
rect 5353 21913 5365 21947
rect 5399 21913 5411 21947
rect 5353 21907 5411 21913
rect 1857 21879 1915 21885
rect 1857 21845 1869 21879
rect 1903 21876 1915 21879
rect 1946 21876 1952 21888
rect 1903 21848 1952 21876
rect 1903 21845 1915 21848
rect 1857 21839 1915 21845
rect 1946 21836 1952 21848
rect 2004 21836 2010 21888
rect 3237 21879 3295 21885
rect 3237 21845 3249 21879
rect 3283 21876 3295 21879
rect 3326 21876 3332 21888
rect 3283 21848 3332 21876
rect 3283 21845 3295 21848
rect 3237 21839 3295 21845
rect 3326 21836 3332 21848
rect 3384 21876 3390 21888
rect 3878 21876 3884 21888
rect 3384 21848 3884 21876
rect 3384 21836 3390 21848
rect 3878 21836 3884 21848
rect 3936 21836 3942 21888
rect 4065 21879 4123 21885
rect 4065 21845 4077 21879
rect 4111 21876 4123 21879
rect 4706 21876 4712 21888
rect 4111 21848 4712 21876
rect 4111 21845 4123 21848
rect 4065 21839 4123 21845
rect 4706 21836 4712 21848
rect 4764 21836 4770 21888
rect 4890 21836 4896 21888
rect 4948 21836 4954 21888
rect 5552 21876 5580 22043
rect 7190 22040 7196 22052
rect 7248 22040 7254 22092
rect 7653 22083 7711 22089
rect 7653 22049 7665 22083
rect 7699 22080 7711 22083
rect 7852 22080 7880 22120
rect 8478 22108 8484 22160
rect 8536 22148 8542 22160
rect 9122 22148 9128 22160
rect 8536 22120 9128 22148
rect 8536 22108 8542 22120
rect 9122 22108 9128 22120
rect 9180 22108 9186 22160
rect 9398 22108 9404 22160
rect 9456 22148 9462 22160
rect 9953 22151 10011 22157
rect 9953 22148 9965 22151
rect 9456 22120 9965 22148
rect 9456 22108 9462 22120
rect 9953 22117 9965 22120
rect 9999 22117 10011 22151
rect 9953 22111 10011 22117
rect 10042 22108 10048 22160
rect 10100 22148 10106 22160
rect 10153 22151 10211 22157
rect 10153 22148 10165 22151
rect 10100 22120 10165 22148
rect 10100 22108 10106 22120
rect 10153 22117 10165 22120
rect 10199 22117 10211 22151
rect 10244 22148 10272 22188
rect 10321 22185 10333 22219
rect 10367 22216 10379 22219
rect 10962 22216 10968 22228
rect 10367 22188 10968 22216
rect 10367 22185 10379 22188
rect 10321 22179 10379 22185
rect 10962 22176 10968 22188
rect 11020 22176 11026 22228
rect 11514 22216 11520 22228
rect 11072 22188 11520 22216
rect 10244 22120 10364 22148
rect 10153 22111 10211 22117
rect 10336 22092 10364 22120
rect 7699 22052 7880 22080
rect 7929 22083 7987 22089
rect 7699 22049 7711 22052
rect 7653 22043 7711 22049
rect 7929 22049 7941 22083
rect 7975 22080 7987 22083
rect 8205 22084 8263 22089
rect 8205 22083 8340 22084
rect 8205 22080 8217 22083
rect 7975 22052 8217 22080
rect 7975 22049 7987 22052
rect 7929 22043 7987 22049
rect 8205 22049 8217 22052
rect 8251 22056 8340 22083
rect 8251 22049 8263 22056
rect 8205 22043 8263 22049
rect 6089 22015 6147 22021
rect 6089 21981 6101 22015
rect 6135 22012 6147 22015
rect 6454 22012 6460 22024
rect 6135 21984 6460 22012
rect 6135 21981 6147 21984
rect 6089 21975 6147 21981
rect 6454 21972 6460 21984
rect 6512 21972 6518 22024
rect 6825 22015 6883 22021
rect 6825 21981 6837 22015
rect 6871 22012 6883 22015
rect 8110 22012 8116 22024
rect 6871 21984 8116 22012
rect 6871 21981 6883 21984
rect 6825 21975 6883 21981
rect 5810 21904 5816 21956
rect 5868 21944 5874 21956
rect 6840 21944 6868 21975
rect 8110 21972 8116 21984
rect 8168 21972 8174 22024
rect 8312 22012 8340 22056
rect 8386 22040 8392 22092
rect 8444 22040 8450 22092
rect 8496 22052 9904 22080
rect 8496 22012 8524 22052
rect 8312 21984 8524 22012
rect 5868 21916 6868 21944
rect 6917 21947 6975 21953
rect 5868 21904 5874 21916
rect 6917 21913 6929 21947
rect 6963 21944 6975 21947
rect 7377 21947 7435 21953
rect 7377 21944 7389 21947
rect 6963 21916 7389 21944
rect 6963 21913 6975 21916
rect 6917 21907 6975 21913
rect 7377 21913 7389 21916
rect 7423 21944 7435 21947
rect 7926 21944 7932 21956
rect 7423 21916 7932 21944
rect 7423 21913 7435 21916
rect 7377 21907 7435 21913
rect 7926 21904 7932 21916
rect 7984 21904 7990 21956
rect 8018 21904 8024 21956
rect 8076 21904 8082 21956
rect 8404 21888 8432 21984
rect 9490 21972 9496 22024
rect 9548 21972 9554 22024
rect 9582 21972 9588 22024
rect 9640 21972 9646 22024
rect 9674 21972 9680 22024
rect 9732 21972 9738 22024
rect 9769 22015 9827 22021
rect 9769 21981 9781 22015
rect 9815 21981 9827 22015
rect 9876 22012 9904 22052
rect 10318 22040 10324 22092
rect 10376 22080 10382 22092
rect 10597 22083 10655 22089
rect 10597 22080 10609 22083
rect 10376 22052 10609 22080
rect 10376 22040 10382 22052
rect 10597 22049 10609 22052
rect 10643 22049 10655 22083
rect 10597 22043 10655 22049
rect 10778 22040 10784 22092
rect 10836 22040 10842 22092
rect 11072 22012 11100 22188
rect 11514 22176 11520 22188
rect 11572 22216 11578 22228
rect 11701 22219 11759 22225
rect 11701 22216 11713 22219
rect 11572 22188 11713 22216
rect 11572 22176 11578 22188
rect 11701 22185 11713 22188
rect 11747 22185 11759 22219
rect 11701 22179 11759 22185
rect 15565 22219 15623 22225
rect 15565 22185 15577 22219
rect 15611 22216 15623 22219
rect 15654 22216 15660 22228
rect 15611 22188 15660 22216
rect 15611 22185 15623 22188
rect 15565 22179 15623 22185
rect 15654 22176 15660 22188
rect 15712 22176 15718 22228
rect 15838 22176 15844 22228
rect 15896 22216 15902 22228
rect 16022 22216 16028 22228
rect 15896 22188 16028 22216
rect 15896 22176 15902 22188
rect 16022 22176 16028 22188
rect 16080 22176 16086 22228
rect 16206 22176 16212 22228
rect 16264 22216 16270 22228
rect 16301 22219 16359 22225
rect 16301 22216 16313 22219
rect 16264 22188 16313 22216
rect 16264 22176 16270 22188
rect 16301 22185 16313 22188
rect 16347 22185 16359 22219
rect 16301 22179 16359 22185
rect 17218 22176 17224 22228
rect 17276 22216 17282 22228
rect 17313 22219 17371 22225
rect 17313 22216 17325 22219
rect 17276 22188 17325 22216
rect 17276 22176 17282 22188
rect 17313 22185 17325 22188
rect 17359 22216 17371 22219
rect 19153 22219 19211 22225
rect 19153 22216 19165 22219
rect 17359 22188 19165 22216
rect 17359 22185 17371 22188
rect 17313 22179 17371 22185
rect 19153 22185 19165 22188
rect 19199 22185 19211 22219
rect 20162 22216 20168 22228
rect 19153 22179 19211 22185
rect 19306 22188 20168 22216
rect 11238 22108 11244 22160
rect 11296 22148 11302 22160
rect 12250 22148 12256 22160
rect 11296 22120 12256 22148
rect 11296 22108 11302 22120
rect 11422 22040 11428 22092
rect 11480 22040 11486 22092
rect 11992 22089 12020 22120
rect 12250 22108 12256 22120
rect 12308 22108 12314 22160
rect 13446 22148 13452 22160
rect 12360 22120 13452 22148
rect 11885 22083 11943 22089
rect 11885 22049 11897 22083
rect 11931 22080 11943 22083
rect 11977 22083 12035 22089
rect 11977 22080 11989 22083
rect 11931 22052 11989 22080
rect 11931 22049 11943 22052
rect 11885 22043 11943 22049
rect 11977 22049 11989 22052
rect 12023 22080 12035 22083
rect 12161 22083 12219 22089
rect 12023 22052 12057 22080
rect 12023 22049 12035 22052
rect 11977 22043 12035 22049
rect 12161 22049 12173 22083
rect 12207 22080 12219 22083
rect 12360 22080 12388 22120
rect 13446 22108 13452 22120
rect 13504 22108 13510 22160
rect 13630 22108 13636 22160
rect 13688 22108 13694 22160
rect 14366 22148 14372 22160
rect 13924 22120 14372 22148
rect 12207 22052 12388 22080
rect 12207 22049 12219 22052
rect 12161 22043 12219 22049
rect 9876 21984 11100 22012
rect 11440 22012 11468 22040
rect 12176 22012 12204 22043
rect 12526 22040 12532 22092
rect 12584 22080 12590 22092
rect 12897 22083 12955 22089
rect 12897 22080 12909 22083
rect 12584 22052 12909 22080
rect 12584 22040 12590 22052
rect 12897 22049 12909 22052
rect 12943 22049 12955 22083
rect 12897 22043 12955 22049
rect 13541 22083 13599 22089
rect 13541 22049 13553 22083
rect 13587 22080 13599 22083
rect 13722 22080 13728 22092
rect 13587 22052 13728 22080
rect 13587 22049 13599 22052
rect 13541 22043 13599 22049
rect 13722 22040 13728 22052
rect 13780 22040 13786 22092
rect 13924 22089 13952 22120
rect 14366 22108 14372 22120
rect 14424 22148 14430 22160
rect 14645 22151 14703 22157
rect 14645 22148 14657 22151
rect 14424 22120 14657 22148
rect 14424 22108 14430 22120
rect 14645 22117 14657 22120
rect 14691 22117 14703 22151
rect 14645 22111 14703 22117
rect 14826 22108 14832 22160
rect 14884 22108 14890 22160
rect 15010 22108 15016 22160
rect 15068 22108 15074 22160
rect 17954 22108 17960 22160
rect 18012 22148 18018 22160
rect 19306 22148 19334 22188
rect 20162 22176 20168 22188
rect 20220 22176 20226 22228
rect 20254 22176 20260 22228
rect 20312 22176 20318 22228
rect 20622 22216 20628 22228
rect 20548 22188 20628 22216
rect 18012 22120 19334 22148
rect 18012 22108 18018 22120
rect 19426 22108 19432 22160
rect 19484 22148 19490 22160
rect 20548 22157 20576 22188
rect 20622 22176 20628 22188
rect 20680 22176 20686 22228
rect 20533 22151 20591 22157
rect 20533 22148 20545 22151
rect 19484 22120 20545 22148
rect 19484 22108 19490 22120
rect 20533 22117 20545 22120
rect 20579 22117 20591 22151
rect 20533 22111 20591 22117
rect 20714 22108 20720 22160
rect 20772 22148 20778 22160
rect 20772 22120 21680 22148
rect 20772 22108 20778 22120
rect 13817 22083 13875 22089
rect 13817 22049 13829 22083
rect 13863 22049 13875 22083
rect 13817 22043 13875 22049
rect 13909 22083 13967 22089
rect 13909 22049 13921 22083
rect 13955 22049 13967 22083
rect 13909 22043 13967 22049
rect 11440 21984 12204 22012
rect 13832 22012 13860 22043
rect 14182 22040 14188 22092
rect 14240 22040 14246 22092
rect 15105 22083 15163 22089
rect 15105 22049 15117 22083
rect 15151 22080 15163 22083
rect 15286 22080 15292 22092
rect 15151 22052 15292 22080
rect 15151 22049 15163 22052
rect 15105 22043 15163 22049
rect 15286 22040 15292 22052
rect 15344 22040 15350 22092
rect 15378 22040 15384 22092
rect 15436 22040 15442 22092
rect 15654 22040 15660 22092
rect 15712 22040 15718 22092
rect 16114 22040 16120 22092
rect 16172 22040 16178 22092
rect 16850 22040 16856 22092
rect 16908 22040 16914 22092
rect 17862 22080 17868 22092
rect 16960 22052 17868 22080
rect 14200 22012 14228 22040
rect 13832 21984 14228 22012
rect 9769 21975 9827 21981
rect 8570 21904 8576 21956
rect 8628 21944 8634 21956
rect 8665 21947 8723 21953
rect 8665 21944 8677 21947
rect 8628 21916 8677 21944
rect 8628 21904 8634 21916
rect 8665 21913 8677 21916
rect 8711 21913 8723 21947
rect 8665 21907 8723 21913
rect 9214 21904 9220 21956
rect 9272 21904 9278 21956
rect 6178 21876 6184 21888
rect 5552 21848 6184 21876
rect 6178 21836 6184 21848
rect 6236 21836 6242 21888
rect 6365 21879 6423 21885
rect 6365 21845 6377 21879
rect 6411 21876 6423 21879
rect 6546 21876 6552 21888
rect 6411 21848 6552 21876
rect 6411 21845 6423 21848
rect 6365 21839 6423 21845
rect 6546 21836 6552 21848
rect 6604 21836 6610 21888
rect 7098 21836 7104 21888
rect 7156 21876 7162 21888
rect 7561 21879 7619 21885
rect 7561 21876 7573 21879
rect 7156 21848 7573 21876
rect 7156 21836 7162 21848
rect 7561 21845 7573 21848
rect 7607 21845 7619 21879
rect 7561 21839 7619 21845
rect 8386 21836 8392 21888
rect 8444 21836 8450 21888
rect 9030 21836 9036 21888
rect 9088 21836 9094 21888
rect 9398 21836 9404 21888
rect 9456 21876 9462 21888
rect 9784 21876 9812 21975
rect 14274 21972 14280 22024
rect 14332 21972 14338 22024
rect 16960 22021 16988 22052
rect 17862 22040 17868 22052
rect 17920 22040 17926 22092
rect 18437 22083 18495 22089
rect 18437 22049 18449 22083
rect 18483 22080 18495 22083
rect 18598 22080 18604 22092
rect 18483 22052 18604 22080
rect 18483 22049 18495 22052
rect 18437 22043 18495 22049
rect 18598 22040 18604 22052
rect 18656 22040 18662 22092
rect 18690 22040 18696 22092
rect 18748 22040 18754 22092
rect 19150 22040 19156 22092
rect 19208 22080 19214 22092
rect 19797 22083 19855 22089
rect 19797 22080 19809 22083
rect 19208 22052 19809 22080
rect 19208 22040 19214 22052
rect 19797 22049 19809 22052
rect 19843 22049 19855 22083
rect 19797 22043 19855 22049
rect 19889 22083 19947 22089
rect 19889 22049 19901 22083
rect 19935 22049 19947 22083
rect 19889 22043 19947 22049
rect 16945 22015 17003 22021
rect 16945 21981 16957 22015
rect 16991 21981 17003 22015
rect 16945 21975 17003 21981
rect 17126 21972 17132 22024
rect 17184 22012 17190 22024
rect 17310 22012 17316 22024
rect 17184 21984 17316 22012
rect 17184 21972 17190 21984
rect 17310 21972 17316 21984
rect 17368 21972 17374 22024
rect 18966 21972 18972 22024
rect 19024 21972 19030 22024
rect 19061 22015 19119 22021
rect 19061 21981 19073 22015
rect 19107 21981 19119 22015
rect 19904 22012 19932 22043
rect 19978 22040 19984 22092
rect 20036 22040 20042 22092
rect 20162 22040 20168 22092
rect 20220 22040 20226 22092
rect 20254 22040 20260 22092
rect 20312 22080 20318 22092
rect 20824 22089 20852 22120
rect 21542 22089 21548 22092
rect 20441 22083 20499 22089
rect 20441 22080 20453 22083
rect 20312 22052 20453 22080
rect 20312 22040 20318 22052
rect 20441 22049 20453 22052
rect 20487 22049 20499 22083
rect 20441 22043 20499 22049
rect 20625 22083 20683 22089
rect 20625 22049 20637 22083
rect 20671 22049 20683 22083
rect 20625 22043 20683 22049
rect 20809 22083 20867 22089
rect 20809 22049 20821 22083
rect 20855 22049 20867 22083
rect 20809 22043 20867 22049
rect 21085 22083 21143 22089
rect 21085 22049 21097 22083
rect 21131 22049 21143 22083
rect 21536 22080 21548 22089
rect 21503 22052 21548 22080
rect 21085 22043 21143 22049
rect 21536 22043 21548 22052
rect 20346 22012 20352 22024
rect 19904 21984 20352 22012
rect 19061 21975 19119 21981
rect 9858 21904 9864 21956
rect 9916 21944 9922 21956
rect 11057 21947 11115 21953
rect 11057 21944 11069 21947
rect 9916 21916 11069 21944
rect 9916 21904 9922 21916
rect 11057 21913 11069 21916
rect 11103 21913 11115 21947
rect 11057 21907 11115 21913
rect 12710 21904 12716 21956
rect 12768 21944 12774 21956
rect 13081 21947 13139 21953
rect 13081 21944 13093 21947
rect 12768 21916 13093 21944
rect 12768 21904 12774 21916
rect 13081 21913 13093 21916
rect 13127 21913 13139 21947
rect 13081 21907 13139 21913
rect 13262 21904 13268 21956
rect 13320 21944 13326 21956
rect 13357 21947 13415 21953
rect 13357 21944 13369 21947
rect 13320 21916 13369 21944
rect 13320 21904 13326 21916
rect 13357 21913 13369 21916
rect 13403 21913 13415 21947
rect 13357 21907 13415 21913
rect 15289 21947 15347 21953
rect 15289 21913 15301 21947
rect 15335 21944 15347 21947
rect 19076 21944 19104 21975
rect 20346 21972 20352 21984
rect 20404 21972 20410 22024
rect 20530 21972 20536 22024
rect 20588 22012 20594 22024
rect 20640 22012 20668 22043
rect 20588 21984 20668 22012
rect 20588 21972 20594 21984
rect 19613 21947 19671 21953
rect 19613 21944 19625 21947
rect 15335 21916 17356 21944
rect 19076 21916 19625 21944
rect 15335 21913 15347 21916
rect 15289 21907 15347 21913
rect 9456 21848 9812 21876
rect 10137 21879 10195 21885
rect 9456 21836 9462 21848
rect 10137 21845 10149 21879
rect 10183 21876 10195 21879
rect 10413 21879 10471 21885
rect 10413 21876 10425 21879
rect 10183 21848 10425 21876
rect 10183 21845 10195 21848
rect 10137 21839 10195 21845
rect 10413 21845 10425 21848
rect 10459 21845 10471 21879
rect 10413 21839 10471 21845
rect 12066 21836 12072 21888
rect 12124 21836 12130 21888
rect 12526 21836 12532 21888
rect 12584 21836 12590 21888
rect 12618 21836 12624 21888
rect 12676 21876 12682 21888
rect 13633 21879 13691 21885
rect 13633 21876 13645 21879
rect 12676 21848 13645 21876
rect 12676 21836 12682 21848
rect 13633 21845 13645 21848
rect 13679 21845 13691 21879
rect 13633 21839 13691 21845
rect 14553 21879 14611 21885
rect 14553 21845 14565 21879
rect 14599 21876 14611 21879
rect 15010 21876 15016 21888
rect 14599 21848 15016 21876
rect 14599 21845 14611 21848
rect 14553 21839 14611 21845
rect 15010 21836 15016 21848
rect 15068 21836 15074 21888
rect 15841 21879 15899 21885
rect 15841 21845 15853 21879
rect 15887 21876 15899 21879
rect 16390 21876 16396 21888
rect 15887 21848 16396 21876
rect 15887 21845 15899 21848
rect 15841 21839 15899 21845
rect 16390 21836 16396 21848
rect 16448 21836 16454 21888
rect 16485 21879 16543 21885
rect 16485 21845 16497 21879
rect 16531 21876 16543 21879
rect 16850 21876 16856 21888
rect 16531 21848 16856 21876
rect 16531 21845 16543 21848
rect 16485 21839 16543 21845
rect 16850 21836 16856 21848
rect 16908 21836 16914 21888
rect 17328 21876 17356 21916
rect 19613 21913 19625 21916
rect 19659 21913 19671 21947
rect 19613 21907 19671 21913
rect 19794 21904 19800 21956
rect 19852 21944 19858 21956
rect 21100 21944 21128 22043
rect 21542 22040 21548 22043
rect 21600 22040 21606 22092
rect 21652 22080 21680 22120
rect 22922 22108 22928 22160
rect 22980 22108 22986 22160
rect 21652 22052 22692 22080
rect 21266 21972 21272 22024
rect 21324 21972 21330 22024
rect 22664 21953 22692 22052
rect 19852 21916 21128 21944
rect 22649 21947 22707 21953
rect 19852 21904 19858 21916
rect 22649 21913 22661 21947
rect 22695 21913 22707 21947
rect 22649 21907 22707 21913
rect 19426 21876 19432 21888
rect 17328 21848 19432 21876
rect 19426 21836 19432 21848
rect 19484 21836 19490 21888
rect 19521 21879 19579 21885
rect 19521 21845 19533 21879
rect 19567 21876 19579 21879
rect 20806 21876 20812 21888
rect 19567 21848 20812 21876
rect 19567 21845 19579 21848
rect 19521 21839 19579 21845
rect 20806 21836 20812 21848
rect 20864 21836 20870 21888
rect 20901 21879 20959 21885
rect 20901 21845 20913 21879
rect 20947 21876 20959 21879
rect 21174 21876 21180 21888
rect 20947 21848 21180 21876
rect 20947 21845 20959 21848
rect 20901 21839 20959 21845
rect 21174 21836 21180 21848
rect 21232 21836 21238 21888
rect 21266 21836 21272 21888
rect 21324 21876 21330 21888
rect 22186 21876 22192 21888
rect 21324 21848 22192 21876
rect 21324 21836 21330 21848
rect 22186 21836 22192 21848
rect 22244 21836 22250 21888
rect 22278 21836 22284 21888
rect 22336 21876 22342 21888
rect 22833 21879 22891 21885
rect 22833 21876 22845 21879
rect 22336 21848 22845 21876
rect 22336 21836 22342 21848
rect 22833 21845 22845 21848
rect 22879 21845 22891 21879
rect 22833 21839 22891 21845
rect 552 21786 23368 21808
rect 552 21734 1366 21786
rect 1418 21734 1430 21786
rect 1482 21734 1494 21786
rect 1546 21734 1558 21786
rect 1610 21734 1622 21786
rect 1674 21734 1686 21786
rect 1738 21734 7366 21786
rect 7418 21734 7430 21786
rect 7482 21734 7494 21786
rect 7546 21734 7558 21786
rect 7610 21734 7622 21786
rect 7674 21734 7686 21786
rect 7738 21734 13366 21786
rect 13418 21734 13430 21786
rect 13482 21734 13494 21786
rect 13546 21734 13558 21786
rect 13610 21734 13622 21786
rect 13674 21734 13686 21786
rect 13738 21734 19366 21786
rect 19418 21734 19430 21786
rect 19482 21734 19494 21786
rect 19546 21734 19558 21786
rect 19610 21734 19622 21786
rect 19674 21734 19686 21786
rect 19738 21734 23368 21786
rect 552 21712 23368 21734
rect 1854 21632 1860 21684
rect 1912 21672 1918 21684
rect 2869 21675 2927 21681
rect 2869 21672 2881 21675
rect 1912 21644 2881 21672
rect 1912 21632 1918 21644
rect 2869 21641 2881 21644
rect 2915 21641 2927 21675
rect 2869 21635 2927 21641
rect 3418 21632 3424 21684
rect 3476 21632 3482 21684
rect 5166 21632 5172 21684
rect 5224 21672 5230 21684
rect 5902 21672 5908 21684
rect 5224 21644 5908 21672
rect 5224 21632 5230 21644
rect 5902 21632 5908 21644
rect 5960 21632 5966 21684
rect 6365 21675 6423 21681
rect 6365 21641 6377 21675
rect 6411 21672 6423 21675
rect 6822 21672 6828 21684
rect 6411 21644 6828 21672
rect 6411 21641 6423 21644
rect 6365 21635 6423 21641
rect 3234 21604 3240 21616
rect 2240 21576 3240 21604
rect 2240 21545 2268 21576
rect 3234 21564 3240 21576
rect 3292 21564 3298 21616
rect 3436 21604 3464 21632
rect 4341 21607 4399 21613
rect 3436 21576 4108 21604
rect 2225 21539 2283 21545
rect 2225 21505 2237 21539
rect 2271 21505 2283 21539
rect 2225 21499 2283 21505
rect 2774 21496 2780 21548
rect 2832 21496 2838 21548
rect 2958 21496 2964 21548
rect 3016 21536 3022 21548
rect 4080 21545 4108 21576
rect 4341 21573 4353 21607
rect 4387 21604 4399 21607
rect 5258 21604 5264 21616
rect 4387 21576 5264 21604
rect 4387 21573 4399 21576
rect 4341 21567 4399 21573
rect 5258 21564 5264 21576
rect 5316 21564 5322 21616
rect 3697 21539 3755 21545
rect 3697 21536 3709 21539
rect 3016 21508 3709 21536
rect 3016 21496 3022 21508
rect 3697 21505 3709 21508
rect 3743 21505 3755 21539
rect 3697 21499 3755 21505
rect 4065 21539 4123 21545
rect 4065 21505 4077 21539
rect 4111 21536 4123 21539
rect 4890 21536 4896 21548
rect 4111 21508 4896 21536
rect 4111 21505 4123 21508
rect 4065 21499 4123 21505
rect 1946 21428 1952 21480
rect 2004 21477 2010 21480
rect 2004 21468 2016 21477
rect 2004 21440 2049 21468
rect 2004 21431 2016 21440
rect 2004 21428 2010 21431
rect 2498 21428 2504 21480
rect 2556 21428 2562 21480
rect 3053 21471 3111 21477
rect 3053 21437 3065 21471
rect 3099 21468 3111 21471
rect 3142 21468 3148 21480
rect 3099 21440 3148 21468
rect 3099 21437 3111 21440
rect 3053 21431 3111 21437
rect 3142 21428 3148 21440
rect 3200 21468 3206 21480
rect 3200 21440 3648 21468
rect 3200 21428 3206 21440
rect 2130 21360 2136 21412
rect 2188 21400 2194 21412
rect 2866 21400 2872 21412
rect 2188 21372 2872 21400
rect 2188 21360 2194 21372
rect 2866 21360 2872 21372
rect 2924 21360 2930 21412
rect 3326 21360 3332 21412
rect 3384 21409 3390 21412
rect 3620 21409 3648 21440
rect 3878 21428 3884 21480
rect 3936 21428 3942 21480
rect 4246 21428 4252 21480
rect 4304 21468 4310 21480
rect 4724 21477 4752 21508
rect 4890 21496 4896 21508
rect 4948 21496 4954 21548
rect 6380 21536 6408 21635
rect 6822 21632 6828 21644
rect 6880 21672 6886 21684
rect 6880 21644 7328 21672
rect 6880 21632 6886 21644
rect 6638 21564 6644 21616
rect 6696 21604 6702 21616
rect 7193 21607 7251 21613
rect 7193 21604 7205 21607
rect 6696 21576 7205 21604
rect 6696 21564 6702 21576
rect 7193 21573 7205 21576
rect 7239 21573 7251 21607
rect 7300 21604 7328 21644
rect 7466 21632 7472 21684
rect 7524 21632 7530 21684
rect 8846 21632 8852 21684
rect 8904 21672 8910 21684
rect 9033 21675 9091 21681
rect 9033 21672 9045 21675
rect 8904 21644 9045 21672
rect 8904 21632 8910 21644
rect 9033 21641 9045 21644
rect 9079 21641 9091 21675
rect 9033 21635 9091 21641
rect 9416 21644 9628 21672
rect 8018 21604 8024 21616
rect 7300 21576 8024 21604
rect 7193 21567 7251 21573
rect 8018 21564 8024 21576
rect 8076 21564 8082 21616
rect 8757 21607 8815 21613
rect 8757 21573 8769 21607
rect 8803 21604 8815 21607
rect 9306 21604 9312 21616
rect 8803 21576 9312 21604
rect 8803 21573 8815 21576
rect 8757 21567 8815 21573
rect 9306 21564 9312 21576
rect 9364 21564 9370 21616
rect 5000 21508 5856 21536
rect 4525 21471 4583 21477
rect 4525 21468 4537 21471
rect 4304 21440 4537 21468
rect 4304 21428 4310 21440
rect 4525 21437 4537 21440
rect 4571 21437 4583 21471
rect 4525 21431 4583 21437
rect 4709 21471 4767 21477
rect 4709 21437 4721 21471
rect 4755 21437 4767 21471
rect 5000 21468 5028 21508
rect 4709 21431 4767 21437
rect 4816 21440 5028 21468
rect 3384 21403 3447 21409
rect 3384 21369 3401 21403
rect 3435 21369 3447 21403
rect 3384 21363 3447 21369
rect 3605 21403 3663 21409
rect 3605 21369 3617 21403
rect 3651 21369 3663 21403
rect 3605 21363 3663 21369
rect 3384 21360 3390 21363
rect 845 21335 903 21341
rect 845 21301 857 21335
rect 891 21332 903 21335
rect 2038 21332 2044 21344
rect 891 21304 2044 21332
rect 891 21301 903 21304
rect 845 21295 903 21301
rect 2038 21292 2044 21304
rect 2096 21292 2102 21344
rect 2590 21292 2596 21344
rect 2648 21332 2654 21344
rect 2685 21335 2743 21341
rect 2685 21332 2697 21335
rect 2648 21304 2697 21332
rect 2648 21292 2654 21304
rect 2685 21301 2697 21304
rect 2731 21301 2743 21335
rect 2685 21295 2743 21301
rect 2958 21292 2964 21344
rect 3016 21332 3022 21344
rect 3237 21335 3295 21341
rect 3237 21332 3249 21335
rect 3016 21304 3249 21332
rect 3016 21292 3022 21304
rect 3237 21301 3249 21304
rect 3283 21301 3295 21335
rect 3620 21332 3648 21363
rect 4617 21335 4675 21341
rect 4617 21332 4629 21335
rect 3620 21304 4629 21332
rect 3237 21295 3295 21301
rect 4617 21301 4629 21304
rect 4663 21332 4675 21335
rect 4816 21332 4844 21440
rect 5166 21428 5172 21480
rect 5224 21428 5230 21480
rect 5445 21471 5503 21477
rect 5445 21437 5457 21471
rect 5491 21468 5503 21471
rect 5626 21468 5632 21480
rect 5491 21440 5632 21468
rect 5491 21437 5503 21440
rect 5445 21431 5503 21437
rect 5626 21428 5632 21440
rect 5684 21428 5690 21480
rect 5828 21477 5856 21508
rect 6104 21508 6408 21536
rect 6779 21539 6837 21545
rect 6104 21477 6132 21508
rect 6779 21505 6791 21539
rect 6825 21536 6837 21539
rect 7926 21536 7932 21548
rect 6825 21508 7932 21536
rect 6825 21505 6837 21508
rect 6779 21499 6837 21505
rect 7926 21496 7932 21508
rect 7984 21496 7990 21548
rect 8312 21508 8800 21536
rect 5813 21471 5871 21477
rect 5813 21437 5825 21471
rect 5859 21437 5871 21471
rect 5813 21431 5871 21437
rect 6089 21471 6147 21477
rect 6089 21437 6101 21471
rect 6135 21437 6147 21471
rect 6089 21431 6147 21437
rect 6178 21428 6184 21480
rect 6236 21470 6242 21480
rect 6236 21442 6316 21470
rect 6236 21428 6242 21442
rect 6288 21400 6316 21442
rect 6638 21428 6644 21480
rect 6696 21428 6702 21480
rect 6914 21428 6920 21480
rect 6972 21428 6978 21480
rect 7006 21428 7012 21480
rect 7064 21428 7070 21480
rect 7101 21471 7159 21477
rect 7101 21437 7113 21471
rect 7147 21468 7159 21471
rect 7190 21468 7196 21480
rect 7147 21440 7196 21468
rect 7147 21437 7159 21440
rect 7101 21431 7159 21437
rect 7190 21428 7196 21440
rect 7248 21428 7254 21480
rect 7374 21428 7380 21480
rect 7432 21428 7438 21480
rect 7469 21471 7527 21477
rect 7469 21437 7481 21471
rect 7515 21437 7527 21471
rect 7469 21431 7527 21437
rect 7484 21400 7512 21431
rect 7650 21428 7656 21480
rect 7708 21468 7714 21480
rect 8312 21468 8340 21508
rect 7708 21440 8340 21468
rect 7708 21428 7714 21440
rect 8386 21428 8392 21480
rect 8444 21468 8450 21480
rect 8573 21471 8631 21477
rect 8573 21468 8585 21471
rect 8444 21440 8585 21468
rect 8444 21428 8450 21440
rect 8573 21437 8585 21440
rect 8619 21437 8631 21471
rect 8573 21431 8631 21437
rect 8665 21471 8723 21477
rect 8665 21437 8677 21471
rect 8711 21437 8723 21471
rect 8665 21431 8723 21437
rect 8680 21400 8708 21431
rect 6288 21372 7512 21400
rect 8312 21372 8708 21400
rect 8772 21400 8800 21508
rect 8846 21496 8852 21548
rect 8904 21536 8910 21548
rect 9416 21536 9444 21644
rect 9490 21564 9496 21616
rect 9548 21564 9554 21616
rect 9600 21604 9628 21644
rect 10042 21632 10048 21684
rect 10100 21672 10106 21684
rect 10137 21675 10195 21681
rect 10137 21672 10149 21675
rect 10100 21644 10149 21672
rect 10100 21632 10106 21644
rect 10137 21641 10149 21644
rect 10183 21641 10195 21675
rect 10137 21635 10195 21641
rect 14001 21675 14059 21681
rect 14001 21641 14013 21675
rect 14047 21672 14059 21675
rect 14182 21672 14188 21684
rect 14047 21644 14188 21672
rect 14047 21641 14059 21644
rect 14001 21635 14059 21641
rect 14182 21632 14188 21644
rect 14240 21632 14246 21684
rect 14829 21675 14887 21681
rect 14829 21641 14841 21675
rect 14875 21672 14887 21675
rect 15378 21672 15384 21684
rect 14875 21644 15384 21672
rect 14875 21641 14887 21644
rect 14829 21635 14887 21641
rect 15378 21632 15384 21644
rect 15436 21632 15442 21684
rect 15746 21632 15752 21684
rect 15804 21672 15810 21684
rect 18141 21675 18199 21681
rect 18141 21672 18153 21675
rect 15804 21644 18153 21672
rect 15804 21632 15810 21644
rect 18141 21641 18153 21644
rect 18187 21641 18199 21675
rect 18141 21635 18199 21641
rect 19242 21632 19248 21684
rect 19300 21632 19306 21684
rect 19518 21632 19524 21684
rect 19576 21672 19582 21684
rect 19889 21675 19947 21681
rect 19889 21672 19901 21675
rect 19576 21644 19901 21672
rect 19576 21632 19582 21644
rect 19889 21641 19901 21644
rect 19935 21641 19947 21675
rect 20533 21675 20591 21681
rect 20533 21672 20545 21675
rect 19889 21635 19947 21641
rect 19996 21644 20545 21672
rect 10873 21607 10931 21613
rect 10873 21604 10885 21607
rect 9600 21576 10885 21604
rect 10873 21573 10885 21576
rect 10919 21573 10931 21607
rect 10873 21567 10931 21573
rect 13357 21607 13415 21613
rect 13357 21573 13369 21607
rect 13403 21604 13415 21607
rect 16022 21604 16028 21616
rect 13403 21576 16028 21604
rect 13403 21573 13415 21576
rect 13357 21567 13415 21573
rect 16022 21564 16028 21576
rect 16080 21564 16086 21616
rect 19260 21604 19288 21632
rect 19996 21604 20024 21644
rect 20533 21641 20545 21644
rect 20579 21641 20591 21675
rect 20533 21635 20591 21641
rect 20806 21632 20812 21684
rect 20864 21672 20870 21684
rect 20864 21644 23060 21672
rect 20864 21632 20870 21644
rect 19260 21576 20024 21604
rect 20162 21564 20168 21616
rect 20220 21604 20226 21616
rect 21082 21604 21088 21616
rect 20220 21576 21088 21604
rect 20220 21564 20226 21576
rect 8904 21508 9444 21536
rect 9508 21536 9536 21564
rect 9508 21508 10640 21536
rect 8904 21496 8910 21508
rect 8938 21428 8944 21480
rect 8996 21468 9002 21480
rect 9217 21471 9275 21477
rect 9217 21468 9229 21471
rect 8996 21440 9229 21468
rect 8996 21428 9002 21440
rect 9217 21437 9229 21440
rect 9263 21437 9275 21471
rect 9217 21431 9275 21437
rect 9306 21428 9312 21480
rect 9364 21428 9370 21480
rect 9416 21468 9444 21508
rect 9769 21471 9827 21477
rect 9769 21468 9781 21471
rect 9416 21440 9781 21468
rect 9769 21437 9781 21440
rect 9815 21437 9827 21471
rect 9769 21431 9827 21437
rect 9858 21428 9864 21480
rect 9916 21428 9922 21480
rect 10060 21477 10088 21508
rect 10045 21471 10103 21477
rect 10045 21437 10057 21471
rect 10091 21437 10103 21471
rect 10045 21431 10103 21437
rect 10229 21471 10287 21477
rect 10229 21437 10241 21471
rect 10275 21468 10287 21471
rect 10318 21468 10324 21480
rect 10275 21440 10324 21468
rect 10275 21437 10287 21440
rect 10229 21431 10287 21437
rect 9876 21400 9904 21428
rect 10244 21400 10272 21431
rect 10318 21428 10324 21440
rect 10376 21428 10382 21480
rect 10612 21477 10640 21508
rect 11974 21496 11980 21548
rect 12032 21536 12038 21548
rect 12529 21539 12587 21545
rect 12529 21536 12541 21539
rect 12032 21508 12541 21536
rect 12032 21496 12038 21508
rect 12529 21505 12541 21508
rect 12575 21505 12587 21539
rect 15286 21536 15292 21548
rect 12529 21499 12587 21505
rect 14660 21508 15292 21536
rect 10597 21471 10655 21477
rect 10597 21437 10609 21471
rect 10643 21468 10655 21471
rect 10778 21468 10784 21480
rect 10643 21440 10784 21468
rect 10643 21437 10655 21440
rect 10597 21431 10655 21437
rect 10778 21428 10784 21440
rect 10836 21428 10842 21480
rect 11057 21471 11115 21477
rect 11057 21437 11069 21471
rect 11103 21468 11115 21471
rect 11422 21468 11428 21480
rect 11103 21440 11428 21468
rect 11103 21437 11115 21440
rect 11057 21431 11115 21437
rect 11422 21428 11428 21440
rect 11480 21428 11486 21480
rect 11514 21428 11520 21480
rect 11572 21468 11578 21480
rect 11609 21471 11667 21477
rect 11609 21468 11621 21471
rect 11572 21440 11621 21468
rect 11572 21428 11578 21440
rect 11609 21437 11621 21440
rect 11655 21437 11667 21471
rect 11609 21431 11667 21437
rect 11885 21471 11943 21477
rect 11885 21437 11897 21471
rect 11931 21437 11943 21471
rect 11885 21431 11943 21437
rect 12437 21471 12495 21477
rect 12437 21437 12449 21471
rect 12483 21468 12495 21471
rect 12618 21468 12624 21480
rect 12483 21440 12624 21468
rect 12483 21437 12495 21440
rect 12437 21431 12495 21437
rect 8772 21372 9904 21400
rect 9968 21372 10272 21400
rect 11900 21400 11928 21431
rect 12618 21428 12624 21440
rect 12676 21428 12682 21480
rect 13170 21428 13176 21480
rect 13228 21428 13234 21480
rect 13725 21471 13783 21477
rect 13725 21437 13737 21471
rect 13771 21468 13783 21471
rect 13771 21440 14044 21468
rect 13771 21437 13783 21440
rect 13725 21431 13783 21437
rect 11974 21400 11980 21412
rect 11900 21372 11980 21400
rect 8312 21344 8340 21372
rect 4663 21304 4844 21332
rect 4663 21301 4675 21304
rect 4617 21295 4675 21301
rect 4890 21292 4896 21344
rect 4948 21292 4954 21344
rect 5074 21292 5080 21344
rect 5132 21292 5138 21344
rect 5629 21335 5687 21341
rect 5629 21301 5641 21335
rect 5675 21332 5687 21335
rect 5810 21332 5816 21344
rect 5675 21304 5816 21332
rect 5675 21301 5687 21304
rect 5629 21295 5687 21301
rect 5810 21292 5816 21304
rect 5868 21292 5874 21344
rect 5902 21292 5908 21344
rect 5960 21332 5966 21344
rect 7466 21332 7472 21344
rect 5960 21304 7472 21332
rect 5960 21292 5966 21304
rect 7466 21292 7472 21304
rect 7524 21292 7530 21344
rect 8294 21292 8300 21344
rect 8352 21292 8358 21344
rect 8389 21335 8447 21341
rect 8389 21301 8401 21335
rect 8435 21332 8447 21335
rect 9674 21332 9680 21344
rect 8435 21304 9680 21332
rect 8435 21301 8447 21304
rect 8389 21295 8447 21301
rect 9674 21292 9680 21304
rect 9732 21292 9738 21344
rect 9858 21292 9864 21344
rect 9916 21332 9922 21344
rect 9968 21341 9996 21372
rect 11974 21360 11980 21372
rect 12032 21400 12038 21412
rect 12032 21372 12434 21400
rect 12032 21360 12038 21372
rect 9953 21335 10011 21341
rect 9953 21332 9965 21335
rect 9916 21304 9965 21332
rect 9916 21292 9922 21304
rect 9953 21301 9965 21304
rect 9999 21301 10011 21335
rect 9953 21295 10011 21301
rect 10689 21335 10747 21341
rect 10689 21301 10701 21335
rect 10735 21332 10747 21335
rect 10778 21332 10784 21344
rect 10735 21304 10784 21332
rect 10735 21301 10747 21304
rect 10689 21295 10747 21301
rect 10778 21292 10784 21304
rect 10836 21292 10842 21344
rect 11422 21292 11428 21344
rect 11480 21292 11486 21344
rect 11698 21292 11704 21344
rect 11756 21292 11762 21344
rect 12406 21332 12434 21372
rect 12710 21332 12716 21344
rect 12406 21304 12716 21332
rect 12710 21292 12716 21304
rect 12768 21292 12774 21344
rect 12802 21292 12808 21344
rect 12860 21292 12866 21344
rect 13906 21292 13912 21344
rect 13964 21292 13970 21344
rect 14016 21332 14044 21440
rect 14182 21428 14188 21480
rect 14240 21428 14246 21480
rect 14274 21428 14280 21480
rect 14332 21428 14338 21480
rect 14366 21428 14372 21480
rect 14424 21428 14430 21480
rect 14458 21428 14464 21480
rect 14516 21428 14522 21480
rect 14660 21477 14688 21508
rect 15286 21496 15292 21508
rect 15344 21536 15350 21548
rect 15562 21536 15568 21548
rect 15344 21508 15568 21536
rect 15344 21496 15350 21508
rect 15562 21496 15568 21508
rect 15620 21496 15626 21548
rect 16761 21539 16819 21545
rect 16761 21505 16773 21539
rect 16807 21536 16819 21539
rect 16807 21508 16876 21536
rect 16807 21505 16819 21508
rect 16761 21499 16819 21505
rect 14645 21471 14703 21477
rect 14645 21437 14657 21471
rect 14691 21437 14703 21471
rect 14645 21431 14703 21437
rect 14734 21428 14740 21480
rect 14792 21468 14798 21480
rect 14829 21471 14887 21477
rect 14829 21468 14841 21471
rect 14792 21440 14841 21468
rect 14792 21428 14798 21440
rect 14829 21437 14841 21440
rect 14875 21437 14887 21471
rect 14829 21431 14887 21437
rect 15212 21440 16620 21468
rect 15212 21412 15240 21440
rect 14090 21360 14096 21412
rect 14148 21400 14154 21412
rect 14921 21403 14979 21409
rect 14921 21400 14933 21403
rect 14148 21372 14933 21400
rect 14148 21360 14154 21372
rect 14921 21369 14933 21372
rect 14967 21400 14979 21403
rect 15194 21400 15200 21412
rect 14967 21372 15200 21400
rect 14967 21369 14979 21372
rect 14921 21363 14979 21369
rect 15194 21360 15200 21372
rect 15252 21360 15258 21412
rect 15378 21360 15384 21412
rect 15436 21400 15442 21412
rect 15838 21400 15844 21412
rect 15436 21372 15844 21400
rect 15436 21360 15442 21372
rect 15838 21360 15844 21372
rect 15896 21360 15902 21412
rect 16592 21400 16620 21440
rect 16666 21428 16672 21480
rect 16724 21428 16730 21480
rect 16848 21468 16876 21508
rect 19058 21496 19064 21548
rect 19116 21536 19122 21548
rect 19153 21539 19211 21545
rect 19153 21536 19165 21539
rect 19116 21508 19165 21536
rect 19116 21496 19122 21508
rect 19153 21505 19165 21508
rect 19199 21505 19211 21539
rect 19153 21499 19211 21505
rect 19242 21496 19248 21548
rect 19300 21536 19306 21548
rect 19300 21508 20208 21536
rect 19300 21496 19306 21508
rect 20180 21480 20208 21508
rect 16776 21440 16876 21468
rect 17017 21471 17075 21477
rect 16776 21400 16804 21440
rect 17017 21437 17029 21471
rect 17063 21437 17075 21471
rect 17017 21431 17075 21437
rect 18325 21471 18383 21477
rect 18325 21437 18337 21471
rect 18371 21468 18383 21471
rect 19886 21468 19892 21480
rect 18371 21464 19104 21468
rect 19168 21464 19892 21468
rect 18371 21440 19892 21464
rect 18371 21437 18383 21440
rect 18325 21431 18383 21437
rect 19076 21436 19196 21440
rect 17032 21400 17060 21431
rect 19886 21428 19892 21440
rect 19944 21428 19950 21480
rect 20070 21428 20076 21480
rect 20128 21428 20134 21480
rect 20162 21428 20168 21480
rect 20220 21428 20226 21480
rect 20272 21477 20300 21576
rect 21082 21564 21088 21576
rect 21140 21564 21146 21616
rect 21361 21607 21419 21613
rect 21361 21573 21373 21607
rect 21407 21604 21419 21607
rect 21450 21604 21456 21616
rect 21407 21576 21456 21604
rect 21407 21573 21419 21576
rect 21361 21567 21419 21573
rect 21450 21564 21456 21576
rect 21508 21564 21514 21616
rect 22741 21539 22799 21545
rect 20640 21508 20852 21536
rect 20257 21471 20315 21477
rect 20257 21437 20269 21471
rect 20303 21437 20315 21471
rect 20257 21431 20315 21437
rect 20441 21471 20499 21477
rect 20441 21437 20453 21471
rect 20487 21437 20499 21471
rect 20441 21431 20499 21437
rect 16592 21372 16804 21400
rect 16848 21372 17060 21400
rect 16114 21332 16120 21344
rect 14016 21304 16120 21332
rect 16114 21292 16120 21304
rect 16172 21292 16178 21344
rect 16390 21292 16396 21344
rect 16448 21332 16454 21344
rect 16848 21332 16876 21372
rect 17770 21360 17776 21412
rect 17828 21400 17834 21412
rect 18785 21403 18843 21409
rect 18785 21400 18797 21403
rect 17828 21372 18797 21400
rect 17828 21360 17834 21372
rect 18785 21369 18797 21372
rect 18831 21400 18843 21403
rect 19242 21400 19248 21412
rect 18831 21372 19248 21400
rect 18831 21369 18843 21372
rect 18785 21363 18843 21369
rect 19242 21360 19248 21372
rect 19300 21360 19306 21412
rect 19337 21403 19395 21409
rect 19337 21369 19349 21403
rect 19383 21400 19395 21403
rect 19518 21400 19524 21412
rect 19383 21372 19524 21400
rect 19383 21369 19395 21372
rect 19337 21363 19395 21369
rect 19518 21360 19524 21372
rect 19576 21360 19582 21412
rect 19702 21360 19708 21412
rect 19760 21400 19766 21412
rect 19760 21372 19840 21400
rect 19760 21360 19766 21372
rect 16448 21304 16876 21332
rect 16448 21292 16454 21304
rect 16942 21292 16948 21344
rect 17000 21332 17006 21344
rect 17494 21332 17500 21344
rect 17000 21304 17500 21332
rect 17000 21292 17006 21304
rect 17494 21292 17500 21304
rect 17552 21292 17558 21344
rect 18414 21292 18420 21344
rect 18472 21292 18478 21344
rect 18874 21292 18880 21344
rect 18932 21292 18938 21344
rect 19426 21292 19432 21344
rect 19484 21292 19490 21344
rect 19812 21341 19840 21372
rect 19978 21360 19984 21412
rect 20036 21400 20042 21412
rect 20456 21400 20484 21431
rect 20530 21428 20536 21480
rect 20588 21468 20594 21480
rect 20640 21468 20668 21508
rect 20824 21484 20852 21508
rect 22741 21505 22753 21539
rect 22787 21536 22799 21539
rect 22830 21536 22836 21548
rect 22787 21508 22836 21536
rect 22787 21505 22799 21508
rect 22741 21499 22799 21505
rect 22830 21496 22836 21508
rect 22888 21496 22894 21548
rect 20824 21477 20944 21484
rect 21100 21477 21220 21484
rect 20588 21440 20668 21468
rect 20717 21471 20775 21477
rect 20588 21428 20594 21440
rect 20717 21437 20729 21471
rect 20763 21437 20775 21471
rect 20824 21471 20959 21477
rect 20824 21456 20913 21471
rect 20717 21431 20775 21437
rect 20901 21437 20913 21456
rect 20947 21437 20959 21471
rect 20901 21431 20959 21437
rect 21085 21471 21220 21477
rect 21085 21437 21097 21471
rect 21131 21468 21220 21471
rect 21358 21468 21364 21480
rect 21131 21456 21364 21468
rect 21131 21437 21143 21456
rect 21192 21440 21364 21456
rect 21085 21431 21143 21437
rect 20036 21372 20484 21400
rect 20036 21360 20042 21372
rect 19797 21335 19855 21341
rect 19797 21301 19809 21335
rect 19843 21301 19855 21335
rect 20732 21332 20760 21431
rect 21358 21428 21364 21440
rect 21416 21428 21422 21480
rect 23032 21477 23060 21644
rect 23017 21471 23075 21477
rect 23017 21437 23029 21471
rect 23063 21437 23075 21471
rect 23017 21431 23075 21437
rect 20806 21360 20812 21412
rect 20864 21360 20870 21412
rect 22002 21400 22008 21412
rect 21192 21372 22008 21400
rect 21192 21332 21220 21372
rect 22002 21360 22008 21372
rect 22060 21360 22066 21412
rect 22278 21360 22284 21412
rect 22336 21400 22342 21412
rect 22474 21403 22532 21409
rect 22474 21400 22486 21403
rect 22336 21372 22486 21400
rect 22336 21360 22342 21372
rect 22474 21369 22486 21372
rect 22520 21369 22532 21403
rect 22474 21363 22532 21369
rect 20732 21304 21220 21332
rect 19797 21295 19855 21301
rect 21450 21292 21456 21344
rect 21508 21332 21514 21344
rect 22833 21335 22891 21341
rect 22833 21332 22845 21335
rect 21508 21304 22845 21332
rect 21508 21292 21514 21304
rect 22833 21301 22845 21304
rect 22879 21301 22891 21335
rect 22833 21295 22891 21301
rect 552 21242 23368 21264
rect 552 21190 4366 21242
rect 4418 21190 4430 21242
rect 4482 21190 4494 21242
rect 4546 21190 4558 21242
rect 4610 21190 4622 21242
rect 4674 21190 4686 21242
rect 4738 21190 10366 21242
rect 10418 21190 10430 21242
rect 10482 21190 10494 21242
rect 10546 21190 10558 21242
rect 10610 21190 10622 21242
rect 10674 21190 10686 21242
rect 10738 21190 16366 21242
rect 16418 21190 16430 21242
rect 16482 21190 16494 21242
rect 16546 21190 16558 21242
rect 16610 21190 16622 21242
rect 16674 21190 16686 21242
rect 16738 21190 22366 21242
rect 22418 21190 22430 21242
rect 22482 21190 22494 21242
rect 22546 21190 22558 21242
rect 22610 21190 22622 21242
rect 22674 21190 22686 21242
rect 22738 21190 23368 21242
rect 552 21168 23368 21190
rect 2222 21128 2228 21140
rect 1596 21100 2228 21128
rect 1596 21001 1624 21100
rect 2222 21088 2228 21100
rect 2280 21128 2286 21140
rect 2280 21100 2452 21128
rect 2280 21088 2286 21100
rect 1673 21063 1731 21069
rect 1673 21029 1685 21063
rect 1719 21060 1731 21063
rect 1719 21032 2084 21060
rect 1719 21029 1731 21032
rect 1673 21023 1731 21029
rect 1581 20995 1639 21001
rect 1581 20961 1593 20995
rect 1627 20961 1639 20995
rect 1581 20955 1639 20961
rect 1765 20995 1823 21001
rect 1765 20961 1777 20995
rect 1811 20961 1823 20995
rect 1765 20955 1823 20961
rect 1780 20924 1808 20955
rect 1854 20952 1860 21004
rect 1912 20952 1918 21004
rect 2056 20992 2084 21032
rect 2130 21020 2136 21072
rect 2188 21020 2194 21072
rect 2333 21063 2391 21069
rect 2333 21029 2345 21063
rect 2379 21029 2391 21063
rect 2424 21060 2452 21100
rect 2498 21088 2504 21140
rect 2556 21088 2562 21140
rect 2774 21088 2780 21140
rect 2832 21128 2838 21140
rect 3789 21131 3847 21137
rect 3789 21128 3801 21131
rect 2832 21100 3801 21128
rect 2832 21088 2838 21100
rect 3789 21097 3801 21100
rect 3835 21128 3847 21131
rect 5353 21131 5411 21137
rect 5353 21128 5365 21131
rect 3835 21100 5365 21128
rect 3835 21097 3847 21100
rect 3789 21091 3847 21097
rect 5353 21097 5365 21100
rect 5399 21097 5411 21131
rect 5353 21091 5411 21097
rect 5626 21088 5632 21140
rect 5684 21088 5690 21140
rect 6270 21088 6276 21140
rect 6328 21088 6334 21140
rect 6914 21088 6920 21140
rect 6972 21128 6978 21140
rect 7101 21131 7159 21137
rect 7101 21128 7113 21131
rect 6972 21100 7113 21128
rect 6972 21088 6978 21100
rect 7101 21097 7113 21100
rect 7147 21097 7159 21131
rect 7101 21091 7159 21097
rect 7834 21088 7840 21140
rect 7892 21088 7898 21140
rect 8573 21131 8631 21137
rect 8573 21097 8585 21131
rect 8619 21128 8631 21131
rect 9582 21128 9588 21140
rect 8619 21100 9588 21128
rect 8619 21097 8631 21100
rect 8573 21091 8631 21097
rect 9582 21088 9588 21100
rect 9640 21088 9646 21140
rect 9766 21088 9772 21140
rect 9824 21128 9830 21140
rect 11698 21128 11704 21140
rect 9824 21100 11704 21128
rect 9824 21088 9830 21100
rect 2958 21060 2964 21072
rect 2424 21032 2964 21060
rect 2333 21023 2391 21029
rect 2222 20992 2228 21004
rect 2056 20964 2228 20992
rect 2222 20952 2228 20964
rect 2280 20992 2286 21004
rect 2348 20992 2376 21023
rect 2958 21020 2964 21032
rect 3016 21020 3022 21072
rect 4338 21060 4344 21072
rect 3988 21032 4344 21060
rect 2280 20964 2376 20992
rect 2777 20995 2835 21001
rect 2280 20952 2286 20964
rect 2777 20961 2789 20995
rect 2823 20992 2835 20995
rect 3329 20995 3387 21001
rect 2823 20964 2857 20992
rect 2823 20961 2835 20964
rect 2777 20955 2835 20961
rect 3329 20961 3341 20995
rect 3375 20992 3387 20995
rect 3510 20992 3516 21004
rect 3375 20964 3516 20992
rect 3375 20961 3387 20964
rect 3329 20955 3387 20961
rect 2792 20924 2820 20955
rect 3510 20952 3516 20964
rect 3568 20952 3574 21004
rect 3988 21001 4016 21032
rect 4338 21020 4344 21032
rect 4396 21020 4402 21072
rect 4890 21060 4896 21072
rect 4540 21032 4896 21060
rect 4540 21001 4568 21032
rect 4890 21020 4896 21032
rect 4948 21060 4954 21072
rect 8456 21063 8514 21069
rect 4948 21032 6592 21060
rect 4948 21020 4954 21032
rect 3973 20995 4031 21001
rect 3973 20961 3985 20995
rect 4019 20961 4031 20995
rect 3973 20955 4031 20961
rect 4249 20995 4307 21001
rect 4249 20961 4261 20995
rect 4295 20961 4307 20995
rect 4249 20955 4307 20961
rect 4433 20995 4491 21001
rect 4433 20961 4445 20995
rect 4479 20961 4491 20995
rect 4433 20955 4491 20961
rect 4525 20995 4583 21001
rect 4525 20961 4537 20995
rect 4571 20961 4583 20995
rect 4525 20955 4583 20961
rect 4154 20924 4160 20936
rect 1780 20896 4160 20924
rect 2056 20865 2084 20896
rect 4154 20884 4160 20896
rect 4212 20884 4218 20936
rect 2041 20859 2099 20865
rect 2041 20825 2053 20859
rect 2087 20825 2099 20859
rect 2041 20819 2099 20825
rect 3142 20816 3148 20868
rect 3200 20816 3206 20868
rect 4264 20856 4292 20955
rect 4448 20924 4476 20955
rect 4614 20952 4620 21004
rect 4672 20952 4678 21004
rect 4706 20952 4712 21004
rect 4764 20992 4770 21004
rect 4764 20964 4936 20992
rect 4764 20952 4770 20964
rect 4798 20924 4804 20936
rect 4448 20896 4804 20924
rect 4798 20884 4804 20896
rect 4856 20884 4862 20936
rect 4908 20924 4936 20964
rect 4982 20952 4988 21004
rect 5040 20952 5046 21004
rect 5258 20952 5264 21004
rect 5316 20952 5322 21004
rect 5445 20995 5503 21001
rect 5445 20961 5457 20995
rect 5491 20992 5503 20995
rect 5534 20992 5540 21004
rect 5491 20964 5540 20992
rect 5491 20961 5503 20964
rect 5445 20955 5503 20961
rect 5534 20952 5540 20964
rect 5592 20952 5598 21004
rect 5810 20952 5816 21004
rect 5868 20952 5874 21004
rect 6086 20952 6092 21004
rect 6144 20952 6150 21004
rect 6454 20952 6460 21004
rect 6512 20952 6518 21004
rect 6564 21001 6592 21032
rect 8456 21029 8468 21063
rect 8502 21060 8514 21063
rect 9125 21063 9183 21069
rect 9125 21060 9137 21063
rect 8502 21032 9137 21060
rect 8502 21029 8514 21032
rect 8456 21023 8514 21029
rect 9125 21029 9137 21032
rect 9171 21029 9183 21063
rect 9674 21060 9680 21072
rect 9125 21023 9183 21029
rect 9508 21032 9680 21060
rect 6549 20995 6607 21001
rect 6549 20961 6561 20995
rect 6595 20961 6607 20995
rect 6549 20955 6607 20961
rect 7098 20952 7104 21004
rect 7156 20992 7162 21004
rect 7193 20995 7251 21001
rect 7193 20992 7205 20995
rect 7156 20964 7205 20992
rect 7156 20952 7162 20964
rect 7193 20961 7205 20964
rect 7239 20961 7251 20995
rect 7193 20955 7251 20961
rect 7653 20995 7711 21001
rect 7653 20961 7665 20995
rect 7699 20992 7711 20995
rect 7834 20992 7840 21004
rect 7699 20964 7840 20992
rect 7699 20961 7711 20964
rect 7653 20955 7711 20961
rect 7834 20952 7840 20964
rect 7892 20952 7898 21004
rect 7926 20952 7932 21004
rect 7984 20952 7990 21004
rect 8110 20952 8116 21004
rect 8168 20992 8174 21004
rect 9033 20995 9091 21001
rect 9033 20992 9045 20995
rect 8168 20964 9045 20992
rect 8168 20952 8174 20964
rect 9033 20961 9045 20964
rect 9079 20961 9091 20995
rect 9033 20955 9091 20961
rect 6825 20927 6883 20933
rect 4908 20896 6040 20924
rect 4982 20856 4988 20868
rect 4264 20828 4988 20856
rect 4982 20816 4988 20828
rect 5040 20856 5046 20868
rect 5077 20859 5135 20865
rect 5077 20856 5089 20859
rect 5040 20828 5089 20856
rect 5040 20816 5046 20828
rect 5077 20825 5089 20828
rect 5123 20825 5135 20859
rect 6012 20856 6040 20896
rect 6825 20893 6837 20927
rect 6871 20893 6883 20927
rect 6825 20887 6883 20893
rect 6840 20856 6868 20887
rect 7006 20884 7012 20936
rect 7064 20924 7070 20936
rect 7282 20924 7288 20936
rect 7064 20896 7288 20924
rect 7064 20884 7070 20896
rect 7282 20884 7288 20896
rect 7340 20924 7346 20936
rect 7377 20927 7435 20933
rect 7377 20924 7389 20927
rect 7340 20896 7389 20924
rect 7340 20884 7346 20896
rect 7377 20893 7389 20896
rect 7423 20893 7435 20927
rect 7377 20887 7435 20893
rect 7469 20927 7527 20933
rect 7469 20893 7481 20927
rect 7515 20924 7527 20927
rect 8021 20927 8079 20933
rect 8021 20924 8033 20927
rect 7515 20896 8033 20924
rect 7515 20893 7527 20896
rect 7469 20887 7527 20893
rect 8021 20893 8033 20896
rect 8067 20893 8079 20927
rect 8021 20887 8079 20893
rect 8662 20884 8668 20936
rect 8720 20884 8726 20936
rect 8941 20927 8999 20933
rect 8941 20893 8953 20927
rect 8987 20924 8999 20927
rect 9508 20924 9536 21032
rect 9674 21020 9680 21032
rect 9732 21060 9738 21072
rect 9732 21032 9996 21060
rect 9732 21020 9738 21032
rect 9858 20952 9864 21004
rect 9916 20952 9922 21004
rect 8987 20896 9536 20924
rect 8987 20893 8999 20896
rect 8941 20887 8999 20893
rect 9582 20884 9588 20936
rect 9640 20924 9646 20936
rect 9677 20927 9735 20933
rect 9677 20924 9689 20927
rect 9640 20896 9689 20924
rect 9640 20884 9646 20896
rect 9677 20893 9689 20896
rect 9723 20893 9735 20927
rect 9677 20887 9735 20893
rect 9766 20884 9772 20936
rect 9824 20884 9830 20936
rect 9968 20933 9996 21032
rect 10778 21020 10784 21072
rect 10836 21060 10842 21072
rect 10836 21032 11192 21060
rect 10836 21020 10842 21032
rect 10042 20952 10048 21004
rect 10100 20992 10106 21004
rect 10686 20992 10692 21004
rect 10100 20964 10692 20992
rect 10100 20952 10106 20964
rect 10686 20952 10692 20964
rect 10744 20992 10750 21004
rect 11164 21001 11192 21032
rect 10965 20995 11023 21001
rect 10965 20992 10977 20995
rect 10744 20964 10977 20992
rect 10744 20952 10750 20964
rect 10965 20961 10977 20964
rect 11011 20961 11023 20995
rect 10965 20955 11023 20961
rect 11149 20995 11207 21001
rect 11149 20961 11161 20995
rect 11195 20961 11207 20995
rect 11149 20955 11207 20961
rect 11238 20952 11244 21004
rect 11296 20952 11302 21004
rect 11348 21001 11376 21100
rect 11698 21088 11704 21100
rect 11756 21088 11762 21140
rect 12158 21088 12164 21140
rect 12216 21128 12222 21140
rect 15197 21131 15255 21137
rect 12216 21100 14504 21128
rect 12216 21088 12222 21100
rect 11790 21020 11796 21072
rect 11848 21060 11854 21072
rect 14090 21060 14096 21072
rect 11848 21032 14096 21060
rect 11848 21020 11854 21032
rect 11333 20995 11391 21001
rect 11333 20961 11345 20995
rect 11379 20961 11391 20995
rect 11333 20955 11391 20961
rect 11974 20952 11980 21004
rect 12032 20952 12038 21004
rect 12066 20952 12072 21004
rect 12124 20952 12130 21004
rect 13262 20952 13268 21004
rect 13320 21001 13326 21004
rect 13556 21001 13584 21032
rect 14090 21020 14096 21032
rect 14148 21020 14154 21072
rect 14476 21060 14504 21100
rect 15197 21097 15209 21131
rect 15243 21128 15255 21131
rect 15378 21128 15384 21140
rect 15243 21100 15384 21128
rect 15243 21097 15255 21100
rect 15197 21091 15255 21097
rect 15378 21088 15384 21100
rect 15436 21088 15442 21140
rect 15746 21128 15752 21140
rect 15672 21100 15752 21128
rect 14734 21060 14740 21072
rect 14476 21032 14740 21060
rect 13320 20955 13332 21001
rect 13541 20995 13599 21001
rect 13541 20961 13553 20995
rect 13587 20961 13599 20995
rect 13541 20955 13599 20961
rect 13320 20952 13326 20955
rect 13814 20952 13820 21004
rect 13872 20952 13878 21004
rect 14476 21001 14504 21032
rect 14734 21020 14740 21032
rect 14792 21060 14798 21072
rect 15672 21069 15700 21100
rect 15746 21088 15752 21100
rect 15804 21088 15810 21140
rect 15933 21131 15991 21137
rect 15933 21097 15945 21131
rect 15979 21128 15991 21131
rect 19058 21128 19064 21140
rect 15979 21100 19064 21128
rect 15979 21097 15991 21100
rect 15933 21091 15991 21097
rect 19058 21088 19064 21100
rect 19116 21088 19122 21140
rect 19978 21088 19984 21140
rect 20036 21128 20042 21140
rect 20036 21100 20392 21128
rect 20036 21088 20042 21100
rect 15473 21063 15531 21069
rect 15473 21060 15485 21063
rect 14792 21032 15485 21060
rect 14792 21020 14798 21032
rect 15473 21029 15485 21032
rect 15519 21029 15531 21063
rect 15473 21023 15531 21029
rect 15657 21063 15715 21069
rect 15657 21029 15669 21063
rect 15703 21029 15715 21063
rect 17586 21060 17592 21072
rect 15657 21023 15715 21029
rect 15764 21032 17592 21060
rect 14461 20995 14519 21001
rect 14461 20961 14473 20995
rect 14507 20961 14519 20995
rect 14461 20955 14519 20961
rect 14826 20952 14832 21004
rect 14884 20952 14890 21004
rect 15764 21001 15792 21032
rect 17586 21020 17592 21032
rect 17644 21020 17650 21072
rect 18598 21020 18604 21072
rect 18656 21060 18662 21072
rect 20070 21060 20076 21072
rect 18656 21032 20076 21060
rect 18656 21020 18662 21032
rect 20070 21020 20076 21032
rect 20128 21020 20134 21072
rect 20364 21060 20392 21100
rect 20438 21088 20444 21140
rect 20496 21128 20502 21140
rect 20533 21131 20591 21137
rect 20533 21128 20545 21131
rect 20496 21100 20545 21128
rect 20496 21088 20502 21100
rect 20533 21097 20545 21100
rect 20579 21097 20591 21131
rect 21637 21131 21695 21137
rect 21637 21128 21649 21131
rect 20533 21091 20591 21097
rect 20640 21100 21649 21128
rect 20640 21060 20668 21100
rect 21637 21097 21649 21100
rect 21683 21097 21695 21131
rect 21637 21091 21695 21097
rect 20364 21032 20668 21060
rect 20806 21020 20812 21072
rect 20864 21020 20870 21072
rect 20898 21020 20904 21072
rect 20956 21020 20962 21072
rect 20990 21020 20996 21072
rect 21048 21060 21054 21072
rect 21453 21063 21511 21069
rect 21453 21060 21465 21063
rect 21048 21032 21465 21060
rect 21048 21020 21054 21032
rect 21453 21029 21465 21032
rect 21499 21029 21511 21063
rect 21453 21023 21511 21029
rect 16390 21001 16396 21004
rect 15749 20995 15807 21001
rect 15749 20961 15761 20995
rect 15795 20961 15807 20995
rect 15749 20955 15807 20961
rect 16384 20955 16396 21001
rect 16390 20952 16396 20955
rect 16448 20952 16454 21004
rect 16758 20952 16764 21004
rect 16816 20992 16822 21004
rect 18693 20995 18751 21001
rect 18693 20992 18705 20995
rect 16816 20964 18705 20992
rect 16816 20952 16822 20964
rect 18693 20961 18705 20964
rect 18739 20961 18751 20995
rect 18693 20955 18751 20961
rect 20714 20952 20720 21004
rect 20772 20952 20778 21004
rect 21082 20952 21088 21004
rect 21140 20952 21146 21004
rect 22738 20952 22744 21004
rect 22796 21001 22802 21004
rect 22796 20955 22808 21001
rect 22796 20952 22802 20955
rect 22922 20952 22928 21004
rect 22980 20992 22986 21004
rect 23017 20995 23075 21001
rect 23017 20992 23029 20995
rect 22980 20964 23029 20992
rect 22980 20952 22986 20964
rect 23017 20961 23029 20964
rect 23063 20961 23075 20995
rect 23017 20955 23075 20961
rect 9953 20927 10011 20933
rect 9953 20893 9965 20927
rect 9999 20924 10011 20927
rect 10318 20924 10324 20936
rect 9999 20896 10324 20924
rect 9999 20893 10011 20896
rect 9953 20887 10011 20893
rect 10318 20884 10324 20896
rect 10376 20884 10382 20936
rect 11054 20884 11060 20936
rect 11112 20924 11118 20936
rect 12084 20924 12112 20952
rect 11112 20896 12112 20924
rect 13909 20927 13967 20933
rect 11112 20884 11118 20896
rect 13909 20893 13921 20927
rect 13955 20893 13967 20927
rect 13909 20887 13967 20893
rect 6012 20828 6868 20856
rect 7561 20859 7619 20865
rect 5077 20819 5135 20825
rect 7561 20825 7573 20859
rect 7607 20856 7619 20859
rect 8297 20859 8355 20865
rect 8297 20856 8309 20859
rect 7607 20828 8309 20856
rect 7607 20825 7619 20828
rect 7561 20819 7619 20825
rect 8297 20825 8309 20828
rect 8343 20825 8355 20859
rect 8297 20819 8355 20825
rect 8386 20816 8392 20868
rect 8444 20856 8450 20868
rect 11609 20859 11667 20865
rect 8444 20828 9674 20856
rect 8444 20816 8450 20828
rect 2317 20791 2375 20797
rect 2317 20757 2329 20791
rect 2363 20788 2375 20791
rect 2593 20791 2651 20797
rect 2593 20788 2605 20791
rect 2363 20760 2605 20788
rect 2363 20757 2375 20760
rect 2317 20751 2375 20757
rect 2593 20757 2605 20760
rect 2639 20757 2651 20791
rect 2593 20751 2651 20757
rect 4062 20748 4068 20800
rect 4120 20748 4126 20800
rect 6089 20791 6147 20797
rect 6089 20757 6101 20791
rect 6135 20788 6147 20791
rect 6178 20788 6184 20800
rect 6135 20760 6184 20788
rect 6135 20757 6147 20760
rect 6089 20751 6147 20757
rect 6178 20748 6184 20760
rect 6236 20748 6242 20800
rect 6822 20748 6828 20800
rect 6880 20748 6886 20800
rect 7098 20748 7104 20800
rect 7156 20788 7162 20800
rect 7650 20788 7656 20800
rect 7156 20760 7656 20788
rect 7156 20748 7162 20760
rect 7650 20748 7656 20760
rect 7708 20748 7714 20800
rect 9490 20748 9496 20800
rect 9548 20748 9554 20800
rect 9646 20788 9674 20828
rect 11609 20825 11621 20859
rect 11655 20856 11667 20859
rect 12066 20856 12072 20868
rect 11655 20828 12072 20856
rect 11655 20825 11667 20828
rect 11609 20819 11667 20825
rect 12066 20816 12072 20828
rect 12124 20816 12130 20868
rect 13924 20856 13952 20887
rect 14182 20884 14188 20936
rect 14240 20924 14246 20936
rect 14737 20927 14795 20933
rect 14737 20924 14749 20927
rect 14240 20896 14749 20924
rect 14240 20884 14246 20896
rect 14737 20893 14749 20896
rect 14783 20893 14795 20927
rect 14737 20887 14795 20893
rect 15194 20884 15200 20936
rect 15252 20924 15258 20936
rect 16117 20927 16175 20933
rect 16117 20924 16129 20927
rect 15252 20896 16129 20924
rect 15252 20884 15258 20896
rect 16117 20893 16129 20896
rect 16163 20893 16175 20927
rect 16117 20887 16175 20893
rect 17586 20884 17592 20936
rect 17644 20884 17650 20936
rect 17862 20884 17868 20936
rect 17920 20884 17926 20936
rect 20441 20927 20499 20933
rect 20441 20924 20453 20927
rect 18708 20896 20453 20924
rect 18708 20868 18736 20896
rect 20441 20893 20453 20896
rect 20487 20924 20499 20927
rect 21266 20924 21272 20936
rect 20487 20896 21272 20924
rect 20487 20893 20499 20896
rect 20441 20887 20499 20893
rect 21266 20884 21272 20896
rect 21324 20924 21330 20936
rect 21634 20924 21640 20936
rect 21324 20896 21640 20924
rect 21324 20884 21330 20896
rect 21634 20884 21640 20896
rect 21692 20884 21698 20936
rect 14090 20856 14096 20868
rect 13924 20828 14096 20856
rect 14090 20816 14096 20828
rect 14148 20856 14154 20868
rect 14148 20828 15424 20856
rect 14148 20816 14154 20828
rect 11701 20791 11759 20797
rect 11701 20788 11713 20791
rect 9646 20760 11713 20788
rect 11701 20757 11713 20760
rect 11747 20757 11759 20791
rect 11701 20751 11759 20757
rect 11977 20791 12035 20797
rect 11977 20757 11989 20791
rect 12023 20788 12035 20791
rect 12158 20788 12164 20800
rect 12023 20760 12164 20788
rect 12023 20757 12035 20760
rect 11977 20751 12035 20757
rect 12158 20748 12164 20760
rect 12216 20748 12222 20800
rect 12526 20748 12532 20800
rect 12584 20788 12590 20800
rect 14277 20791 14335 20797
rect 14277 20788 14289 20791
rect 12584 20760 14289 20788
rect 12584 20748 12590 20760
rect 14277 20757 14289 20760
rect 14323 20788 14335 20791
rect 14366 20788 14372 20800
rect 14323 20760 14372 20788
rect 14323 20757 14335 20760
rect 14277 20751 14335 20757
rect 14366 20748 14372 20760
rect 14424 20748 14430 20800
rect 15286 20748 15292 20800
rect 15344 20748 15350 20800
rect 15396 20788 15424 20828
rect 17494 20816 17500 20868
rect 17552 20816 17558 20868
rect 18690 20816 18696 20868
rect 18748 20816 18754 20868
rect 20162 20816 20168 20868
rect 20220 20856 20226 20868
rect 21082 20856 21088 20868
rect 20220 20828 21088 20856
rect 20220 20816 20226 20828
rect 21082 20816 21088 20828
rect 21140 20816 21146 20868
rect 17512 20788 17540 20816
rect 15396 20760 17540 20788
rect 20346 20748 20352 20800
rect 20404 20788 20410 20800
rect 21361 20791 21419 20797
rect 21361 20788 21373 20791
rect 20404 20760 21373 20788
rect 20404 20748 20410 20760
rect 21361 20757 21373 20760
rect 21407 20757 21419 20791
rect 21361 20751 21419 20757
rect 22094 20748 22100 20800
rect 22152 20788 22158 20800
rect 22370 20788 22376 20800
rect 22152 20760 22376 20788
rect 22152 20748 22158 20760
rect 22370 20748 22376 20760
rect 22428 20748 22434 20800
rect 552 20698 23368 20720
rect 552 20646 1366 20698
rect 1418 20646 1430 20698
rect 1482 20646 1494 20698
rect 1546 20646 1558 20698
rect 1610 20646 1622 20698
rect 1674 20646 1686 20698
rect 1738 20646 7366 20698
rect 7418 20646 7430 20698
rect 7482 20646 7494 20698
rect 7546 20646 7558 20698
rect 7610 20646 7622 20698
rect 7674 20646 7686 20698
rect 7738 20646 13366 20698
rect 13418 20646 13430 20698
rect 13482 20646 13494 20698
rect 13546 20646 13558 20698
rect 13610 20646 13622 20698
rect 13674 20646 13686 20698
rect 13738 20646 19366 20698
rect 19418 20646 19430 20698
rect 19482 20646 19494 20698
rect 19546 20646 19558 20698
rect 19610 20646 19622 20698
rect 19674 20646 19686 20698
rect 19738 20646 23368 20698
rect 552 20624 23368 20646
rect 1854 20544 1860 20596
rect 1912 20584 1918 20596
rect 2682 20584 2688 20596
rect 1912 20556 2688 20584
rect 1912 20544 1918 20556
rect 2682 20544 2688 20556
rect 2740 20544 2746 20596
rect 6362 20544 6368 20596
rect 6420 20544 6426 20596
rect 6638 20544 6644 20596
rect 6696 20584 6702 20596
rect 6825 20587 6883 20593
rect 6825 20584 6837 20587
rect 6696 20556 6837 20584
rect 6696 20544 6702 20556
rect 6825 20553 6837 20556
rect 6871 20553 6883 20587
rect 6825 20547 6883 20553
rect 7190 20544 7196 20596
rect 7248 20544 7254 20596
rect 7926 20544 7932 20596
rect 7984 20544 7990 20596
rect 8570 20544 8576 20596
rect 8628 20584 8634 20596
rect 9766 20584 9772 20596
rect 8628 20556 9772 20584
rect 8628 20544 8634 20556
rect 9766 20544 9772 20556
rect 9824 20544 9830 20596
rect 10226 20544 10232 20596
rect 10284 20584 10290 20596
rect 10597 20587 10655 20593
rect 10597 20584 10609 20587
rect 10284 20556 10609 20584
rect 10284 20544 10290 20556
rect 10597 20553 10609 20556
rect 10643 20553 10655 20587
rect 10597 20547 10655 20553
rect 10686 20544 10692 20596
rect 10744 20584 10750 20596
rect 10781 20587 10839 20593
rect 10781 20584 10793 20587
rect 10744 20556 10793 20584
rect 10744 20544 10750 20556
rect 10781 20553 10793 20556
rect 10827 20553 10839 20587
rect 10781 20547 10839 20553
rect 11422 20544 11428 20596
rect 11480 20544 11486 20596
rect 12802 20544 12808 20596
rect 12860 20584 12866 20596
rect 13173 20587 13231 20593
rect 13173 20584 13185 20587
rect 12860 20556 13185 20584
rect 12860 20544 12866 20556
rect 13173 20553 13185 20556
rect 13219 20553 13231 20587
rect 13173 20547 13231 20553
rect 5534 20476 5540 20528
rect 5592 20516 5598 20528
rect 6656 20516 6684 20544
rect 5592 20488 6684 20516
rect 5592 20476 5598 20488
rect 6914 20476 6920 20528
rect 6972 20516 6978 20528
rect 7561 20519 7619 20525
rect 7561 20516 7573 20519
rect 6972 20488 7573 20516
rect 6972 20476 6978 20488
rect 7561 20485 7573 20488
rect 7607 20485 7619 20519
rect 7561 20479 7619 20485
rect 8941 20519 8999 20525
rect 8941 20485 8953 20519
rect 8987 20516 8999 20519
rect 11514 20516 11520 20528
rect 8987 20488 10180 20516
rect 8987 20485 8999 20488
rect 8941 20479 8999 20485
rect 3234 20408 3240 20460
rect 3292 20408 3298 20460
rect 4614 20408 4620 20460
rect 4672 20448 4678 20460
rect 4890 20448 4896 20460
rect 4672 20420 4896 20448
rect 4672 20408 4678 20420
rect 4890 20408 4896 20420
rect 4948 20408 4954 20460
rect 7653 20451 7711 20457
rect 7653 20417 7665 20451
rect 7699 20448 7711 20451
rect 9401 20451 9459 20457
rect 7699 20420 7880 20448
rect 7699 20417 7711 20420
rect 7653 20411 7711 20417
rect 1581 20383 1639 20389
rect 1581 20349 1593 20383
rect 1627 20380 1639 20383
rect 1854 20380 1860 20392
rect 1627 20352 1860 20380
rect 1627 20349 1639 20352
rect 1581 20343 1639 20349
rect 1854 20340 1860 20352
rect 1912 20340 1918 20392
rect 2038 20340 2044 20392
rect 2096 20340 2102 20392
rect 2498 20340 2504 20392
rect 2556 20340 2562 20392
rect 2685 20383 2743 20389
rect 2685 20349 2697 20383
rect 2731 20380 2743 20383
rect 2774 20380 2780 20392
rect 2731 20352 2780 20380
rect 2731 20349 2743 20352
rect 2685 20343 2743 20349
rect 2774 20340 2780 20352
rect 2832 20380 2838 20392
rect 4062 20380 4068 20392
rect 2832 20352 4068 20380
rect 2832 20340 2838 20352
rect 4062 20340 4068 20352
rect 4120 20340 4126 20392
rect 6914 20340 6920 20392
rect 6972 20340 6978 20392
rect 7374 20340 7380 20392
rect 7432 20340 7438 20392
rect 1765 20315 1823 20321
rect 1765 20281 1777 20315
rect 1811 20312 1823 20315
rect 2056 20312 2084 20340
rect 1811 20284 2084 20312
rect 1811 20281 1823 20284
rect 1765 20275 1823 20281
rect 2590 20272 2596 20324
rect 2648 20312 2654 20324
rect 3482 20315 3540 20321
rect 3482 20312 3494 20315
rect 2648 20284 3494 20312
rect 2648 20272 2654 20284
rect 3482 20281 3494 20284
rect 3528 20281 3540 20315
rect 3482 20275 3540 20281
rect 4893 20315 4951 20321
rect 4893 20281 4905 20315
rect 4939 20312 4951 20315
rect 5534 20312 5540 20324
rect 4939 20284 5540 20312
rect 4939 20281 4951 20284
rect 4893 20275 4951 20281
rect 5534 20272 5540 20284
rect 5592 20272 5598 20324
rect 6178 20272 6184 20324
rect 6236 20312 6242 20324
rect 6236 20284 7788 20312
rect 6236 20272 6242 20284
rect 1394 20204 1400 20256
rect 1452 20204 1458 20256
rect 1949 20247 2007 20253
rect 1949 20213 1961 20247
rect 1995 20244 2007 20247
rect 2038 20244 2044 20256
rect 1995 20216 2044 20244
rect 1995 20213 2007 20216
rect 1949 20207 2007 20213
rect 2038 20204 2044 20216
rect 2096 20204 2102 20256
rect 2682 20204 2688 20256
rect 2740 20204 2746 20256
rect 4338 20204 4344 20256
rect 4396 20244 4402 20256
rect 4617 20247 4675 20253
rect 4617 20244 4629 20247
rect 4396 20216 4629 20244
rect 4396 20204 4402 20216
rect 4617 20213 4629 20216
rect 4663 20244 4675 20247
rect 5350 20244 5356 20256
rect 4663 20216 5356 20244
rect 4663 20213 4675 20216
rect 4617 20207 4675 20213
rect 5350 20204 5356 20216
rect 5408 20204 5414 20256
rect 7006 20204 7012 20256
rect 7064 20244 7070 20256
rect 7650 20244 7656 20256
rect 7064 20216 7656 20244
rect 7064 20204 7070 20216
rect 7650 20204 7656 20216
rect 7708 20204 7714 20256
rect 7760 20253 7788 20284
rect 7745 20247 7803 20253
rect 7745 20213 7757 20247
rect 7791 20213 7803 20247
rect 7852 20244 7880 20420
rect 9401 20417 9413 20451
rect 9447 20448 9459 20451
rect 9447 20420 10088 20448
rect 9447 20417 9459 20420
rect 9401 20411 9459 20417
rect 7929 20383 7987 20389
rect 7929 20349 7941 20383
rect 7975 20349 7987 20383
rect 7929 20343 7987 20349
rect 7951 20312 7979 20343
rect 8018 20340 8024 20392
rect 8076 20340 8082 20392
rect 8205 20383 8263 20389
rect 8205 20349 8217 20383
rect 8251 20380 8263 20383
rect 8386 20380 8392 20392
rect 8251 20352 8392 20380
rect 8251 20349 8263 20352
rect 8205 20343 8263 20349
rect 8110 20312 8116 20324
rect 7951 20284 8116 20312
rect 8110 20272 8116 20284
rect 8168 20272 8174 20324
rect 8220 20244 8248 20343
rect 8386 20340 8392 20352
rect 8444 20340 8450 20392
rect 8570 20340 8576 20392
rect 8628 20340 8634 20392
rect 8754 20340 8760 20392
rect 8812 20340 8818 20392
rect 9490 20340 9496 20392
rect 9548 20380 9554 20392
rect 9585 20383 9643 20389
rect 9585 20380 9597 20383
rect 9548 20352 9597 20380
rect 9548 20340 9554 20352
rect 9585 20349 9597 20352
rect 9631 20349 9643 20383
rect 9585 20343 9643 20349
rect 9677 20383 9735 20389
rect 9677 20349 9689 20383
rect 9723 20380 9735 20383
rect 9858 20380 9864 20392
rect 9723 20352 9864 20380
rect 9723 20349 9735 20352
rect 9677 20343 9735 20349
rect 9858 20340 9864 20352
rect 9916 20340 9922 20392
rect 9950 20340 9956 20392
rect 10008 20340 10014 20392
rect 10060 20389 10088 20420
rect 10060 20383 10123 20389
rect 10060 20352 10077 20383
rect 10065 20349 10077 20352
rect 10111 20349 10123 20383
rect 10152 20380 10180 20488
rect 10980 20488 11520 20516
rect 10229 20383 10287 20389
rect 10229 20380 10241 20383
rect 10152 20352 10241 20380
rect 10065 20343 10123 20349
rect 10229 20349 10241 20352
rect 10275 20349 10287 20383
rect 10229 20343 10287 20349
rect 10318 20340 10324 20392
rect 10376 20340 10382 20392
rect 10410 20340 10416 20392
rect 10468 20340 10474 20392
rect 10980 20389 11008 20488
rect 11514 20476 11520 20488
rect 11572 20476 11578 20528
rect 11790 20408 11796 20460
rect 11848 20408 11854 20460
rect 13188 20448 13216 20547
rect 13262 20544 13268 20596
rect 13320 20584 13326 20596
rect 13541 20587 13599 20593
rect 13541 20584 13553 20587
rect 13320 20556 13553 20584
rect 13320 20544 13326 20556
rect 13541 20553 13553 20556
rect 13587 20553 13599 20587
rect 13541 20547 13599 20553
rect 14277 20587 14335 20593
rect 14277 20553 14289 20587
rect 14323 20584 14335 20587
rect 14458 20584 14464 20596
rect 14323 20556 14464 20584
rect 14323 20553 14335 20556
rect 14277 20547 14335 20553
rect 14458 20544 14464 20556
rect 14516 20544 14522 20596
rect 14550 20544 14556 20596
rect 14608 20544 14614 20596
rect 14737 20587 14795 20593
rect 14737 20553 14749 20587
rect 14783 20584 14795 20587
rect 14826 20584 14832 20596
rect 14783 20556 14832 20584
rect 14783 20553 14795 20556
rect 14737 20547 14795 20553
rect 14826 20544 14832 20556
rect 14884 20544 14890 20596
rect 15654 20544 15660 20596
rect 15712 20584 15718 20596
rect 15749 20587 15807 20593
rect 15749 20584 15761 20587
rect 15712 20556 15761 20584
rect 15712 20544 15718 20556
rect 15749 20553 15761 20556
rect 15795 20553 15807 20587
rect 15749 20547 15807 20553
rect 16390 20544 16396 20596
rect 16448 20584 16454 20596
rect 16577 20587 16635 20593
rect 16577 20584 16589 20587
rect 16448 20556 16589 20584
rect 16448 20544 16454 20556
rect 16577 20553 16589 20556
rect 16623 20553 16635 20587
rect 17310 20584 17316 20596
rect 16577 20547 16635 20553
rect 16776 20556 17316 20584
rect 16776 20516 16804 20556
rect 17310 20544 17316 20556
rect 17368 20584 17374 20596
rect 17862 20584 17868 20596
rect 17368 20556 17868 20584
rect 17368 20544 17374 20556
rect 17862 20544 17868 20556
rect 17920 20544 17926 20596
rect 18138 20544 18144 20596
rect 18196 20584 18202 20596
rect 20165 20587 20223 20593
rect 20165 20584 20177 20587
rect 18196 20556 20177 20584
rect 18196 20544 18202 20556
rect 20165 20553 20177 20556
rect 20211 20553 20223 20587
rect 20165 20547 20223 20553
rect 21729 20587 21787 20593
rect 21729 20553 21741 20587
rect 21775 20584 21787 20587
rect 22278 20584 22284 20596
rect 21775 20556 22284 20584
rect 21775 20553 21787 20556
rect 21729 20547 21787 20553
rect 22278 20544 22284 20556
rect 22336 20544 22342 20596
rect 22649 20587 22707 20593
rect 22649 20553 22661 20587
rect 22695 20553 22707 20587
rect 22649 20547 22707 20553
rect 14384 20488 16344 20516
rect 13814 20448 13820 20460
rect 13188 20420 13820 20448
rect 13814 20408 13820 20420
rect 13872 20448 13878 20460
rect 13909 20451 13967 20457
rect 13909 20448 13921 20451
rect 13872 20420 13921 20448
rect 13872 20408 13878 20420
rect 13909 20417 13921 20420
rect 13955 20417 13967 20451
rect 13909 20411 13967 20417
rect 10965 20383 11023 20389
rect 10965 20349 10977 20383
rect 11011 20349 11023 20383
rect 10965 20343 11023 20349
rect 11057 20383 11115 20389
rect 11057 20349 11069 20383
rect 11103 20380 11115 20383
rect 11238 20380 11244 20392
rect 11103 20352 11244 20380
rect 11103 20349 11115 20352
rect 11057 20343 11115 20349
rect 11238 20340 11244 20352
rect 11296 20380 11302 20392
rect 11514 20380 11520 20392
rect 11296 20352 11520 20380
rect 11296 20340 11302 20352
rect 11514 20340 11520 20352
rect 11572 20340 11578 20392
rect 13725 20383 13783 20389
rect 13725 20349 13737 20383
rect 13771 20349 13783 20383
rect 13725 20343 13783 20349
rect 12066 20321 12072 20324
rect 9125 20315 9183 20321
rect 9125 20312 9137 20315
rect 8588 20284 9137 20312
rect 7852 20216 8248 20244
rect 7745 20207 7803 20213
rect 8478 20204 8484 20256
rect 8536 20244 8542 20256
rect 8588 20253 8616 20284
rect 9125 20281 9137 20284
rect 9171 20281 9183 20315
rect 9125 20275 9183 20281
rect 9309 20315 9367 20321
rect 9309 20281 9321 20315
rect 9355 20312 9367 20315
rect 12060 20312 12072 20321
rect 9355 20284 10824 20312
rect 12027 20284 12072 20312
rect 9355 20281 9367 20284
rect 9309 20275 9367 20281
rect 8573 20247 8631 20253
rect 8573 20244 8585 20247
rect 8536 20216 8585 20244
rect 8536 20204 8542 20216
rect 8573 20213 8585 20216
rect 8619 20213 8631 20247
rect 8573 20207 8631 20213
rect 9766 20204 9772 20256
rect 9824 20204 9830 20256
rect 10796 20244 10824 20284
rect 12060 20275 12072 20284
rect 12066 20272 12072 20275
rect 12124 20272 12130 20324
rect 13740 20312 13768 20343
rect 14090 20340 14096 20392
rect 14148 20340 14154 20392
rect 14384 20389 14412 20488
rect 14918 20408 14924 20460
rect 14976 20448 14982 20460
rect 15105 20451 15163 20457
rect 15105 20448 15117 20451
rect 14976 20420 15117 20448
rect 14976 20408 14982 20420
rect 15105 20417 15117 20420
rect 15151 20417 15163 20451
rect 15105 20411 15163 20417
rect 16206 20408 16212 20460
rect 16264 20408 16270 20460
rect 14369 20383 14427 20389
rect 14369 20349 14381 20383
rect 14415 20349 14427 20383
rect 14369 20343 14427 20349
rect 14645 20383 14703 20389
rect 14645 20349 14657 20383
rect 14691 20349 14703 20383
rect 14645 20343 14703 20349
rect 12406 20284 13768 20312
rect 11054 20244 11060 20256
rect 10796 20216 11060 20244
rect 11054 20204 11060 20216
rect 11112 20204 11118 20256
rect 11422 20204 11428 20256
rect 11480 20204 11486 20256
rect 11609 20247 11667 20253
rect 11609 20213 11621 20247
rect 11655 20244 11667 20247
rect 12406 20244 12434 20284
rect 14274 20272 14280 20324
rect 14332 20312 14338 20324
rect 14660 20312 14688 20343
rect 14734 20340 14740 20392
rect 14792 20380 14798 20392
rect 14829 20383 14887 20389
rect 14829 20380 14841 20383
rect 14792 20352 14841 20380
rect 14792 20340 14798 20352
rect 14829 20349 14841 20352
rect 14875 20349 14887 20383
rect 14829 20343 14887 20349
rect 15286 20340 15292 20392
rect 15344 20340 15350 20392
rect 15473 20383 15531 20389
rect 15473 20349 15485 20383
rect 15519 20380 15531 20383
rect 15654 20380 15660 20392
rect 15519 20352 15660 20380
rect 15519 20349 15531 20352
rect 15473 20343 15531 20349
rect 15654 20340 15660 20352
rect 15712 20340 15718 20392
rect 15746 20340 15752 20392
rect 15804 20380 15810 20392
rect 16117 20383 16175 20389
rect 16117 20380 16129 20383
rect 15804 20352 16129 20380
rect 15804 20340 15810 20352
rect 16117 20349 16129 20352
rect 16163 20349 16175 20383
rect 16117 20343 16175 20349
rect 15764 20312 15792 20340
rect 14332 20284 15792 20312
rect 16316 20312 16344 20488
rect 16408 20488 16804 20516
rect 16408 20457 16436 20488
rect 16850 20476 16856 20528
rect 16908 20476 16914 20528
rect 17129 20519 17187 20525
rect 17129 20485 17141 20519
rect 17175 20516 17187 20519
rect 17218 20516 17224 20528
rect 17175 20488 17224 20516
rect 17175 20485 17187 20488
rect 17129 20479 17187 20485
rect 17218 20476 17224 20488
rect 17276 20476 17282 20528
rect 20714 20516 20720 20528
rect 19352 20488 20720 20516
rect 16393 20451 16451 20457
rect 16393 20417 16405 20451
rect 16439 20417 16451 20451
rect 16868 20448 16896 20476
rect 16393 20411 16451 20417
rect 16776 20420 16896 20448
rect 16776 20389 16804 20420
rect 16942 20408 16948 20460
rect 17000 20408 17006 20460
rect 19352 20457 19380 20488
rect 20714 20476 20720 20488
rect 20772 20476 20778 20528
rect 20806 20476 20812 20528
rect 20864 20476 20870 20528
rect 21453 20519 21511 20525
rect 21453 20485 21465 20519
rect 21499 20516 21511 20519
rect 21818 20516 21824 20528
rect 21499 20488 21824 20516
rect 21499 20485 21511 20488
rect 21453 20479 21511 20485
rect 21818 20476 21824 20488
rect 21876 20476 21882 20528
rect 22094 20476 22100 20528
rect 22152 20516 22158 20528
rect 22664 20516 22692 20547
rect 22152 20488 22692 20516
rect 22152 20476 22158 20488
rect 19337 20451 19395 20457
rect 19337 20448 19349 20451
rect 18432 20420 19349 20448
rect 16761 20383 16819 20389
rect 16761 20349 16773 20383
rect 16807 20349 16819 20383
rect 16761 20343 16819 20349
rect 16850 20340 16856 20392
rect 16908 20340 16914 20392
rect 18432 20380 18460 20420
rect 19337 20417 19349 20420
rect 19383 20417 19395 20451
rect 21174 20448 21180 20460
rect 19337 20411 19395 20417
rect 19628 20420 21180 20448
rect 17144 20352 18460 20380
rect 17034 20312 17040 20324
rect 16316 20284 17040 20312
rect 14332 20272 14338 20284
rect 17034 20272 17040 20284
rect 17092 20272 17098 20324
rect 11655 20216 12434 20244
rect 11655 20213 11667 20216
rect 11609 20207 11667 20213
rect 12618 20204 12624 20256
rect 12676 20244 12682 20256
rect 15286 20244 15292 20256
rect 12676 20216 15292 20244
rect 12676 20204 12682 20216
rect 15286 20204 15292 20216
rect 15344 20204 15350 20256
rect 15562 20204 15568 20256
rect 15620 20244 15626 20256
rect 17144 20244 17172 20352
rect 18506 20340 18512 20392
rect 18564 20340 18570 20392
rect 19628 20380 19656 20420
rect 21174 20408 21180 20420
rect 21232 20408 21238 20460
rect 22554 20448 22560 20460
rect 22204 20420 22560 20448
rect 18616 20352 19656 20380
rect 20349 20383 20407 20389
rect 18264 20315 18322 20321
rect 18264 20281 18276 20315
rect 18310 20312 18322 20315
rect 18616 20312 18644 20352
rect 20349 20349 20361 20383
rect 20395 20349 20407 20383
rect 20349 20343 20407 20349
rect 20717 20383 20775 20389
rect 20717 20349 20729 20383
rect 20763 20380 20775 20383
rect 20898 20380 20904 20392
rect 20763 20352 20904 20380
rect 20763 20349 20775 20352
rect 20717 20343 20775 20349
rect 18310 20284 18644 20312
rect 18310 20281 18322 20284
rect 18264 20275 18322 20281
rect 18690 20272 18696 20324
rect 18748 20272 18754 20324
rect 18874 20272 18880 20324
rect 18932 20272 18938 20324
rect 15620 20216 17172 20244
rect 15620 20204 15626 20216
rect 17954 20204 17960 20256
rect 18012 20244 18018 20256
rect 19061 20247 19119 20253
rect 19061 20244 19073 20247
rect 18012 20216 19073 20244
rect 18012 20204 18018 20216
rect 19061 20213 19073 20216
rect 19107 20213 19119 20247
rect 19061 20207 19119 20213
rect 19334 20204 19340 20256
rect 19392 20244 19398 20256
rect 19429 20247 19487 20253
rect 19429 20244 19441 20247
rect 19392 20216 19441 20244
rect 19392 20204 19398 20216
rect 19429 20213 19441 20216
rect 19475 20213 19487 20247
rect 19429 20207 19487 20213
rect 19518 20204 19524 20256
rect 19576 20204 19582 20256
rect 19886 20204 19892 20256
rect 19944 20204 19950 20256
rect 20364 20244 20392 20343
rect 20898 20340 20904 20352
rect 20956 20340 20962 20392
rect 20990 20340 20996 20392
rect 21048 20340 21054 20392
rect 21085 20383 21143 20389
rect 21085 20349 21097 20383
rect 21131 20380 21143 20383
rect 21266 20380 21272 20392
rect 21131 20352 21272 20380
rect 21131 20349 21143 20352
rect 21085 20343 21143 20349
rect 21266 20340 21272 20352
rect 21324 20340 21330 20392
rect 21358 20340 21364 20392
rect 21416 20340 21422 20392
rect 21542 20340 21548 20392
rect 21600 20380 21606 20392
rect 21729 20383 21787 20389
rect 21729 20380 21741 20383
rect 21600 20352 21741 20380
rect 21600 20340 21606 20352
rect 21729 20349 21741 20352
rect 21775 20349 21787 20383
rect 21729 20343 21787 20349
rect 21818 20340 21824 20392
rect 21876 20380 21882 20392
rect 22204 20389 22232 20420
rect 22554 20408 22560 20420
rect 22612 20408 22618 20460
rect 21913 20383 21971 20389
rect 21913 20380 21925 20383
rect 21876 20352 21925 20380
rect 21876 20340 21882 20352
rect 21913 20349 21925 20352
rect 21959 20349 21971 20383
rect 21913 20343 21971 20349
rect 22189 20383 22247 20389
rect 22189 20349 22201 20383
rect 22235 20349 22247 20383
rect 22189 20343 22247 20349
rect 20438 20272 20444 20324
rect 20496 20272 20502 20324
rect 20530 20272 20536 20324
rect 20588 20312 20594 20324
rect 21177 20315 21235 20321
rect 21177 20312 21189 20315
rect 20588 20284 21189 20312
rect 20588 20272 20594 20284
rect 21177 20281 21189 20284
rect 21223 20312 21235 20315
rect 21450 20312 21456 20324
rect 21223 20284 21456 20312
rect 21223 20281 21235 20284
rect 21177 20275 21235 20281
rect 21450 20272 21456 20284
rect 21508 20272 21514 20324
rect 21928 20312 21956 20343
rect 22370 20340 22376 20392
rect 22428 20380 22434 20392
rect 23474 20380 23480 20392
rect 22428 20352 23480 20380
rect 22428 20340 22434 20352
rect 23474 20340 23480 20352
rect 23532 20340 23538 20392
rect 22465 20315 22523 20321
rect 22465 20312 22477 20315
rect 21928 20284 22477 20312
rect 22465 20281 22477 20284
rect 22511 20281 22523 20315
rect 22465 20275 22523 20281
rect 22554 20272 22560 20324
rect 22612 20312 22618 20324
rect 22681 20315 22739 20321
rect 22681 20312 22693 20315
rect 22612 20284 22693 20312
rect 22612 20272 22618 20284
rect 22681 20281 22693 20284
rect 22727 20312 22739 20315
rect 23290 20312 23296 20324
rect 22727 20284 23296 20312
rect 22727 20281 22739 20284
rect 22681 20275 22739 20281
rect 23290 20272 23296 20284
rect 23348 20272 23354 20324
rect 20714 20244 20720 20256
rect 20364 20216 20720 20244
rect 20714 20204 20720 20216
rect 20772 20204 20778 20256
rect 21910 20204 21916 20256
rect 21968 20244 21974 20256
rect 22005 20247 22063 20253
rect 22005 20244 22017 20247
rect 21968 20216 22017 20244
rect 21968 20204 21974 20216
rect 22005 20213 22017 20216
rect 22051 20213 22063 20247
rect 22005 20207 22063 20213
rect 22833 20247 22891 20253
rect 22833 20213 22845 20247
rect 22879 20244 22891 20247
rect 23014 20244 23020 20256
rect 22879 20216 23020 20244
rect 22879 20213 22891 20216
rect 22833 20207 22891 20213
rect 23014 20204 23020 20216
rect 23072 20204 23078 20256
rect 552 20154 23368 20176
rect 552 20102 4366 20154
rect 4418 20102 4430 20154
rect 4482 20102 4494 20154
rect 4546 20102 4558 20154
rect 4610 20102 4622 20154
rect 4674 20102 4686 20154
rect 4738 20102 10366 20154
rect 10418 20102 10430 20154
rect 10482 20102 10494 20154
rect 10546 20102 10558 20154
rect 10610 20102 10622 20154
rect 10674 20102 10686 20154
rect 10738 20102 16366 20154
rect 16418 20102 16430 20154
rect 16482 20102 16494 20154
rect 16546 20102 16558 20154
rect 16610 20102 16622 20154
rect 16674 20102 16686 20154
rect 16738 20102 22366 20154
rect 22418 20102 22430 20154
rect 22482 20102 22494 20154
rect 22546 20102 22558 20154
rect 22610 20102 22622 20154
rect 22674 20102 22686 20154
rect 22738 20102 23368 20154
rect 552 20080 23368 20102
rect 1765 20043 1823 20049
rect 1765 20009 1777 20043
rect 1811 20040 1823 20043
rect 1946 20040 1952 20052
rect 1811 20012 1952 20040
rect 1811 20009 1823 20012
rect 1765 20003 1823 20009
rect 1946 20000 1952 20012
rect 2004 20000 2010 20052
rect 2682 20000 2688 20052
rect 2740 20040 2746 20052
rect 2793 20043 2851 20049
rect 2793 20040 2805 20043
rect 2740 20012 2805 20040
rect 2740 20000 2746 20012
rect 2793 20009 2805 20012
rect 2839 20009 2851 20043
rect 2793 20003 2851 20009
rect 4617 20043 4675 20049
rect 4617 20009 4629 20043
rect 4663 20040 4675 20043
rect 4798 20040 4804 20052
rect 4663 20012 4804 20040
rect 4663 20009 4675 20012
rect 4617 20003 4675 20009
rect 4798 20000 4804 20012
rect 4856 20000 4862 20052
rect 5077 20043 5135 20049
rect 5077 20009 5089 20043
rect 5123 20040 5135 20043
rect 5258 20040 5264 20052
rect 5123 20012 5264 20040
rect 5123 20009 5135 20012
rect 5077 20003 5135 20009
rect 5258 20000 5264 20012
rect 5316 20000 5322 20052
rect 5810 20000 5816 20052
rect 5868 20000 5874 20052
rect 6178 20000 6184 20052
rect 6236 20000 6242 20052
rect 6273 20043 6331 20049
rect 6273 20009 6285 20043
rect 6319 20040 6331 20043
rect 6641 20043 6699 20049
rect 6641 20040 6653 20043
rect 6319 20012 6653 20040
rect 6319 20009 6331 20012
rect 6273 20003 6331 20009
rect 6641 20009 6653 20012
rect 6687 20009 6699 20043
rect 6641 20003 6699 20009
rect 7926 20000 7932 20052
rect 7984 20000 7990 20052
rect 9766 20040 9772 20052
rect 8772 20012 9772 20040
rect 1121 19975 1179 19981
rect 1121 19941 1133 19975
rect 1167 19972 1179 19975
rect 1167 19944 2084 19972
rect 1167 19941 1179 19944
rect 1121 19935 1179 19941
rect 2056 19916 2084 19944
rect 2498 19932 2504 19984
rect 2556 19932 2562 19984
rect 2593 19975 2651 19981
rect 2593 19941 2605 19975
rect 2639 19972 2651 19975
rect 2958 19972 2964 19984
rect 2639 19944 2964 19972
rect 2639 19941 2651 19944
rect 2593 19935 2651 19941
rect 2958 19932 2964 19944
rect 3016 19932 3022 19984
rect 4246 19932 4252 19984
rect 4304 19972 4310 19984
rect 5169 19975 5227 19981
rect 5169 19972 5181 19975
rect 4304 19944 5181 19972
rect 4304 19932 4310 19944
rect 5169 19941 5181 19944
rect 5215 19941 5227 19975
rect 5169 19935 5227 19941
rect 5350 19932 5356 19984
rect 5408 19972 5414 19984
rect 7944 19972 7972 20000
rect 5408 19944 7972 19972
rect 5408 19932 5414 19944
rect 1394 19864 1400 19916
rect 1452 19904 1458 19916
rect 1581 19907 1639 19913
rect 1581 19904 1593 19907
rect 1452 19876 1593 19904
rect 1452 19864 1458 19876
rect 1581 19873 1593 19876
rect 1627 19904 1639 19907
rect 1857 19907 1915 19913
rect 1857 19904 1869 19907
rect 1627 19876 1869 19904
rect 1627 19873 1639 19876
rect 1581 19867 1639 19873
rect 1857 19873 1869 19876
rect 1903 19873 1915 19907
rect 1857 19867 1915 19873
rect 2038 19864 2044 19916
rect 2096 19864 2102 19916
rect 2317 19907 2375 19913
rect 2317 19873 2329 19907
rect 2363 19904 2375 19907
rect 2774 19904 2780 19916
rect 2363 19876 2780 19904
rect 2363 19873 2375 19876
rect 2317 19867 2375 19873
rect 2774 19864 2780 19876
rect 2832 19864 2838 19916
rect 3145 19907 3203 19913
rect 3145 19873 3157 19907
rect 3191 19904 3203 19907
rect 3234 19904 3240 19916
rect 3191 19876 3240 19904
rect 3191 19873 3203 19876
rect 3145 19867 3203 19873
rect 3234 19864 3240 19876
rect 3292 19864 3298 19916
rect 3418 19913 3424 19916
rect 3412 19867 3424 19913
rect 3418 19864 3424 19867
rect 3476 19864 3482 19916
rect 4801 19907 4859 19913
rect 4801 19873 4813 19907
rect 4847 19904 4859 19907
rect 5074 19904 5080 19916
rect 4847 19876 5080 19904
rect 4847 19873 4859 19876
rect 4801 19867 4859 19873
rect 5074 19864 5080 19876
rect 5132 19864 5138 19916
rect 5442 19864 5448 19916
rect 5500 19864 5506 19916
rect 5644 19913 5672 19944
rect 5629 19907 5687 19913
rect 5629 19873 5641 19907
rect 5675 19873 5687 19907
rect 5629 19867 5687 19873
rect 6178 19864 6184 19916
rect 6236 19904 6242 19916
rect 6825 19907 6883 19913
rect 6825 19904 6837 19907
rect 6236 19876 6837 19904
rect 6236 19864 6242 19876
rect 6825 19873 6837 19876
rect 6871 19873 6883 19907
rect 6825 19867 6883 19873
rect 7101 19907 7159 19913
rect 7101 19873 7113 19907
rect 7147 19873 7159 19907
rect 7101 19867 7159 19873
rect 1489 19839 1547 19845
rect 1489 19805 1501 19839
rect 1535 19836 1547 19839
rect 1762 19836 1768 19848
rect 1535 19808 1768 19836
rect 1535 19805 1547 19808
rect 1489 19799 1547 19805
rect 1762 19796 1768 19808
rect 1820 19796 1826 19848
rect 4893 19839 4951 19845
rect 4893 19805 4905 19839
rect 4939 19836 4951 19839
rect 4982 19836 4988 19848
rect 4939 19808 4988 19836
rect 4939 19805 4951 19808
rect 4893 19799 4951 19805
rect 4982 19796 4988 19808
rect 5040 19796 5046 19848
rect 5261 19839 5319 19845
rect 5261 19805 5273 19839
rect 5307 19805 5319 19839
rect 5261 19799 5319 19805
rect 1854 19660 1860 19712
rect 1912 19700 1918 19712
rect 1949 19703 2007 19709
rect 1949 19700 1961 19703
rect 1912 19672 1961 19700
rect 1912 19660 1918 19672
rect 1949 19669 1961 19672
rect 1995 19669 2007 19703
rect 1949 19663 2007 19669
rect 2133 19703 2191 19709
rect 2133 19669 2145 19703
rect 2179 19700 2191 19703
rect 2777 19703 2835 19709
rect 2777 19700 2789 19703
rect 2179 19672 2789 19700
rect 2179 19669 2191 19672
rect 2133 19663 2191 19669
rect 2777 19669 2789 19672
rect 2823 19669 2835 19703
rect 2777 19663 2835 19669
rect 2961 19703 3019 19709
rect 2961 19669 2973 19703
rect 3007 19700 3019 19703
rect 3510 19700 3516 19712
rect 3007 19672 3516 19700
rect 3007 19669 3019 19672
rect 2961 19663 3019 19669
rect 3510 19660 3516 19672
rect 3568 19660 3574 19712
rect 4522 19660 4528 19712
rect 4580 19660 4586 19712
rect 5276 19700 5304 19799
rect 5902 19796 5908 19848
rect 5960 19836 5966 19848
rect 6365 19839 6423 19845
rect 6365 19836 6377 19839
rect 5960 19808 6377 19836
rect 5960 19796 5966 19808
rect 6365 19805 6377 19808
rect 6411 19805 6423 19839
rect 6365 19799 6423 19805
rect 6917 19839 6975 19845
rect 6917 19805 6929 19839
rect 6963 19805 6975 19839
rect 7116 19836 7144 19867
rect 7282 19864 7288 19916
rect 7340 19904 7346 19916
rect 7377 19907 7435 19913
rect 7377 19904 7389 19907
rect 7340 19876 7389 19904
rect 7340 19864 7346 19876
rect 7377 19873 7389 19876
rect 7423 19873 7435 19907
rect 7377 19867 7435 19873
rect 7650 19864 7656 19916
rect 7708 19904 7714 19916
rect 7745 19907 7803 19913
rect 7745 19904 7757 19907
rect 7708 19876 7757 19904
rect 7708 19864 7714 19876
rect 7745 19873 7757 19876
rect 7791 19873 7803 19907
rect 7745 19867 7803 19873
rect 7926 19864 7932 19916
rect 7984 19864 7990 19916
rect 8202 19864 8208 19916
rect 8260 19904 8266 19916
rect 8772 19913 8800 20012
rect 9766 20000 9772 20012
rect 9824 20000 9830 20052
rect 10134 20000 10140 20052
rect 10192 20040 10198 20052
rect 10321 20043 10379 20049
rect 10321 20040 10333 20043
rect 10192 20012 10333 20040
rect 10192 20000 10198 20012
rect 10321 20009 10333 20012
rect 10367 20009 10379 20043
rect 10321 20003 10379 20009
rect 10410 20000 10416 20052
rect 10468 20040 10474 20052
rect 10468 20012 11284 20040
rect 10468 20000 10474 20012
rect 8846 19932 8852 19984
rect 8904 19972 8910 19984
rect 9033 19975 9091 19981
rect 9033 19972 9045 19975
rect 8904 19944 9045 19972
rect 8904 19932 8910 19944
rect 9033 19941 9045 19944
rect 9079 19972 9091 19975
rect 10870 19972 10876 19984
rect 9079 19944 10876 19972
rect 9079 19941 9091 19944
rect 9033 19935 9091 19941
rect 10870 19932 10876 19944
rect 10928 19932 10934 19984
rect 11256 19972 11284 20012
rect 11422 20000 11428 20052
rect 11480 20000 11486 20052
rect 11514 20000 11520 20052
rect 11572 20000 11578 20052
rect 11790 20000 11796 20052
rect 11848 20040 11854 20052
rect 11848 20012 12020 20040
rect 11848 20000 11854 20012
rect 11256 19944 11836 19972
rect 8389 19907 8447 19913
rect 8389 19904 8401 19907
rect 8260 19876 8401 19904
rect 8260 19864 8266 19876
rect 8389 19873 8401 19876
rect 8435 19873 8447 19907
rect 8389 19867 8447 19873
rect 8573 19907 8631 19913
rect 8573 19873 8585 19907
rect 8619 19873 8631 19907
rect 8573 19867 8631 19873
rect 8757 19907 8815 19913
rect 8757 19873 8769 19907
rect 8803 19873 8815 19907
rect 8757 19867 8815 19873
rect 8941 19907 8999 19913
rect 8941 19873 8953 19907
rect 8987 19904 8999 19907
rect 8987 19876 9444 19904
rect 8987 19873 8999 19876
rect 8941 19867 8999 19873
rect 8478 19836 8484 19848
rect 7116 19808 8484 19836
rect 6917 19799 6975 19805
rect 5537 19771 5595 19777
rect 5537 19737 5549 19771
rect 5583 19768 5595 19771
rect 6932 19768 6960 19799
rect 8478 19796 8484 19808
rect 8536 19796 8542 19848
rect 8588 19836 8616 19867
rect 8846 19836 8852 19848
rect 8588 19808 8852 19836
rect 8846 19796 8852 19808
rect 8904 19796 8910 19848
rect 9416 19780 9444 19876
rect 9858 19864 9864 19916
rect 9916 19904 9922 19916
rect 10962 19904 10968 19916
rect 9916 19876 10968 19904
rect 9916 19864 9922 19876
rect 10962 19864 10968 19876
rect 11020 19864 11026 19916
rect 11256 19913 11284 19944
rect 11808 19913 11836 19944
rect 11992 19913 12020 20012
rect 13078 20000 13084 20052
rect 13136 20040 13142 20052
rect 13633 20043 13691 20049
rect 13633 20040 13645 20043
rect 13136 20012 13645 20040
rect 13136 20000 13142 20012
rect 13633 20009 13645 20012
rect 13679 20009 13691 20043
rect 13633 20003 13691 20009
rect 14366 20000 14372 20052
rect 14424 20040 14430 20052
rect 15197 20043 15255 20049
rect 15197 20040 15209 20043
rect 14424 20012 15209 20040
rect 14424 20000 14430 20012
rect 15197 20009 15209 20012
rect 15243 20009 15255 20043
rect 15197 20003 15255 20009
rect 15930 20000 15936 20052
rect 15988 20000 15994 20052
rect 16022 20000 16028 20052
rect 16080 20040 16086 20052
rect 16603 20043 16661 20049
rect 16080 20012 16436 20040
rect 16080 20000 16086 20012
rect 12268 19944 13768 19972
rect 11057 19907 11115 19913
rect 11057 19873 11069 19907
rect 11103 19873 11115 19907
rect 11057 19867 11115 19873
rect 11241 19907 11299 19913
rect 11241 19873 11253 19907
rect 11287 19873 11299 19907
rect 11241 19867 11299 19873
rect 11701 19907 11759 19913
rect 11701 19873 11713 19907
rect 11747 19873 11759 19907
rect 11701 19867 11759 19873
rect 11793 19907 11851 19913
rect 11793 19873 11805 19907
rect 11839 19873 11851 19907
rect 11793 19867 11851 19873
rect 11977 19907 12035 19913
rect 11977 19873 11989 19907
rect 12023 19873 12035 19907
rect 11977 19867 12035 19873
rect 9766 19796 9772 19848
rect 9824 19836 9830 19848
rect 11072 19836 11100 19867
rect 11716 19836 11744 19867
rect 12066 19864 12072 19916
rect 12124 19904 12130 19916
rect 12161 19907 12219 19913
rect 12161 19904 12173 19907
rect 12124 19876 12173 19904
rect 12124 19864 12130 19876
rect 12161 19873 12173 19876
rect 12207 19873 12219 19907
rect 12161 19867 12219 19873
rect 9824 19808 11744 19836
rect 9824 19796 9830 19808
rect 11882 19796 11888 19848
rect 11940 19836 11946 19848
rect 12268 19845 12296 19944
rect 12526 19913 12532 19916
rect 12520 19867 12532 19913
rect 12526 19864 12532 19867
rect 12584 19864 12590 19916
rect 13740 19913 13768 19944
rect 14734 19932 14740 19984
rect 14792 19972 14798 19984
rect 16408 19981 16436 20012
rect 16603 20009 16615 20043
rect 16649 20040 16661 20043
rect 16942 20040 16948 20052
rect 16649 20012 16948 20040
rect 16649 20009 16661 20012
rect 16603 20003 16661 20009
rect 16942 20000 16948 20012
rect 17000 20000 17006 20052
rect 17586 20000 17592 20052
rect 17644 20040 17650 20052
rect 19245 20043 19303 20049
rect 19245 20040 19257 20043
rect 17644 20012 19257 20040
rect 17644 20000 17650 20012
rect 19245 20009 19257 20012
rect 19291 20009 19303 20043
rect 19245 20003 19303 20009
rect 19518 20000 19524 20052
rect 19576 20040 19582 20052
rect 20346 20040 20352 20052
rect 19576 20012 20352 20040
rect 19576 20000 19582 20012
rect 20346 20000 20352 20012
rect 20404 20000 20410 20052
rect 20438 20000 20444 20052
rect 20496 20040 20502 20052
rect 21266 20040 21272 20052
rect 20496 20012 21272 20040
rect 20496 20000 20502 20012
rect 21266 20000 21272 20012
rect 21324 20000 21330 20052
rect 21358 20000 21364 20052
rect 21416 20040 21422 20052
rect 23017 20043 23075 20049
rect 23017 20040 23029 20043
rect 21416 20012 23029 20040
rect 21416 20000 21422 20012
rect 23017 20009 23029 20012
rect 23063 20009 23075 20043
rect 23017 20003 23075 20009
rect 16393 19975 16451 19981
rect 14792 19944 16160 19972
rect 14792 19932 14798 19944
rect 13725 19907 13783 19913
rect 13725 19873 13737 19907
rect 13771 19873 13783 19907
rect 13725 19867 13783 19873
rect 13814 19864 13820 19916
rect 13872 19904 13878 19916
rect 13981 19907 14039 19913
rect 13981 19904 13993 19907
rect 13872 19876 13993 19904
rect 13872 19864 13878 19876
rect 13981 19873 13993 19876
rect 14027 19873 14039 19907
rect 13981 19867 14039 19873
rect 15102 19864 15108 19916
rect 15160 19904 15166 19916
rect 15381 19907 15439 19913
rect 15381 19904 15393 19907
rect 15160 19876 15393 19904
rect 15160 19864 15166 19876
rect 15381 19873 15393 19876
rect 15427 19904 15439 19907
rect 15562 19904 15568 19916
rect 15427 19876 15568 19904
rect 15427 19873 15439 19876
rect 15381 19867 15439 19873
rect 15562 19864 15568 19876
rect 15620 19864 15626 19916
rect 15657 19907 15715 19913
rect 15657 19873 15669 19907
rect 15703 19873 15715 19907
rect 15657 19867 15715 19873
rect 15749 19907 15807 19913
rect 15749 19873 15761 19907
rect 15795 19904 15807 19907
rect 15838 19904 15844 19916
rect 15795 19876 15844 19904
rect 15795 19873 15807 19876
rect 15749 19867 15807 19873
rect 12253 19839 12311 19845
rect 12253 19836 12265 19839
rect 11940 19808 12265 19836
rect 11940 19796 11946 19808
rect 12253 19805 12265 19808
rect 12299 19805 12311 19839
rect 12253 19799 12311 19805
rect 14826 19796 14832 19848
rect 14884 19836 14890 19848
rect 15672 19836 15700 19867
rect 15838 19864 15844 19876
rect 15896 19864 15902 19916
rect 16132 19913 16160 19944
rect 16393 19941 16405 19975
rect 16439 19941 16451 19975
rect 17034 19972 17040 19984
rect 16393 19935 16451 19941
rect 16684 19944 17040 19972
rect 16117 19907 16175 19913
rect 16117 19873 16129 19907
rect 16163 19873 16175 19907
rect 16117 19867 16175 19873
rect 16301 19907 16359 19913
rect 16301 19873 16313 19907
rect 16347 19904 16359 19907
rect 16684 19904 16712 19944
rect 17034 19932 17040 19944
rect 17092 19972 17098 19984
rect 18690 19972 18696 19984
rect 17092 19944 18696 19972
rect 17092 19932 17098 19944
rect 18690 19932 18696 19944
rect 18748 19932 18754 19984
rect 23382 19972 23388 19984
rect 20548 19944 23388 19972
rect 16347 19876 16712 19904
rect 16347 19873 16359 19876
rect 16301 19867 16359 19873
rect 14884 19808 15700 19836
rect 16132 19836 16160 19867
rect 16758 19864 16764 19916
rect 16816 19904 16822 19916
rect 16853 19907 16911 19913
rect 16853 19904 16865 19907
rect 16816 19876 16865 19904
rect 16816 19864 16822 19876
rect 16853 19873 16865 19876
rect 16899 19873 16911 19907
rect 16853 19867 16911 19873
rect 19521 19907 19579 19913
rect 19521 19873 19533 19907
rect 19567 19904 19579 19907
rect 20162 19904 20168 19916
rect 19567 19876 20168 19904
rect 19567 19873 19579 19876
rect 19521 19867 19579 19873
rect 20162 19864 20168 19876
rect 20220 19864 20226 19916
rect 20349 19907 20407 19913
rect 20349 19873 20361 19907
rect 20395 19904 20407 19907
rect 20548 19904 20576 19944
rect 23382 19932 23388 19944
rect 23440 19932 23446 19984
rect 20395 19876 20576 19904
rect 20395 19873 20407 19876
rect 20349 19867 20407 19873
rect 20622 19864 20628 19916
rect 20680 19864 20686 19916
rect 20806 19864 20812 19916
rect 20864 19864 20870 19916
rect 21082 19864 21088 19916
rect 21140 19864 21146 19916
rect 21358 19864 21364 19916
rect 21416 19904 21422 19916
rect 21453 19907 21511 19913
rect 21453 19904 21465 19907
rect 21416 19876 21465 19904
rect 21416 19864 21422 19876
rect 21453 19873 21465 19876
rect 21499 19873 21511 19907
rect 21453 19867 21511 19873
rect 21634 19864 21640 19916
rect 21692 19864 21698 19916
rect 21726 19864 21732 19916
rect 21784 19904 21790 19916
rect 21893 19907 21951 19913
rect 21893 19904 21905 19907
rect 21784 19876 21905 19904
rect 21784 19864 21790 19876
rect 21893 19873 21905 19876
rect 21939 19873 21951 19907
rect 21893 19867 21951 19873
rect 18785 19839 18843 19845
rect 18785 19836 18797 19839
rect 16132 19808 18797 19836
rect 14884 19796 14890 19808
rect 18785 19805 18797 19808
rect 18831 19805 18843 19839
rect 18785 19799 18843 19805
rect 18877 19839 18935 19845
rect 18877 19805 18889 19839
rect 18923 19805 18935 19839
rect 18877 19799 18935 19805
rect 5583 19740 6960 19768
rect 5583 19737 5595 19740
rect 5537 19731 5595 19737
rect 7742 19728 7748 19780
rect 7800 19768 7806 19780
rect 7837 19771 7895 19777
rect 7837 19768 7849 19771
rect 7800 19740 7849 19768
rect 7800 19728 7806 19740
rect 7837 19737 7849 19740
rect 7883 19768 7895 19771
rect 9030 19768 9036 19780
rect 7883 19740 9036 19768
rect 7883 19737 7895 19740
rect 7837 19731 7895 19737
rect 9030 19728 9036 19740
rect 9088 19728 9094 19780
rect 9398 19728 9404 19780
rect 9456 19768 9462 19780
rect 9456 19740 12204 19768
rect 9456 19728 9462 19740
rect 6730 19700 6736 19712
rect 5276 19672 6736 19700
rect 6730 19660 6736 19672
rect 6788 19660 6794 19712
rect 7098 19660 7104 19712
rect 7156 19660 7162 19712
rect 7190 19660 7196 19712
rect 7248 19660 7254 19712
rect 8478 19660 8484 19712
rect 8536 19660 8542 19712
rect 8757 19703 8815 19709
rect 8757 19669 8769 19703
rect 8803 19700 8815 19703
rect 8938 19700 8944 19712
rect 8803 19672 8944 19700
rect 8803 19669 8815 19672
rect 8757 19663 8815 19669
rect 8938 19660 8944 19672
rect 8996 19660 9002 19712
rect 9674 19660 9680 19712
rect 9732 19700 9738 19712
rect 10410 19700 10416 19712
rect 9732 19672 10416 19700
rect 9732 19660 9738 19672
rect 10410 19660 10416 19672
rect 10468 19660 10474 19712
rect 12066 19660 12072 19712
rect 12124 19660 12130 19712
rect 12176 19700 12204 19740
rect 14918 19728 14924 19780
rect 14976 19768 14982 19780
rect 15473 19771 15531 19777
rect 15473 19768 15485 19771
rect 14976 19740 15485 19768
rect 14976 19728 14982 19740
rect 15473 19737 15485 19740
rect 15519 19737 15531 19771
rect 15473 19731 15531 19737
rect 16114 19728 16120 19780
rect 16172 19768 16178 19780
rect 16172 19740 18276 19768
rect 16172 19728 16178 19740
rect 14734 19700 14740 19712
rect 12176 19672 14740 19700
rect 14734 19660 14740 19672
rect 14792 19660 14798 19712
rect 15102 19660 15108 19712
rect 15160 19660 15166 19712
rect 15562 19660 15568 19712
rect 15620 19700 15626 19712
rect 16206 19700 16212 19712
rect 15620 19672 16212 19700
rect 15620 19660 15626 19672
rect 16206 19660 16212 19672
rect 16264 19660 16270 19712
rect 16298 19660 16304 19712
rect 16356 19660 16362 19712
rect 16574 19660 16580 19712
rect 16632 19660 16638 19712
rect 16761 19703 16819 19709
rect 16761 19669 16773 19703
rect 16807 19700 16819 19703
rect 17586 19700 17592 19712
rect 16807 19672 17592 19700
rect 16807 19669 16819 19672
rect 16761 19663 16819 19669
rect 17586 19660 17592 19672
rect 17644 19660 17650 19712
rect 18138 19660 18144 19712
rect 18196 19660 18202 19712
rect 18248 19700 18276 19740
rect 18690 19728 18696 19780
rect 18748 19768 18754 19780
rect 18892 19768 18920 19799
rect 18966 19796 18972 19848
rect 19024 19796 19030 19848
rect 19058 19796 19064 19848
rect 19116 19796 19122 19848
rect 19150 19796 19156 19848
rect 19208 19836 19214 19848
rect 19613 19839 19671 19845
rect 19613 19836 19625 19839
rect 19208 19808 19625 19836
rect 19208 19796 19214 19808
rect 19613 19805 19625 19808
rect 19659 19836 19671 19839
rect 19794 19836 19800 19848
rect 19659 19808 19800 19836
rect 19659 19805 19671 19808
rect 19613 19799 19671 19805
rect 19794 19796 19800 19808
rect 19852 19796 19858 19848
rect 20530 19796 20536 19848
rect 20588 19796 20594 19848
rect 20824 19836 20852 19864
rect 21174 19836 21180 19848
rect 20824 19808 21180 19836
rect 21174 19796 21180 19808
rect 21232 19836 21238 19848
rect 21232 19808 21404 19836
rect 21232 19796 21238 19808
rect 18748 19740 18920 19768
rect 19889 19771 19947 19777
rect 18748 19728 18754 19740
rect 19889 19737 19901 19771
rect 19935 19768 19947 19771
rect 20254 19768 20260 19780
rect 19935 19740 20260 19768
rect 19935 19737 19947 19740
rect 19889 19731 19947 19737
rect 20254 19728 20260 19740
rect 20312 19728 20318 19780
rect 20806 19728 20812 19780
rect 20864 19728 20870 19780
rect 21269 19771 21327 19777
rect 21269 19737 21281 19771
rect 21315 19768 21327 19771
rect 21376 19768 21404 19808
rect 21315 19740 21404 19768
rect 21315 19737 21327 19740
rect 21269 19731 21327 19737
rect 20165 19703 20223 19709
rect 20165 19700 20177 19703
rect 18248 19672 20177 19700
rect 20165 19669 20177 19672
rect 20211 19669 20223 19703
rect 20165 19663 20223 19669
rect 20530 19660 20536 19712
rect 20588 19700 20594 19712
rect 20901 19703 20959 19709
rect 20901 19700 20913 19703
rect 20588 19672 20913 19700
rect 20588 19660 20594 19672
rect 20901 19669 20913 19672
rect 20947 19669 20959 19703
rect 20901 19663 20959 19669
rect 552 19610 23368 19632
rect 552 19558 1366 19610
rect 1418 19558 1430 19610
rect 1482 19558 1494 19610
rect 1546 19558 1558 19610
rect 1610 19558 1622 19610
rect 1674 19558 1686 19610
rect 1738 19558 7366 19610
rect 7418 19558 7430 19610
rect 7482 19558 7494 19610
rect 7546 19558 7558 19610
rect 7610 19558 7622 19610
rect 7674 19558 7686 19610
rect 7738 19558 13366 19610
rect 13418 19558 13430 19610
rect 13482 19558 13494 19610
rect 13546 19558 13558 19610
rect 13610 19558 13622 19610
rect 13674 19558 13686 19610
rect 13738 19558 19366 19610
rect 19418 19558 19430 19610
rect 19482 19558 19494 19610
rect 19546 19558 19558 19610
rect 19610 19558 19622 19610
rect 19674 19558 19686 19610
rect 19738 19558 23368 19610
rect 552 19536 23368 19558
rect 2869 19499 2927 19505
rect 2869 19465 2881 19499
rect 2915 19496 2927 19499
rect 3326 19496 3332 19508
rect 2915 19468 3332 19496
rect 2915 19465 2927 19468
rect 2869 19459 2927 19465
rect 3326 19456 3332 19468
rect 3384 19456 3390 19508
rect 3418 19456 3424 19508
rect 3476 19496 3482 19508
rect 3513 19499 3571 19505
rect 3513 19496 3525 19499
rect 3476 19468 3525 19496
rect 3476 19456 3482 19468
rect 3513 19465 3525 19468
rect 3559 19465 3571 19499
rect 3513 19459 3571 19465
rect 4893 19499 4951 19505
rect 4893 19465 4905 19499
rect 4939 19496 4951 19499
rect 4982 19496 4988 19508
rect 4939 19468 4988 19496
rect 4939 19465 4951 19468
rect 4893 19459 4951 19465
rect 4982 19456 4988 19468
rect 5040 19456 5046 19508
rect 5353 19499 5411 19505
rect 5353 19465 5365 19499
rect 5399 19496 5411 19499
rect 5442 19496 5448 19508
rect 5399 19468 5448 19496
rect 5399 19465 5411 19468
rect 5353 19459 5411 19465
rect 2498 19388 2504 19440
rect 2556 19428 2562 19440
rect 3789 19431 3847 19437
rect 3789 19428 3801 19431
rect 2556 19400 3801 19428
rect 2556 19388 2562 19400
rect 3789 19397 3801 19400
rect 3835 19397 3847 19431
rect 3789 19391 3847 19397
rect 4617 19431 4675 19437
rect 4617 19397 4629 19431
rect 4663 19428 4675 19431
rect 5258 19428 5264 19440
rect 4663 19400 5264 19428
rect 4663 19397 4675 19400
rect 4617 19391 4675 19397
rect 566 19320 572 19372
rect 624 19360 630 19372
rect 845 19363 903 19369
rect 845 19360 857 19363
rect 624 19332 857 19360
rect 624 19320 630 19332
rect 845 19329 857 19332
rect 891 19329 903 19363
rect 4632 19360 4660 19391
rect 5258 19388 5264 19400
rect 5316 19388 5322 19440
rect 2792 19334 3924 19360
rect 845 19323 903 19329
rect 2700 19332 3924 19334
rect 2700 19306 2820 19332
rect 1673 19295 1731 19301
rect 1673 19261 1685 19295
rect 1719 19292 1731 19295
rect 1762 19292 1768 19304
rect 1719 19264 1768 19292
rect 1719 19261 1731 19264
rect 1673 19255 1731 19261
rect 1762 19252 1768 19264
rect 1820 19252 1826 19304
rect 1854 19252 1860 19304
rect 1912 19252 1918 19304
rect 2222 19252 2228 19304
rect 2280 19252 2286 19304
rect 2406 19252 2412 19304
rect 2464 19252 2470 19304
rect 2424 19224 2452 19252
rect 2700 19224 2728 19306
rect 3418 19252 3424 19304
rect 3476 19252 3482 19304
rect 3510 19252 3516 19304
rect 3568 19292 3574 19304
rect 3697 19295 3755 19301
rect 3697 19292 3709 19295
rect 3568 19264 3709 19292
rect 3568 19252 3574 19264
rect 3697 19261 3709 19264
rect 3743 19261 3755 19295
rect 3697 19255 3755 19261
rect 3786 19252 3792 19304
rect 3844 19252 3850 19304
rect 3896 19292 3924 19332
rect 4356 19332 4660 19360
rect 3970 19292 3976 19304
rect 3896 19264 3976 19292
rect 3970 19252 3976 19264
rect 4028 19252 4034 19304
rect 4062 19252 4068 19304
rect 4120 19292 4126 19304
rect 4356 19301 4384 19332
rect 4157 19295 4215 19301
rect 4157 19292 4169 19295
rect 4120 19264 4169 19292
rect 4120 19252 4126 19264
rect 4157 19261 4169 19264
rect 4203 19261 4215 19295
rect 4157 19255 4215 19261
rect 4341 19295 4399 19301
rect 4341 19261 4353 19295
rect 4387 19261 4399 19295
rect 4341 19255 4399 19261
rect 4433 19295 4491 19301
rect 4433 19261 4445 19295
rect 4479 19261 4491 19295
rect 4433 19255 4491 19261
rect 2424 19196 2728 19224
rect 2958 19184 2964 19236
rect 3016 19224 3022 19236
rect 4448 19224 4476 19255
rect 4522 19252 4528 19304
rect 4580 19292 4586 19304
rect 4709 19295 4767 19301
rect 4709 19292 4721 19295
rect 4580 19264 4721 19292
rect 4580 19252 4586 19264
rect 4709 19261 4721 19264
rect 4755 19261 4767 19295
rect 4709 19255 4767 19261
rect 5169 19295 5227 19301
rect 5169 19261 5181 19295
rect 5215 19292 5227 19295
rect 5368 19292 5396 19459
rect 5442 19456 5448 19468
rect 5500 19456 5506 19508
rect 5534 19456 5540 19508
rect 5592 19496 5598 19508
rect 8662 19496 8668 19508
rect 5592 19468 8668 19496
rect 5592 19456 5598 19468
rect 8662 19456 8668 19468
rect 8720 19456 8726 19508
rect 8757 19499 8815 19505
rect 8757 19465 8769 19499
rect 8803 19496 8815 19499
rect 8846 19496 8852 19508
rect 8803 19468 8852 19496
rect 8803 19465 8815 19468
rect 8757 19459 8815 19465
rect 8846 19456 8852 19468
rect 8904 19456 8910 19508
rect 9766 19456 9772 19508
rect 9824 19496 9830 19508
rect 10137 19499 10195 19505
rect 10137 19496 10149 19499
rect 9824 19468 10149 19496
rect 9824 19456 9830 19468
rect 10137 19465 10149 19468
rect 10183 19465 10195 19499
rect 10137 19459 10195 19465
rect 10410 19456 10416 19508
rect 10468 19456 10474 19508
rect 11425 19499 11483 19505
rect 11425 19465 11437 19499
rect 11471 19496 11483 19499
rect 12069 19499 12127 19505
rect 12069 19496 12081 19499
rect 11471 19468 12081 19496
rect 11471 19465 11483 19468
rect 11425 19459 11483 19465
rect 12069 19465 12081 19468
rect 12115 19465 12127 19499
rect 12069 19459 12127 19465
rect 12802 19456 12808 19508
rect 12860 19496 12866 19508
rect 12897 19499 12955 19505
rect 12897 19496 12909 19499
rect 12860 19468 12909 19496
rect 12860 19456 12866 19468
rect 12897 19465 12909 19468
rect 12943 19465 12955 19499
rect 12897 19459 12955 19465
rect 13725 19499 13783 19505
rect 13725 19465 13737 19499
rect 13771 19496 13783 19499
rect 13814 19496 13820 19508
rect 13771 19468 13820 19496
rect 13771 19465 13783 19468
rect 13725 19459 13783 19465
rect 8941 19431 8999 19437
rect 8941 19397 8953 19431
rect 8987 19428 8999 19431
rect 8987 19400 9904 19428
rect 8987 19397 8999 19400
rect 8941 19391 8999 19397
rect 7926 19320 7932 19372
rect 7984 19360 7990 19372
rect 8202 19360 8208 19372
rect 7984 19332 8208 19360
rect 7984 19320 7990 19332
rect 8202 19320 8208 19332
rect 8260 19360 8266 19372
rect 8260 19334 8432 19360
rect 8260 19332 8616 19334
rect 8260 19320 8266 19332
rect 8404 19306 8616 19332
rect 9398 19320 9404 19372
rect 9456 19320 9462 19372
rect 9582 19320 9588 19372
rect 9640 19360 9646 19372
rect 9674 19360 9680 19372
rect 9640 19332 9680 19360
rect 9640 19320 9646 19332
rect 9674 19320 9680 19332
rect 9732 19320 9738 19372
rect 9876 19360 9904 19400
rect 10778 19388 10784 19440
rect 10836 19428 10842 19440
rect 11882 19428 11888 19440
rect 10836 19400 11888 19428
rect 10836 19388 10842 19400
rect 11882 19388 11888 19400
rect 11940 19388 11946 19440
rect 12912 19428 12940 19459
rect 13814 19456 13820 19468
rect 13872 19456 13878 19508
rect 14366 19456 14372 19508
rect 14424 19456 14430 19508
rect 14553 19499 14611 19505
rect 14553 19465 14565 19499
rect 14599 19496 14611 19499
rect 14826 19496 14832 19508
rect 14599 19468 14832 19496
rect 14599 19465 14611 19468
rect 14553 19459 14611 19465
rect 14826 19456 14832 19468
rect 14884 19456 14890 19508
rect 15286 19456 15292 19508
rect 15344 19496 15350 19508
rect 20438 19496 20444 19508
rect 15344 19468 20444 19496
rect 15344 19456 15350 19468
rect 20438 19456 20444 19468
rect 20496 19456 20502 19508
rect 20714 19456 20720 19508
rect 20772 19456 20778 19508
rect 20809 19499 20867 19505
rect 20809 19465 20821 19499
rect 20855 19465 20867 19499
rect 20809 19459 20867 19465
rect 21637 19499 21695 19505
rect 21637 19465 21649 19499
rect 21683 19465 21695 19499
rect 21637 19459 21695 19465
rect 14384 19428 14412 19456
rect 12912 19400 14412 19428
rect 16025 19431 16083 19437
rect 16025 19397 16037 19431
rect 16071 19397 16083 19431
rect 16025 19391 16083 19397
rect 10502 19360 10508 19372
rect 9876 19332 10180 19360
rect 5215 19264 5396 19292
rect 6733 19295 6791 19301
rect 5215 19261 5227 19264
rect 5169 19255 5227 19261
rect 6733 19261 6745 19295
rect 6779 19292 6791 19295
rect 6822 19292 6828 19304
rect 6779 19264 6828 19292
rect 6779 19261 6791 19264
rect 6733 19255 6791 19261
rect 4724 19224 4752 19255
rect 6822 19252 6828 19264
rect 6880 19252 6886 19304
rect 5810 19224 5816 19236
rect 3016 19196 3188 19224
rect 4448 19196 4568 19224
rect 4724 19196 5816 19224
rect 3016 19184 3022 19196
rect 2409 19159 2467 19165
rect 2409 19125 2421 19159
rect 2455 19156 2467 19159
rect 2869 19159 2927 19165
rect 2869 19156 2881 19159
rect 2455 19128 2881 19156
rect 2455 19125 2467 19128
rect 2409 19119 2467 19125
rect 2869 19125 2881 19128
rect 2915 19125 2927 19159
rect 2869 19119 2927 19125
rect 3050 19116 3056 19168
rect 3108 19116 3114 19168
rect 3160 19156 3188 19196
rect 3237 19159 3295 19165
rect 3237 19156 3249 19159
rect 3160 19128 3249 19156
rect 3237 19125 3249 19128
rect 3283 19125 3295 19159
rect 3237 19119 3295 19125
rect 4246 19116 4252 19168
rect 4304 19116 4310 19168
rect 4540 19156 4568 19196
rect 5810 19184 5816 19196
rect 5868 19224 5874 19236
rect 6362 19224 6368 19236
rect 5868 19196 6368 19224
rect 5868 19184 5874 19196
rect 6362 19184 6368 19196
rect 6420 19184 6426 19236
rect 6488 19227 6546 19233
rect 6488 19193 6500 19227
rect 6534 19224 6546 19227
rect 6914 19224 6920 19236
rect 6534 19196 6920 19224
rect 6534 19193 6546 19196
rect 6488 19187 6546 19193
rect 6914 19184 6920 19196
rect 6972 19184 6978 19236
rect 7092 19227 7150 19233
rect 7092 19193 7104 19227
rect 7138 19224 7150 19227
rect 7190 19224 7196 19236
rect 7138 19196 7196 19224
rect 7138 19193 7150 19196
rect 7092 19187 7150 19193
rect 7190 19184 7196 19196
rect 7248 19184 7254 19236
rect 8588 19233 8616 19306
rect 9493 19295 9551 19301
rect 9493 19261 9505 19295
rect 9539 19292 9551 19295
rect 9858 19292 9864 19304
rect 9539 19264 9864 19292
rect 9539 19261 9551 19264
rect 9493 19255 9551 19261
rect 9858 19252 9864 19264
rect 9916 19252 9922 19304
rect 9950 19252 9956 19304
rect 10008 19252 10014 19304
rect 10042 19252 10048 19304
rect 10100 19252 10106 19304
rect 10152 19292 10180 19332
rect 10428 19332 10508 19360
rect 10321 19295 10379 19301
rect 10321 19292 10333 19295
rect 10152 19264 10333 19292
rect 8573 19227 8631 19233
rect 8573 19193 8585 19227
rect 8619 19193 8631 19227
rect 8573 19187 8631 19193
rect 8662 19184 8668 19236
rect 8720 19224 8726 19236
rect 8720 19196 9168 19224
rect 8720 19184 8726 19196
rect 4798 19156 4804 19168
rect 4540 19128 4804 19156
rect 4798 19116 4804 19128
rect 4856 19116 4862 19168
rect 4985 19159 5043 19165
rect 4985 19125 4997 19159
rect 5031 19156 5043 19159
rect 5166 19156 5172 19168
rect 5031 19128 5172 19156
rect 5031 19125 5043 19128
rect 4985 19119 5043 19125
rect 5166 19116 5172 19128
rect 5224 19116 5230 19168
rect 8202 19116 8208 19168
rect 8260 19116 8266 19168
rect 8754 19116 8760 19168
rect 8812 19165 8818 19168
rect 8812 19159 8831 19165
rect 8819 19125 8831 19159
rect 8812 19119 8831 19125
rect 8812 19116 8818 19119
rect 9030 19116 9036 19168
rect 9088 19116 9094 19168
rect 9140 19156 9168 19196
rect 9214 19184 9220 19236
rect 9272 19224 9278 19236
rect 10134 19224 10140 19236
rect 9272 19196 10140 19224
rect 9272 19184 9278 19196
rect 10134 19184 10140 19196
rect 10192 19184 10198 19236
rect 10244 19224 10272 19264
rect 10321 19261 10333 19264
rect 10367 19261 10379 19295
rect 10428 19292 10456 19332
rect 10502 19320 10508 19332
rect 10560 19320 10566 19372
rect 11790 19320 11796 19372
rect 11848 19360 11854 19372
rect 12529 19363 12587 19369
rect 12529 19360 12541 19363
rect 11848 19332 12541 19360
rect 11848 19320 11854 19332
rect 12529 19329 12541 19332
rect 12575 19329 12587 19363
rect 12529 19323 12587 19329
rect 13464 19332 13676 19360
rect 10597 19295 10655 19301
rect 10597 19292 10609 19295
rect 10428 19264 10609 19292
rect 10321 19255 10379 19261
rect 10597 19261 10609 19264
rect 10643 19261 10655 19295
rect 13464 19292 13492 19332
rect 10597 19255 10655 19261
rect 10704 19264 13492 19292
rect 13541 19295 13599 19301
rect 10704 19224 10732 19264
rect 13541 19261 13553 19295
rect 13587 19261 13599 19295
rect 13541 19255 13599 19261
rect 10244 19196 10732 19224
rect 11609 19227 11667 19233
rect 11609 19193 11621 19227
rect 11655 19193 11667 19227
rect 11609 19187 11667 19193
rect 9677 19159 9735 19165
rect 9677 19156 9689 19159
rect 9140 19128 9689 19156
rect 9677 19125 9689 19128
rect 9723 19125 9735 19159
rect 9677 19119 9735 19125
rect 9858 19116 9864 19168
rect 9916 19156 9922 19168
rect 11146 19156 11152 19168
rect 9916 19128 11152 19156
rect 9916 19116 9922 19128
rect 11146 19116 11152 19128
rect 11204 19116 11210 19168
rect 11624 19156 11652 19187
rect 11790 19184 11796 19236
rect 11848 19184 11854 19236
rect 11882 19184 11888 19236
rect 11940 19184 11946 19236
rect 12066 19184 12072 19236
rect 12124 19233 12130 19236
rect 12124 19227 12143 19233
rect 12131 19193 12143 19227
rect 12124 19187 12143 19193
rect 12124 19184 12130 19187
rect 11974 19156 11980 19168
rect 11624 19128 11980 19156
rect 11974 19116 11980 19128
rect 12032 19116 12038 19168
rect 12253 19159 12311 19165
rect 12253 19125 12265 19159
rect 12299 19156 12311 19159
rect 12434 19156 12440 19168
rect 12299 19128 12440 19156
rect 12299 19125 12311 19128
rect 12253 19119 12311 19125
rect 12434 19116 12440 19128
rect 12492 19116 12498 19168
rect 12894 19116 12900 19168
rect 12952 19116 12958 19168
rect 13081 19159 13139 19165
rect 13081 19125 13093 19159
rect 13127 19156 13139 19159
rect 13556 19156 13584 19255
rect 13648 19224 13676 19332
rect 13998 19252 14004 19304
rect 14056 19252 14062 19304
rect 14645 19295 14703 19301
rect 14645 19261 14657 19295
rect 14691 19292 14703 19295
rect 15194 19292 15200 19304
rect 14691 19264 15200 19292
rect 14691 19261 14703 19264
rect 14645 19255 14703 19261
rect 15194 19252 15200 19264
rect 15252 19252 15258 19304
rect 16040 19292 16068 19391
rect 20254 19388 20260 19440
rect 20312 19428 20318 19440
rect 20824 19428 20852 19459
rect 20312 19400 20852 19428
rect 20312 19388 20318 19400
rect 18138 19360 18144 19372
rect 17512 19332 18144 19360
rect 15580 19264 16068 19292
rect 15580 19236 15608 19264
rect 16114 19252 16120 19304
rect 16172 19292 16178 19304
rect 17512 19292 17540 19332
rect 18138 19320 18144 19332
rect 18196 19320 18202 19372
rect 20441 19363 20499 19369
rect 20441 19329 20453 19363
rect 20487 19329 20499 19363
rect 20441 19323 20499 19329
rect 16172 19264 17540 19292
rect 17589 19295 17647 19301
rect 16172 19252 16178 19264
rect 17589 19261 17601 19295
rect 17635 19261 17647 19295
rect 17589 19255 17647 19261
rect 14918 19233 14924 19236
rect 14912 19224 14924 19233
rect 13648 19196 14780 19224
rect 14879 19196 14924 19224
rect 13127 19128 13584 19156
rect 13127 19125 13139 19128
rect 13081 19119 13139 19125
rect 14366 19116 14372 19168
rect 14424 19116 14430 19168
rect 14752 19156 14780 19196
rect 14912 19187 14924 19196
rect 14918 19184 14924 19187
rect 14976 19184 14982 19236
rect 15562 19184 15568 19236
rect 15620 19184 15626 19236
rect 15746 19184 15752 19236
rect 15804 19224 15810 19236
rect 16362 19227 16420 19233
rect 16362 19224 16374 19227
rect 15804 19196 16374 19224
rect 15804 19184 15810 19196
rect 16362 19193 16374 19196
rect 16408 19193 16420 19227
rect 16362 19187 16420 19193
rect 16482 19184 16488 19236
rect 16540 19224 16546 19236
rect 17604 19224 17632 19255
rect 17862 19252 17868 19304
rect 17920 19252 17926 19304
rect 18156 19292 18184 19320
rect 18506 19292 18512 19304
rect 18156 19264 18512 19292
rect 18506 19252 18512 19264
rect 18564 19292 18570 19304
rect 18693 19295 18751 19301
rect 18693 19292 18705 19295
rect 18564 19264 18705 19292
rect 18564 19252 18570 19264
rect 18693 19261 18705 19264
rect 18739 19261 18751 19295
rect 18693 19255 18751 19261
rect 18708 19224 18736 19255
rect 20254 19252 20260 19304
rect 20312 19292 20318 19304
rect 20349 19295 20407 19301
rect 20349 19292 20361 19295
rect 20312 19264 20361 19292
rect 20312 19252 20318 19264
rect 20349 19261 20361 19264
rect 20395 19261 20407 19295
rect 20456 19292 20484 19323
rect 20530 19320 20536 19372
rect 20588 19360 20594 19372
rect 21174 19360 21180 19372
rect 20588 19332 21180 19360
rect 20588 19320 20594 19332
rect 21174 19320 21180 19332
rect 21232 19320 21238 19372
rect 21652 19360 21680 19459
rect 22002 19456 22008 19508
rect 22060 19496 22066 19508
rect 22741 19499 22799 19505
rect 22741 19496 22753 19499
rect 22060 19468 22753 19496
rect 22060 19456 22066 19468
rect 22741 19465 22753 19468
rect 22787 19465 22799 19499
rect 22741 19459 22799 19465
rect 21818 19388 21824 19440
rect 21876 19428 21882 19440
rect 21876 19400 22232 19428
rect 21876 19388 21882 19400
rect 21726 19360 21732 19372
rect 21652 19332 21732 19360
rect 21726 19320 21732 19332
rect 21784 19320 21790 19372
rect 22204 19369 22232 19400
rect 22005 19363 22063 19369
rect 22005 19360 22017 19363
rect 21928 19334 22017 19360
rect 21919 19332 22017 19334
rect 21919 19306 21956 19332
rect 22005 19329 22017 19332
rect 22051 19329 22063 19363
rect 22005 19323 22063 19329
rect 22189 19363 22247 19369
rect 22189 19329 22201 19363
rect 22235 19329 22247 19363
rect 22189 19323 22247 19329
rect 20622 19292 20628 19304
rect 20456 19264 20628 19292
rect 20349 19255 20407 19261
rect 20622 19252 20628 19264
rect 20680 19252 20686 19304
rect 20714 19252 20720 19304
rect 20772 19292 20778 19304
rect 20809 19295 20867 19301
rect 20809 19292 20821 19295
rect 20772 19264 20821 19292
rect 20772 19252 20778 19264
rect 20809 19261 20821 19264
rect 20855 19261 20867 19295
rect 20809 19255 20867 19261
rect 20990 19252 20996 19304
rect 21048 19252 21054 19304
rect 21082 19252 21088 19304
rect 21140 19292 21146 19304
rect 21453 19295 21511 19301
rect 21453 19292 21465 19295
rect 21140 19264 21465 19292
rect 21140 19252 21146 19264
rect 21453 19261 21465 19264
rect 21499 19261 21511 19295
rect 21453 19255 21511 19261
rect 21542 19252 21548 19304
rect 21600 19292 21606 19304
rect 21821 19295 21879 19301
rect 21821 19292 21833 19295
rect 21600 19264 21833 19292
rect 21600 19252 21606 19264
rect 18782 19224 18788 19236
rect 16540 19196 18644 19224
rect 18708 19196 18788 19224
rect 16540 19184 16546 19196
rect 16574 19156 16580 19168
rect 14752 19128 16580 19156
rect 16574 19116 16580 19128
rect 16632 19156 16638 19168
rect 16850 19156 16856 19168
rect 16632 19128 16856 19156
rect 16632 19116 16638 19128
rect 16850 19116 16856 19128
rect 16908 19116 16914 19168
rect 17497 19159 17555 19165
rect 17497 19125 17509 19159
rect 17543 19156 17555 19159
rect 17678 19156 17684 19168
rect 17543 19128 17684 19156
rect 17543 19125 17555 19128
rect 17497 19119 17555 19125
rect 17678 19116 17684 19128
rect 17736 19116 17742 19168
rect 18616 19156 18644 19196
rect 18782 19184 18788 19196
rect 18840 19184 18846 19236
rect 18966 19233 18972 19236
rect 18960 19187 18972 19233
rect 18966 19184 18972 19187
rect 19024 19184 19030 19236
rect 19058 19184 19064 19236
rect 19116 19224 19122 19236
rect 19116 19196 20208 19224
rect 19116 19184 19122 19196
rect 19242 19156 19248 19168
rect 18616 19128 19248 19156
rect 19242 19116 19248 19128
rect 19300 19116 19306 19168
rect 19426 19116 19432 19168
rect 19484 19156 19490 19168
rect 19702 19156 19708 19168
rect 19484 19128 19708 19156
rect 19484 19116 19490 19128
rect 19702 19116 19708 19128
rect 19760 19156 19766 19168
rect 20073 19159 20131 19165
rect 20073 19156 20085 19159
rect 19760 19128 20085 19156
rect 19760 19116 19766 19128
rect 20073 19125 20085 19128
rect 20119 19125 20131 19159
rect 20180 19156 20208 19196
rect 20364 19196 21220 19224
rect 20364 19156 20392 19196
rect 21192 19165 21220 19196
rect 20180 19128 20392 19156
rect 21177 19159 21235 19165
rect 20073 19119 20131 19125
rect 21177 19125 21189 19159
rect 21223 19125 21235 19159
rect 21177 19119 21235 19125
rect 21269 19159 21327 19165
rect 21269 19125 21281 19159
rect 21315 19156 21327 19159
rect 21358 19156 21364 19168
rect 21315 19128 21364 19156
rect 21315 19125 21327 19128
rect 21269 19119 21327 19125
rect 21358 19116 21364 19128
rect 21416 19116 21422 19168
rect 21652 19156 21680 19264
rect 21821 19261 21833 19264
rect 21867 19261 21879 19295
rect 21821 19255 21879 19261
rect 21726 19184 21732 19236
rect 21784 19224 21790 19236
rect 21919 19224 21947 19306
rect 22094 19252 22100 19304
rect 22152 19252 22158 19304
rect 22373 19295 22431 19301
rect 22373 19261 22385 19295
rect 22419 19261 22431 19295
rect 22373 19255 22431 19261
rect 21784 19196 21947 19224
rect 21784 19184 21790 19196
rect 22388 19168 22416 19255
rect 22462 19252 22468 19304
rect 22520 19292 22526 19304
rect 22833 19295 22891 19301
rect 22833 19292 22845 19295
rect 22520 19264 22845 19292
rect 22520 19252 22526 19264
rect 22833 19261 22845 19264
rect 22879 19261 22891 19295
rect 22833 19255 22891 19261
rect 22002 19156 22008 19168
rect 21652 19128 22008 19156
rect 22002 19116 22008 19128
rect 22060 19156 22066 19168
rect 22186 19156 22192 19168
rect 22060 19128 22192 19156
rect 22060 19116 22066 19128
rect 22186 19116 22192 19128
rect 22244 19116 22250 19168
rect 22370 19116 22376 19168
rect 22428 19116 22434 19168
rect 22557 19159 22615 19165
rect 22557 19125 22569 19159
rect 22603 19156 22615 19159
rect 23106 19156 23112 19168
rect 22603 19128 23112 19156
rect 22603 19125 22615 19128
rect 22557 19119 22615 19125
rect 23106 19116 23112 19128
rect 23164 19116 23170 19168
rect 552 19066 23368 19088
rect 552 19014 4366 19066
rect 4418 19014 4430 19066
rect 4482 19014 4494 19066
rect 4546 19014 4558 19066
rect 4610 19014 4622 19066
rect 4674 19014 4686 19066
rect 4738 19014 10366 19066
rect 10418 19014 10430 19066
rect 10482 19014 10494 19066
rect 10546 19014 10558 19066
rect 10610 19014 10622 19066
rect 10674 19014 10686 19066
rect 10738 19014 16366 19066
rect 16418 19014 16430 19066
rect 16482 19014 16494 19066
rect 16546 19014 16558 19066
rect 16610 19014 16622 19066
rect 16674 19014 16686 19066
rect 16738 19014 22366 19066
rect 22418 19014 22430 19066
rect 22482 19014 22494 19066
rect 22546 19014 22558 19066
rect 22610 19014 22622 19066
rect 22674 19014 22686 19066
rect 22738 19014 23368 19066
rect 552 18992 23368 19014
rect 3050 18952 3056 18964
rect 2700 18924 3056 18952
rect 1857 18819 1915 18825
rect 1857 18785 1869 18819
rect 1903 18816 1915 18819
rect 2406 18816 2412 18828
rect 1903 18788 2412 18816
rect 1903 18785 1915 18788
rect 1857 18779 1915 18785
rect 2406 18776 2412 18788
rect 2464 18776 2470 18828
rect 2700 18825 2728 18924
rect 3050 18912 3056 18924
rect 3108 18912 3114 18964
rect 3234 18912 3240 18964
rect 3292 18912 3298 18964
rect 3970 18912 3976 18964
rect 4028 18952 4034 18964
rect 6178 18952 6184 18964
rect 4028 18924 6184 18952
rect 4028 18912 4034 18924
rect 6178 18912 6184 18924
rect 6236 18912 6242 18964
rect 7282 18912 7288 18964
rect 7340 18952 7346 18964
rect 7653 18955 7711 18961
rect 7653 18952 7665 18955
rect 7340 18924 7665 18952
rect 7340 18912 7346 18924
rect 7653 18921 7665 18924
rect 7699 18921 7711 18955
rect 7653 18915 7711 18921
rect 8757 18955 8815 18961
rect 8757 18921 8769 18955
rect 8803 18952 8815 18955
rect 9306 18952 9312 18964
rect 8803 18924 9312 18952
rect 8803 18921 8815 18924
rect 8757 18915 8815 18921
rect 9306 18912 9312 18924
rect 9364 18912 9370 18964
rect 10042 18912 10048 18964
rect 10100 18952 10106 18964
rect 10100 18924 12480 18952
rect 10100 18912 10106 18924
rect 3252 18884 3280 18912
rect 2976 18856 3280 18884
rect 2976 18825 3004 18856
rect 4890 18844 4896 18896
rect 4948 18884 4954 18896
rect 5258 18884 5264 18896
rect 4948 18856 5264 18884
rect 4948 18844 4954 18856
rect 5258 18844 5264 18856
rect 5316 18884 5322 18896
rect 7834 18884 7840 18896
rect 5316 18856 5396 18884
rect 5316 18844 5322 18856
rect 2685 18819 2743 18825
rect 2685 18785 2697 18819
rect 2731 18785 2743 18819
rect 2685 18779 2743 18785
rect 2961 18819 3019 18825
rect 2961 18785 2973 18819
rect 3007 18785 3019 18819
rect 3217 18819 3275 18825
rect 3217 18816 3229 18819
rect 2961 18779 3019 18785
rect 3068 18788 3229 18816
rect 1946 18708 1952 18760
rect 2004 18708 2010 18760
rect 2501 18751 2559 18757
rect 2501 18717 2513 18751
rect 2547 18748 2559 18751
rect 2590 18748 2596 18760
rect 2547 18720 2596 18748
rect 2547 18717 2559 18720
rect 2501 18711 2559 18717
rect 2590 18708 2596 18720
rect 2648 18708 2654 18760
rect 3068 18748 3096 18788
rect 3217 18785 3229 18788
rect 3263 18785 3275 18819
rect 3217 18779 3275 18785
rect 4617 18819 4675 18825
rect 4617 18785 4629 18819
rect 4663 18816 4675 18819
rect 4982 18816 4988 18828
rect 4663 18788 4988 18816
rect 4663 18785 4675 18788
rect 4617 18779 4675 18785
rect 4982 18776 4988 18788
rect 5040 18776 5046 18828
rect 5077 18819 5135 18825
rect 5077 18785 5089 18819
rect 5123 18816 5135 18819
rect 5166 18816 5172 18828
rect 5123 18788 5172 18816
rect 5123 18785 5135 18788
rect 5077 18779 5135 18785
rect 5166 18776 5172 18788
rect 5224 18776 5230 18828
rect 5368 18825 5396 18856
rect 6564 18856 7840 18884
rect 5353 18819 5411 18825
rect 5353 18785 5365 18819
rect 5399 18816 5411 18819
rect 5626 18816 5632 18828
rect 5399 18788 5632 18816
rect 5399 18785 5411 18788
rect 5353 18779 5411 18785
rect 5626 18776 5632 18788
rect 5684 18776 5690 18828
rect 5810 18776 5816 18828
rect 5868 18825 5874 18828
rect 5868 18816 5877 18825
rect 5997 18819 6055 18825
rect 5868 18788 5913 18816
rect 5868 18779 5877 18788
rect 5997 18785 6009 18819
rect 6043 18816 6055 18819
rect 6273 18819 6331 18825
rect 6273 18816 6285 18819
rect 6043 18788 6285 18816
rect 6043 18785 6055 18788
rect 5997 18779 6055 18785
rect 6273 18785 6285 18788
rect 6319 18816 6331 18819
rect 6564 18816 6592 18856
rect 7834 18844 7840 18856
rect 7892 18844 7898 18896
rect 8478 18844 8484 18896
rect 8536 18844 8542 18896
rect 8662 18844 8668 18896
rect 8720 18884 8726 18896
rect 8720 18856 8892 18884
rect 8720 18844 8726 18856
rect 6319 18788 6592 18816
rect 7285 18819 7343 18825
rect 6319 18785 6331 18788
rect 6273 18779 6331 18785
rect 7285 18785 7297 18819
rect 7331 18816 7343 18819
rect 7745 18819 7803 18825
rect 7745 18816 7757 18819
rect 7331 18788 7757 18816
rect 7331 18785 7343 18788
rect 7285 18779 7343 18785
rect 7745 18785 7757 18788
rect 7791 18785 7803 18819
rect 7745 18779 7803 18785
rect 5868 18776 5874 18779
rect 2884 18720 3096 18748
rect 2884 18689 2912 18720
rect 4246 18708 4252 18760
rect 4304 18748 4310 18760
rect 4525 18751 4583 18757
rect 4525 18748 4537 18751
rect 4304 18720 4537 18748
rect 4304 18708 4310 18720
rect 4525 18717 4537 18720
rect 4571 18717 4583 18751
rect 4798 18748 4804 18760
rect 4525 18711 4583 18717
rect 4632 18720 4804 18748
rect 2869 18683 2927 18689
rect 2869 18649 2881 18683
rect 2915 18649 2927 18683
rect 2869 18643 2927 18649
rect 4341 18683 4399 18689
rect 4341 18649 4353 18683
rect 4387 18680 4399 18683
rect 4632 18680 4660 18720
rect 4798 18708 4804 18720
rect 4856 18748 4862 18760
rect 6012 18748 6040 18779
rect 8294 18776 8300 18828
rect 8352 18776 8358 18828
rect 8570 18776 8576 18828
rect 8628 18816 8634 18828
rect 8864 18825 8892 18856
rect 10134 18844 10140 18896
rect 10192 18884 10198 18896
rect 11149 18887 11207 18893
rect 10192 18856 10824 18884
rect 10192 18844 10198 18856
rect 8757 18819 8815 18825
rect 8757 18816 8769 18819
rect 8628 18788 8769 18816
rect 8628 18776 8634 18788
rect 8757 18785 8769 18788
rect 8803 18785 8815 18819
rect 8757 18779 8815 18785
rect 8849 18819 8907 18825
rect 8849 18785 8861 18819
rect 8895 18816 8907 18819
rect 8938 18816 8944 18828
rect 8895 18788 8944 18816
rect 8895 18785 8907 18788
rect 8849 18779 8907 18785
rect 8938 18776 8944 18788
rect 8996 18776 9002 18828
rect 9214 18776 9220 18828
rect 9272 18816 9278 18828
rect 9309 18819 9367 18825
rect 9309 18816 9321 18819
rect 9272 18788 9321 18816
rect 9272 18776 9278 18788
rect 9309 18785 9321 18788
rect 9355 18816 9367 18819
rect 9950 18816 9956 18828
rect 9355 18788 9956 18816
rect 9355 18785 9367 18788
rect 9309 18779 9367 18785
rect 9950 18776 9956 18788
rect 10008 18776 10014 18828
rect 10502 18776 10508 18828
rect 10560 18825 10566 18828
rect 10796 18825 10824 18856
rect 11149 18853 11161 18887
rect 11195 18884 11207 18887
rect 11609 18887 11667 18893
rect 11609 18884 11621 18887
rect 11195 18856 11621 18884
rect 11195 18853 11207 18856
rect 11149 18847 11207 18853
rect 11609 18853 11621 18856
rect 11655 18853 11667 18887
rect 12452 18884 12480 18924
rect 12526 18912 12532 18964
rect 12584 18952 12590 18964
rect 12621 18955 12679 18961
rect 12621 18952 12633 18955
rect 12584 18924 12633 18952
rect 12584 18912 12590 18924
rect 12621 18921 12633 18924
rect 12667 18921 12679 18955
rect 12621 18915 12679 18921
rect 12894 18912 12900 18964
rect 12952 18912 12958 18964
rect 13446 18912 13452 18964
rect 13504 18952 13510 18964
rect 13909 18955 13967 18961
rect 13909 18952 13921 18955
rect 13504 18924 13921 18952
rect 13504 18912 13510 18924
rect 13909 18921 13921 18924
rect 13955 18952 13967 18955
rect 13998 18952 14004 18964
rect 13955 18924 14004 18952
rect 13955 18921 13967 18924
rect 13909 18915 13967 18921
rect 13998 18912 14004 18924
rect 14056 18912 14062 18964
rect 14366 18912 14372 18964
rect 14424 18912 14430 18964
rect 15212 18924 15700 18952
rect 15212 18884 15240 18924
rect 12452 18856 15240 18884
rect 11609 18847 11667 18853
rect 15286 18844 15292 18896
rect 15344 18844 15350 18896
rect 10560 18779 10572 18825
rect 10781 18819 10839 18825
rect 10781 18785 10793 18819
rect 10827 18816 10839 18819
rect 10962 18816 10968 18828
rect 10827 18788 10968 18816
rect 10827 18785 10839 18788
rect 10781 18779 10839 18785
rect 10560 18776 10566 18779
rect 10962 18776 10968 18788
rect 11020 18776 11026 18828
rect 11054 18776 11060 18828
rect 11112 18816 11118 18828
rect 11793 18819 11851 18825
rect 11793 18816 11805 18819
rect 11112 18788 11805 18816
rect 11112 18776 11118 18788
rect 11793 18785 11805 18788
rect 11839 18785 11851 18819
rect 11793 18779 11851 18785
rect 11974 18776 11980 18828
rect 12032 18776 12038 18828
rect 12066 18776 12072 18828
rect 12124 18776 12130 18828
rect 12342 18776 12348 18828
rect 12400 18776 12406 18828
rect 12434 18776 12440 18828
rect 12492 18776 12498 18828
rect 12526 18776 12532 18828
rect 12584 18816 12590 18828
rect 13081 18819 13139 18825
rect 13081 18816 13093 18819
rect 12584 18788 13093 18816
rect 12584 18776 12590 18788
rect 13081 18785 13093 18788
rect 13127 18816 13139 18819
rect 13170 18816 13176 18828
rect 13127 18788 13176 18816
rect 13127 18785 13139 18788
rect 13081 18779 13139 18785
rect 13170 18776 13176 18788
rect 13228 18776 13234 18828
rect 13265 18819 13323 18825
rect 13265 18785 13277 18819
rect 13311 18816 13323 18819
rect 13446 18816 13452 18828
rect 13311 18788 13452 18816
rect 13311 18785 13323 18788
rect 13265 18779 13323 18785
rect 13446 18776 13452 18788
rect 13504 18776 13510 18828
rect 13541 18819 13599 18825
rect 13541 18785 13553 18819
rect 13587 18816 13599 18819
rect 13906 18816 13912 18828
rect 13587 18788 13912 18816
rect 13587 18785 13599 18788
rect 13541 18779 13599 18785
rect 13906 18776 13912 18788
rect 13964 18776 13970 18828
rect 14093 18819 14151 18825
rect 14093 18785 14105 18819
rect 14139 18785 14151 18819
rect 14093 18779 14151 18785
rect 14277 18819 14335 18825
rect 14277 18785 14289 18819
rect 14323 18816 14335 18819
rect 14366 18816 14372 18828
rect 14323 18788 14372 18816
rect 14323 18785 14335 18788
rect 14277 18779 14335 18785
rect 4856 18720 6040 18748
rect 4856 18708 4862 18720
rect 6454 18708 6460 18760
rect 6512 18748 6518 18760
rect 7009 18751 7067 18757
rect 7009 18748 7021 18751
rect 6512 18720 7021 18748
rect 6512 18708 6518 18720
rect 7009 18717 7021 18720
rect 7055 18717 7067 18751
rect 7009 18711 7067 18717
rect 7190 18708 7196 18760
rect 7248 18708 7254 18760
rect 9398 18708 9404 18760
rect 9456 18708 9462 18760
rect 11164 18720 12434 18748
rect 4387 18652 4660 18680
rect 4387 18649 4399 18652
rect 4341 18643 4399 18649
rect 5258 18640 5264 18692
rect 5316 18640 5322 18692
rect 5442 18640 5448 18692
rect 5500 18680 5506 18692
rect 8018 18680 8024 18692
rect 5500 18652 8024 18680
rect 5500 18640 5506 18652
rect 8018 18640 8024 18652
rect 8076 18680 8082 18692
rect 8665 18683 8723 18689
rect 8665 18680 8677 18683
rect 8076 18652 8677 18680
rect 8076 18640 8082 18652
rect 8665 18649 8677 18652
rect 8711 18649 8723 18683
rect 8665 18643 8723 18649
rect 9125 18683 9183 18689
rect 9125 18649 9137 18683
rect 9171 18680 9183 18683
rect 9416 18680 9444 18708
rect 9171 18652 9444 18680
rect 9171 18649 9183 18652
rect 9125 18643 9183 18649
rect 4890 18572 4896 18624
rect 4948 18572 4954 18624
rect 5537 18615 5595 18621
rect 5537 18581 5549 18615
rect 5583 18612 5595 18615
rect 5718 18612 5724 18624
rect 5583 18584 5724 18612
rect 5583 18581 5595 18584
rect 5537 18575 5595 18581
rect 5718 18572 5724 18584
rect 5776 18572 5782 18624
rect 5997 18615 6055 18621
rect 5997 18581 6009 18615
rect 6043 18612 6055 18615
rect 6086 18612 6092 18624
rect 6043 18584 6092 18612
rect 6043 18581 6055 18584
rect 5997 18575 6055 18581
rect 6086 18572 6092 18584
rect 6144 18572 6150 18624
rect 6178 18572 6184 18624
rect 6236 18612 6242 18624
rect 8570 18612 8576 18624
rect 6236 18584 8576 18612
rect 6236 18572 6242 18584
rect 8570 18572 8576 18584
rect 8628 18572 8634 18624
rect 9033 18615 9091 18621
rect 9033 18581 9045 18615
rect 9079 18612 9091 18615
rect 9306 18612 9312 18624
rect 9079 18584 9312 18612
rect 9079 18581 9091 18584
rect 9033 18575 9091 18581
rect 9306 18572 9312 18584
rect 9364 18572 9370 18624
rect 9398 18572 9404 18624
rect 9456 18572 9462 18624
rect 10410 18572 10416 18624
rect 10468 18612 10474 18624
rect 11164 18621 11192 18720
rect 11514 18640 11520 18692
rect 11572 18640 11578 18692
rect 11790 18640 11796 18692
rect 11848 18680 11854 18692
rect 12066 18680 12072 18692
rect 11848 18652 12072 18680
rect 11848 18640 11854 18652
rect 12066 18640 12072 18652
rect 12124 18680 12130 18692
rect 12161 18683 12219 18689
rect 12161 18680 12173 18683
rect 12124 18652 12173 18680
rect 12124 18640 12130 18652
rect 12161 18649 12173 18652
rect 12207 18649 12219 18683
rect 12161 18643 12219 18649
rect 10965 18615 11023 18621
rect 10965 18612 10977 18615
rect 10468 18584 10977 18612
rect 10468 18572 10474 18584
rect 10965 18581 10977 18584
rect 11011 18581 11023 18615
rect 10965 18575 11023 18581
rect 11149 18615 11207 18621
rect 11149 18581 11161 18615
rect 11195 18581 11207 18615
rect 12406 18612 12434 18720
rect 13814 18708 13820 18760
rect 13872 18748 13878 18760
rect 14108 18748 14136 18779
rect 14366 18776 14372 18788
rect 14424 18816 14430 18828
rect 14553 18819 14611 18825
rect 14553 18816 14565 18819
rect 14424 18788 14565 18816
rect 14424 18776 14430 18788
rect 14553 18785 14565 18788
rect 14599 18785 14611 18819
rect 14553 18779 14611 18785
rect 14737 18819 14795 18825
rect 14737 18785 14749 18819
rect 14783 18816 14795 18819
rect 15565 18819 15623 18825
rect 15565 18816 15577 18819
rect 14783 18788 14964 18816
rect 14783 18785 14795 18788
rect 14737 18779 14795 18785
rect 14936 18748 14964 18788
rect 13872 18720 14964 18748
rect 13872 18708 13878 18720
rect 14936 18689 14964 18720
rect 15488 18788 15577 18816
rect 15488 18689 15516 18788
rect 15565 18785 15577 18788
rect 15611 18785 15623 18819
rect 15565 18779 15623 18785
rect 14921 18683 14979 18689
rect 12820 18652 14044 18680
rect 12820 18624 12848 18652
rect 12802 18612 12808 18624
rect 12406 18584 12808 18612
rect 11149 18575 11207 18581
rect 12802 18572 12808 18584
rect 12860 18572 12866 18624
rect 13170 18572 13176 18624
rect 13228 18612 13234 18624
rect 13357 18615 13415 18621
rect 13357 18612 13369 18615
rect 13228 18584 13369 18612
rect 13228 18572 13234 18584
rect 13357 18581 13369 18584
rect 13403 18581 13415 18615
rect 14016 18612 14044 18652
rect 14921 18649 14933 18683
rect 14967 18680 14979 18683
rect 15473 18683 15531 18689
rect 14967 18652 15424 18680
rect 14967 18649 14979 18652
rect 14921 18643 14979 18649
rect 15289 18615 15347 18621
rect 15289 18612 15301 18615
rect 14016 18584 15301 18612
rect 13357 18575 13415 18581
rect 15289 18581 15301 18584
rect 15335 18581 15347 18615
rect 15396 18612 15424 18652
rect 15473 18649 15485 18683
rect 15519 18649 15531 18683
rect 15672 18680 15700 18924
rect 15746 18912 15752 18964
rect 15804 18912 15810 18964
rect 16850 18912 16856 18964
rect 16908 18912 16914 18964
rect 17034 18912 17040 18964
rect 17092 18912 17098 18964
rect 17497 18955 17555 18961
rect 17497 18921 17509 18955
rect 17543 18952 17555 18955
rect 17770 18952 17776 18964
rect 17543 18924 17776 18952
rect 17543 18921 17555 18924
rect 17497 18915 17555 18921
rect 17770 18912 17776 18924
rect 17828 18912 17834 18964
rect 17954 18912 17960 18964
rect 18012 18912 18018 18964
rect 18141 18955 18199 18961
rect 18141 18921 18153 18955
rect 18187 18921 18199 18955
rect 18141 18915 18199 18921
rect 18417 18955 18475 18961
rect 18417 18921 18429 18955
rect 18463 18952 18475 18955
rect 18966 18952 18972 18964
rect 18463 18924 18972 18952
rect 18463 18921 18475 18924
rect 18417 18915 18475 18921
rect 16868 18884 16896 18912
rect 16776 18856 16896 18884
rect 16776 18825 16804 18856
rect 16761 18819 16819 18825
rect 16761 18785 16773 18819
rect 16807 18785 16819 18819
rect 16761 18779 16819 18785
rect 16853 18819 16911 18825
rect 16853 18785 16865 18819
rect 16899 18816 16911 18819
rect 16942 18816 16948 18828
rect 16899 18788 16948 18816
rect 16899 18785 16911 18788
rect 16853 18779 16911 18785
rect 16942 18776 16948 18788
rect 17000 18776 17006 18828
rect 17310 18776 17316 18828
rect 17368 18776 17374 18828
rect 17586 18776 17592 18828
rect 17644 18776 17650 18828
rect 18156 18816 18184 18915
rect 18966 18912 18972 18924
rect 19024 18912 19030 18964
rect 20438 18952 20444 18964
rect 19076 18924 20444 18952
rect 18322 18844 18328 18896
rect 18380 18884 18386 18896
rect 19076 18884 19104 18924
rect 20438 18912 20444 18924
rect 20496 18912 20502 18964
rect 20898 18912 20904 18964
rect 20956 18952 20962 18964
rect 21637 18955 21695 18961
rect 21637 18952 21649 18955
rect 20956 18924 21649 18952
rect 20956 18912 20962 18924
rect 21637 18921 21649 18924
rect 21683 18921 21695 18955
rect 21637 18915 21695 18921
rect 21726 18912 21732 18964
rect 21784 18952 21790 18964
rect 22278 18952 22284 18964
rect 21784 18924 22284 18952
rect 21784 18912 21790 18924
rect 22278 18912 22284 18924
rect 22336 18952 22342 18964
rect 22922 18952 22928 18964
rect 22336 18924 22928 18952
rect 22336 18912 22342 18924
rect 22922 18912 22928 18924
rect 22980 18912 22986 18964
rect 18380 18856 19104 18884
rect 18380 18844 18386 18856
rect 19242 18844 19248 18896
rect 19300 18884 19306 18896
rect 19300 18856 21036 18884
rect 19300 18844 19306 18856
rect 18233 18819 18291 18825
rect 18233 18816 18245 18819
rect 18156 18788 18245 18816
rect 18233 18785 18245 18788
rect 18279 18785 18291 18819
rect 19426 18816 19432 18828
rect 18233 18779 18291 18785
rect 18892 18788 19432 18816
rect 15930 18708 15936 18760
rect 15988 18748 15994 18760
rect 18892 18748 18920 18788
rect 19426 18776 19432 18788
rect 19484 18776 19490 18828
rect 15988 18720 18920 18748
rect 15988 18708 15994 18720
rect 18966 18708 18972 18760
rect 19024 18748 19030 18760
rect 19628 18757 19656 18856
rect 19886 18776 19892 18828
rect 19944 18776 19950 18828
rect 20530 18776 20536 18828
rect 20588 18776 20594 18828
rect 21008 18816 21036 18856
rect 21082 18844 21088 18896
rect 21140 18884 21146 18896
rect 22094 18884 22100 18896
rect 21140 18856 22100 18884
rect 21140 18844 21146 18856
rect 22094 18844 22100 18856
rect 22152 18844 22158 18896
rect 21174 18816 21180 18828
rect 21008 18788 21180 18816
rect 21174 18776 21180 18788
rect 21232 18776 21238 18828
rect 21453 18819 21511 18825
rect 21453 18785 21465 18819
rect 21499 18785 21511 18819
rect 21453 18779 21511 18785
rect 22761 18819 22819 18825
rect 22761 18785 22773 18819
rect 22807 18816 22819 18819
rect 22922 18816 22928 18828
rect 22807 18788 22928 18816
rect 22807 18785 22819 18788
rect 22761 18779 22819 18785
rect 19153 18751 19211 18757
rect 19153 18748 19165 18751
rect 19024 18720 19165 18748
rect 19024 18708 19030 18720
rect 19153 18717 19165 18720
rect 19199 18717 19211 18751
rect 19153 18711 19211 18717
rect 19613 18751 19671 18757
rect 19613 18717 19625 18751
rect 19659 18717 19671 18751
rect 19613 18711 19671 18717
rect 19797 18751 19855 18757
rect 19797 18717 19809 18751
rect 19843 18748 19855 18751
rect 20162 18748 20168 18760
rect 19843 18720 20168 18748
rect 19843 18717 19855 18720
rect 19797 18711 19855 18717
rect 20162 18708 20168 18720
rect 20220 18708 20226 18760
rect 20438 18708 20444 18760
rect 20496 18708 20502 18760
rect 20901 18751 20959 18757
rect 20901 18717 20913 18751
rect 20947 18748 20959 18751
rect 20990 18748 20996 18760
rect 20947 18720 20996 18748
rect 20947 18717 20959 18720
rect 20901 18711 20959 18717
rect 20990 18708 20996 18720
rect 21048 18708 21054 18760
rect 20070 18680 20076 18692
rect 15672 18652 20076 18680
rect 15473 18643 15531 18649
rect 20070 18640 20076 18652
rect 20128 18640 20134 18692
rect 20257 18683 20315 18689
rect 20257 18649 20269 18683
rect 20303 18680 20315 18683
rect 21468 18680 21496 18779
rect 22922 18776 22928 18788
rect 22980 18776 22986 18828
rect 23017 18751 23075 18757
rect 23017 18717 23029 18751
rect 23063 18717 23075 18751
rect 23017 18711 23075 18717
rect 20303 18652 21496 18680
rect 20303 18649 20315 18652
rect 20257 18643 20315 18649
rect 16942 18612 16948 18624
rect 15396 18584 16948 18612
rect 15289 18575 15347 18581
rect 16942 18572 16948 18584
rect 17000 18572 17006 18624
rect 17586 18572 17592 18624
rect 17644 18612 17650 18624
rect 17862 18612 17868 18624
rect 17644 18584 17868 18612
rect 17644 18572 17650 18584
rect 17862 18572 17868 18584
rect 17920 18612 17926 18624
rect 17957 18615 18015 18621
rect 17957 18612 17969 18615
rect 17920 18584 17969 18612
rect 17920 18572 17926 18584
rect 17957 18581 17969 18584
rect 18003 18581 18015 18615
rect 17957 18575 18015 18581
rect 19978 18572 19984 18624
rect 20036 18612 20042 18624
rect 21269 18615 21327 18621
rect 21269 18612 21281 18615
rect 20036 18584 21281 18612
rect 20036 18572 20042 18584
rect 21269 18581 21281 18584
rect 21315 18581 21327 18615
rect 21269 18575 21327 18581
rect 21726 18572 21732 18624
rect 21784 18612 21790 18624
rect 23032 18612 23060 18711
rect 21784 18584 23060 18612
rect 21784 18572 21790 18584
rect 552 18522 23368 18544
rect 552 18470 1366 18522
rect 1418 18470 1430 18522
rect 1482 18470 1494 18522
rect 1546 18470 1558 18522
rect 1610 18470 1622 18522
rect 1674 18470 1686 18522
rect 1738 18470 7366 18522
rect 7418 18470 7430 18522
rect 7482 18470 7494 18522
rect 7546 18470 7558 18522
rect 7610 18470 7622 18522
rect 7674 18470 7686 18522
rect 7738 18470 13366 18522
rect 13418 18470 13430 18522
rect 13482 18470 13494 18522
rect 13546 18470 13558 18522
rect 13610 18470 13622 18522
rect 13674 18470 13686 18522
rect 13738 18470 19366 18522
rect 19418 18470 19430 18522
rect 19482 18470 19494 18522
rect 19546 18470 19558 18522
rect 19610 18470 19622 18522
rect 19674 18470 19686 18522
rect 19738 18470 23368 18522
rect 552 18448 23368 18470
rect 2314 18368 2320 18420
rect 2372 18408 2378 18420
rect 3970 18408 3976 18420
rect 2372 18380 3976 18408
rect 2372 18368 2378 18380
rect 3970 18368 3976 18380
rect 4028 18408 4034 18420
rect 4249 18411 4307 18417
rect 4249 18408 4261 18411
rect 4028 18380 4261 18408
rect 4028 18368 4034 18380
rect 4249 18377 4261 18380
rect 4295 18377 4307 18411
rect 4249 18371 4307 18377
rect 6454 18368 6460 18420
rect 6512 18368 6518 18420
rect 6917 18411 6975 18417
rect 6917 18377 6929 18411
rect 6963 18408 6975 18411
rect 6963 18380 7236 18408
rect 6963 18377 6975 18380
rect 6917 18371 6975 18377
rect 1949 18343 2007 18349
rect 1949 18309 1961 18343
rect 1995 18340 2007 18343
rect 2038 18340 2044 18352
rect 1995 18312 2044 18340
rect 1995 18309 2007 18312
rect 1949 18303 2007 18309
rect 2038 18300 2044 18312
rect 2096 18300 2102 18352
rect 4890 18300 4896 18352
rect 4948 18340 4954 18352
rect 5810 18340 5816 18352
rect 4948 18312 5816 18340
rect 4948 18300 4954 18312
rect 5810 18300 5816 18312
rect 5868 18300 5874 18352
rect 5902 18300 5908 18352
rect 5960 18300 5966 18352
rect 7208 18340 7236 18380
rect 7282 18368 7288 18420
rect 7340 18408 7346 18420
rect 7745 18411 7803 18417
rect 7745 18408 7757 18411
rect 7340 18380 7757 18408
rect 7340 18368 7346 18380
rect 7745 18377 7757 18380
rect 7791 18377 7803 18411
rect 7745 18371 7803 18377
rect 8113 18411 8171 18417
rect 8113 18377 8125 18411
rect 8159 18408 8171 18411
rect 8754 18408 8760 18420
rect 8159 18380 8760 18408
rect 8159 18377 8171 18380
rect 8113 18371 8171 18377
rect 8754 18368 8760 18380
rect 8812 18368 8818 18420
rect 10413 18411 10471 18417
rect 9048 18380 9812 18408
rect 6656 18312 7144 18340
rect 7208 18312 7972 18340
rect 1765 18275 1823 18281
rect 1765 18241 1777 18275
rect 1811 18241 1823 18275
rect 2958 18272 2964 18284
rect 1765 18235 1823 18241
rect 2056 18244 2964 18272
rect 1780 18136 1808 18235
rect 1946 18164 1952 18216
rect 2004 18204 2010 18216
rect 2056 18213 2084 18244
rect 2958 18232 2964 18244
rect 3016 18232 3022 18284
rect 4154 18232 4160 18284
rect 4212 18272 4218 18284
rect 4341 18275 4399 18281
rect 4341 18272 4353 18275
rect 4212 18244 4353 18272
rect 4212 18232 4218 18244
rect 4341 18241 4353 18244
rect 4387 18241 4399 18275
rect 5166 18272 5172 18284
rect 4341 18235 4399 18241
rect 4540 18244 5172 18272
rect 2041 18207 2099 18213
rect 2041 18204 2053 18207
rect 2004 18176 2053 18204
rect 2004 18164 2010 18176
rect 2041 18173 2053 18176
rect 2087 18173 2099 18207
rect 2041 18167 2099 18173
rect 2774 18164 2780 18216
rect 2832 18204 2838 18216
rect 2869 18207 2927 18213
rect 2869 18204 2881 18207
rect 2832 18176 2881 18204
rect 2832 18164 2838 18176
rect 2869 18173 2881 18176
rect 2915 18173 2927 18207
rect 2869 18167 2927 18173
rect 3053 18207 3111 18213
rect 3053 18173 3065 18207
rect 3099 18173 3111 18207
rect 3053 18167 3111 18173
rect 3973 18207 4031 18213
rect 3973 18173 3985 18207
rect 4019 18204 4031 18207
rect 4062 18204 4068 18216
rect 4019 18176 4068 18204
rect 4019 18173 4031 18176
rect 3973 18167 4031 18173
rect 2222 18136 2228 18148
rect 1780 18108 2228 18136
rect 2222 18096 2228 18108
rect 2280 18096 2286 18148
rect 2682 18096 2688 18148
rect 2740 18136 2746 18148
rect 3068 18136 3096 18167
rect 4062 18164 4068 18176
rect 4120 18164 4126 18216
rect 4540 18213 4568 18244
rect 5166 18232 5172 18244
rect 5224 18232 5230 18284
rect 5258 18232 5264 18284
rect 5316 18272 5322 18284
rect 5316 18244 6224 18272
rect 5316 18232 5322 18244
rect 6196 18216 6224 18244
rect 4525 18207 4583 18213
rect 4525 18173 4537 18207
rect 4571 18173 4583 18207
rect 4525 18167 4583 18173
rect 5077 18207 5135 18213
rect 5077 18173 5089 18207
rect 5123 18173 5135 18207
rect 5077 18167 5135 18173
rect 5353 18207 5411 18213
rect 5353 18173 5365 18207
rect 5399 18173 5411 18207
rect 5353 18167 5411 18173
rect 5629 18207 5687 18213
rect 5629 18173 5641 18207
rect 5675 18204 5687 18207
rect 6086 18204 6092 18216
rect 5675 18176 6092 18204
rect 5675 18173 5687 18176
rect 5629 18167 5687 18173
rect 2740 18108 3096 18136
rect 2740 18096 2746 18108
rect 4246 18096 4252 18148
rect 4304 18136 4310 18148
rect 5092 18136 5120 18167
rect 5261 18139 5319 18145
rect 5261 18136 5273 18139
rect 4304 18108 5273 18136
rect 4304 18096 4310 18108
rect 5261 18105 5273 18108
rect 5307 18105 5319 18139
rect 5261 18099 5319 18105
rect 1762 18028 1768 18080
rect 1820 18028 1826 18080
rect 2961 18071 3019 18077
rect 2961 18037 2973 18071
rect 3007 18068 3019 18071
rect 3050 18068 3056 18080
rect 3007 18040 3056 18068
rect 3007 18037 3019 18040
rect 2961 18031 3019 18037
rect 3050 18028 3056 18040
rect 3108 18028 3114 18080
rect 3878 18028 3884 18080
rect 3936 18068 3942 18080
rect 4157 18071 4215 18077
rect 4157 18068 4169 18071
rect 3936 18040 4169 18068
rect 3936 18028 3942 18040
rect 4157 18037 4169 18040
rect 4203 18037 4215 18071
rect 4157 18031 4215 18037
rect 4709 18071 4767 18077
rect 4709 18037 4721 18071
rect 4755 18068 4767 18071
rect 4798 18068 4804 18080
rect 4755 18040 4804 18068
rect 4755 18037 4767 18040
rect 4709 18031 4767 18037
rect 4798 18028 4804 18040
rect 4856 18028 4862 18080
rect 4890 18028 4896 18080
rect 4948 18028 4954 18080
rect 4982 18028 4988 18080
rect 5040 18068 5046 18080
rect 5368 18068 5396 18167
rect 6086 18164 6092 18176
rect 6144 18164 6150 18216
rect 6178 18164 6184 18216
rect 6236 18164 6242 18216
rect 6656 18213 6684 18312
rect 7116 18281 7144 18312
rect 7101 18275 7159 18281
rect 7101 18241 7113 18275
rect 7147 18272 7159 18275
rect 7147 18244 7788 18272
rect 7147 18241 7159 18244
rect 7101 18235 7159 18241
rect 6641 18207 6699 18213
rect 6641 18173 6653 18207
rect 6687 18173 6699 18207
rect 6641 18167 6699 18173
rect 6733 18207 6791 18213
rect 6733 18173 6745 18207
rect 6779 18204 6791 18207
rect 6914 18204 6920 18216
rect 6779 18176 6920 18204
rect 6779 18173 6791 18176
rect 6733 18167 6791 18173
rect 6914 18164 6920 18176
rect 6972 18164 6978 18216
rect 7009 18207 7067 18213
rect 7009 18173 7021 18207
rect 7055 18204 7067 18207
rect 7190 18204 7196 18216
rect 7055 18176 7196 18204
rect 7055 18173 7067 18176
rect 7009 18167 7067 18173
rect 7190 18164 7196 18176
rect 7248 18164 7254 18216
rect 7285 18207 7343 18213
rect 7285 18173 7297 18207
rect 7331 18173 7343 18207
rect 7285 18167 7343 18173
rect 5905 18139 5963 18145
rect 5905 18105 5917 18139
rect 5951 18136 5963 18139
rect 6362 18136 6368 18148
rect 5951 18108 6368 18136
rect 5951 18105 5963 18108
rect 5905 18099 5963 18105
rect 6362 18096 6368 18108
rect 6420 18096 6426 18148
rect 6822 18096 6828 18148
rect 6880 18136 6886 18148
rect 7300 18136 7328 18167
rect 7374 18164 7380 18216
rect 7432 18164 7438 18216
rect 7466 18164 7472 18216
rect 7524 18164 7530 18216
rect 7561 18207 7619 18213
rect 7561 18173 7573 18207
rect 7607 18204 7619 18207
rect 7650 18204 7656 18216
rect 7607 18176 7656 18204
rect 7607 18173 7619 18176
rect 7561 18167 7619 18173
rect 7650 18164 7656 18176
rect 7708 18164 7714 18216
rect 7760 18213 7788 18244
rect 7944 18216 7972 18312
rect 8386 18300 8392 18352
rect 8444 18340 8450 18352
rect 8481 18343 8539 18349
rect 8481 18340 8493 18343
rect 8444 18312 8493 18340
rect 8444 18300 8450 18312
rect 8481 18309 8493 18312
rect 8527 18309 8539 18343
rect 8481 18303 8539 18309
rect 7745 18207 7803 18213
rect 7745 18173 7757 18207
rect 7791 18173 7803 18207
rect 7745 18167 7803 18173
rect 7926 18164 7932 18216
rect 7984 18164 7990 18216
rect 8018 18164 8024 18216
rect 8076 18164 8082 18216
rect 8849 18207 8907 18213
rect 8849 18173 8861 18207
rect 8895 18204 8907 18207
rect 8941 18207 8999 18213
rect 8941 18204 8953 18207
rect 8895 18176 8953 18204
rect 8895 18173 8907 18176
rect 8849 18167 8907 18173
rect 8941 18173 8953 18176
rect 8987 18204 8999 18207
rect 9048 18204 9076 18380
rect 9585 18343 9643 18349
rect 9585 18309 9597 18343
rect 9631 18340 9643 18343
rect 9674 18340 9680 18352
rect 9631 18312 9680 18340
rect 9631 18309 9643 18312
rect 9585 18303 9643 18309
rect 9674 18300 9680 18312
rect 9732 18300 9738 18352
rect 9784 18340 9812 18380
rect 10413 18377 10425 18411
rect 10459 18408 10471 18411
rect 10502 18408 10508 18420
rect 10459 18380 10508 18408
rect 10459 18377 10471 18380
rect 10413 18371 10471 18377
rect 10502 18368 10508 18380
rect 10560 18368 10566 18420
rect 11149 18411 11207 18417
rect 11149 18377 11161 18411
rect 11195 18408 11207 18411
rect 11698 18408 11704 18420
rect 11195 18380 11704 18408
rect 11195 18377 11207 18380
rect 11149 18371 11207 18377
rect 11698 18368 11704 18380
rect 11756 18368 11762 18420
rect 12342 18408 12348 18420
rect 11808 18380 12348 18408
rect 11422 18340 11428 18352
rect 9784 18312 11428 18340
rect 11422 18300 11428 18312
rect 11480 18300 11486 18352
rect 11330 18272 11336 18284
rect 9140 18244 9720 18272
rect 9140 18213 9168 18244
rect 8987 18176 9076 18204
rect 9125 18207 9183 18213
rect 8987 18173 8999 18176
rect 8941 18167 8999 18173
rect 9125 18173 9137 18207
rect 9171 18173 9183 18207
rect 9125 18167 9183 18173
rect 9309 18207 9367 18213
rect 9309 18173 9321 18207
rect 9355 18204 9367 18207
rect 9490 18204 9496 18216
rect 9355 18176 9496 18204
rect 9355 18173 9367 18176
rect 9309 18167 9367 18173
rect 9490 18164 9496 18176
rect 9548 18164 9554 18216
rect 9692 18213 9720 18244
rect 9876 18244 11336 18272
rect 9876 18213 9904 18244
rect 11330 18232 11336 18244
rect 11388 18232 11394 18284
rect 9677 18207 9735 18213
rect 9677 18173 9689 18207
rect 9723 18173 9735 18207
rect 9677 18167 9735 18173
rect 9861 18207 9919 18213
rect 9861 18173 9873 18207
rect 9907 18173 9919 18207
rect 9861 18167 9919 18173
rect 10229 18207 10287 18213
rect 10229 18173 10241 18207
rect 10275 18204 10287 18207
rect 10410 18204 10416 18216
rect 10275 18176 10416 18204
rect 10275 18173 10287 18176
rect 10229 18167 10287 18173
rect 8754 18136 8760 18148
rect 6880 18108 7328 18136
rect 7944 18108 8760 18136
rect 6880 18096 6886 18108
rect 5040 18040 5396 18068
rect 5040 18028 5046 18040
rect 5718 18028 5724 18080
rect 5776 18028 5782 18080
rect 5810 18028 5816 18080
rect 5868 18068 5874 18080
rect 5997 18071 6055 18077
rect 5997 18068 6009 18071
rect 5868 18040 6009 18068
rect 5868 18028 5874 18040
rect 5997 18037 6009 18040
rect 6043 18037 6055 18071
rect 5997 18031 6055 18037
rect 6270 18028 6276 18080
rect 6328 18068 6334 18080
rect 6914 18068 6920 18080
rect 6328 18040 6920 18068
rect 6328 18028 6334 18040
rect 6914 18028 6920 18040
rect 6972 18028 6978 18080
rect 7190 18028 7196 18080
rect 7248 18068 7254 18080
rect 7944 18068 7972 18108
rect 8754 18096 8760 18108
rect 8812 18096 8818 18148
rect 9582 18096 9588 18148
rect 9640 18096 9646 18148
rect 9692 18136 9720 18167
rect 10410 18164 10416 18176
rect 10468 18164 10474 18216
rect 11698 18164 11704 18216
rect 11756 18164 11762 18216
rect 10134 18136 10140 18148
rect 9692 18108 10140 18136
rect 10134 18096 10140 18108
rect 10192 18096 10198 18148
rect 10965 18139 11023 18145
rect 10965 18105 10977 18139
rect 11011 18136 11023 18139
rect 11054 18136 11060 18148
rect 11011 18108 11060 18136
rect 11011 18105 11023 18108
rect 10965 18099 11023 18105
rect 11054 18096 11060 18108
rect 11112 18096 11118 18148
rect 11181 18139 11239 18145
rect 11181 18105 11193 18139
rect 11227 18136 11239 18139
rect 11808 18136 11836 18380
rect 12342 18368 12348 18380
rect 12400 18408 12406 18420
rect 13541 18411 13599 18417
rect 13541 18408 13553 18411
rect 12400 18380 13553 18408
rect 12400 18368 12406 18380
rect 13541 18377 13553 18380
rect 13587 18377 13599 18411
rect 13541 18371 13599 18377
rect 13725 18411 13783 18417
rect 13725 18377 13737 18411
rect 13771 18408 13783 18411
rect 14182 18408 14188 18420
rect 13771 18380 14188 18408
rect 13771 18377 13783 18380
rect 13725 18371 13783 18377
rect 14182 18368 14188 18380
rect 14240 18368 14246 18420
rect 14660 18380 15240 18408
rect 13357 18343 13415 18349
rect 13357 18309 13369 18343
rect 13403 18340 13415 18343
rect 14660 18340 14688 18380
rect 13403 18312 14688 18340
rect 13403 18309 13415 18312
rect 13357 18303 13415 18309
rect 14734 18300 14740 18352
rect 14792 18340 14798 18352
rect 14921 18343 14979 18349
rect 14921 18340 14933 18343
rect 14792 18312 14933 18340
rect 14792 18300 14798 18312
rect 14921 18309 14933 18312
rect 14967 18309 14979 18343
rect 15212 18340 15240 18380
rect 15286 18368 15292 18420
rect 15344 18408 15350 18420
rect 16761 18411 16819 18417
rect 16761 18408 16773 18411
rect 15344 18380 16773 18408
rect 15344 18368 15350 18380
rect 16761 18377 16773 18380
rect 16807 18377 16819 18411
rect 16761 18371 16819 18377
rect 17586 18368 17592 18420
rect 17644 18408 17650 18420
rect 18049 18411 18107 18417
rect 18049 18408 18061 18411
rect 17644 18380 18061 18408
rect 17644 18368 17650 18380
rect 18049 18377 18061 18380
rect 18095 18377 18107 18411
rect 18049 18371 18107 18377
rect 18156 18380 18368 18408
rect 15212 18312 18092 18340
rect 14921 18303 14979 18309
rect 16114 18272 16120 18284
rect 14108 18244 16120 18272
rect 11977 18207 12035 18213
rect 11977 18173 11989 18207
rect 12023 18204 12035 18207
rect 14108 18204 14136 18244
rect 16114 18232 16120 18244
rect 16172 18232 16178 18284
rect 16224 18281 16252 18312
rect 18064 18284 18092 18312
rect 16209 18275 16267 18281
rect 16209 18241 16221 18275
rect 16255 18241 16267 18275
rect 16209 18235 16267 18241
rect 16669 18275 16727 18281
rect 16669 18241 16681 18275
rect 16715 18272 16727 18275
rect 16850 18272 16856 18284
rect 16715 18244 16856 18272
rect 16715 18241 16727 18244
rect 16669 18235 16727 18241
rect 16850 18232 16856 18244
rect 16908 18232 16914 18284
rect 17221 18275 17279 18281
rect 17221 18272 17233 18275
rect 17144 18244 17233 18272
rect 12023 18176 14136 18204
rect 12023 18173 12035 18176
rect 11977 18167 12035 18173
rect 14182 18164 14188 18216
rect 14240 18164 14246 18216
rect 14829 18207 14887 18213
rect 14829 18173 14841 18207
rect 14875 18204 14887 18207
rect 15102 18204 15108 18216
rect 14875 18176 15108 18204
rect 14875 18173 14887 18176
rect 14829 18167 14887 18173
rect 15102 18164 15108 18176
rect 15160 18164 15166 18216
rect 15562 18164 15568 18216
rect 15620 18204 15626 18216
rect 16301 18207 16359 18213
rect 16301 18204 16313 18207
rect 15620 18176 16313 18204
rect 15620 18164 15626 18176
rect 16301 18173 16313 18176
rect 16347 18204 16359 18207
rect 17034 18204 17040 18216
rect 16347 18176 17040 18204
rect 16347 18173 16359 18176
rect 16301 18167 16359 18173
rect 17034 18164 17040 18176
rect 17092 18164 17098 18216
rect 17144 18213 17172 18244
rect 17221 18241 17233 18244
rect 17267 18272 17279 18275
rect 17681 18275 17739 18281
rect 17681 18272 17693 18275
rect 17267 18244 17693 18272
rect 17267 18241 17279 18244
rect 17221 18235 17279 18241
rect 17681 18241 17693 18244
rect 17727 18241 17739 18275
rect 17681 18235 17739 18241
rect 18046 18232 18052 18284
rect 18104 18232 18110 18284
rect 17129 18207 17187 18213
rect 17129 18173 17141 18207
rect 17175 18173 17187 18207
rect 17129 18167 17187 18173
rect 17405 18207 17463 18213
rect 17405 18173 17417 18207
rect 17451 18204 17463 18207
rect 17494 18204 17500 18216
rect 17451 18176 17500 18204
rect 17451 18173 17463 18176
rect 17405 18167 17463 18173
rect 17494 18164 17500 18176
rect 17552 18164 17558 18216
rect 17589 18207 17647 18213
rect 17589 18173 17601 18207
rect 17635 18204 17647 18207
rect 18156 18204 18184 18380
rect 18340 18349 18368 18380
rect 18414 18368 18420 18420
rect 18472 18408 18478 18420
rect 18472 18380 20392 18408
rect 18472 18368 18478 18380
rect 18233 18343 18291 18349
rect 18233 18309 18245 18343
rect 18279 18309 18291 18343
rect 18233 18303 18291 18309
rect 18325 18343 18383 18349
rect 18325 18309 18337 18343
rect 18371 18340 18383 18343
rect 18874 18340 18880 18352
rect 18371 18312 18880 18340
rect 18371 18309 18383 18312
rect 18325 18303 18383 18309
rect 18248 18272 18276 18303
rect 18874 18300 18880 18312
rect 18932 18300 18938 18352
rect 20364 18340 20392 18380
rect 21082 18368 21088 18420
rect 21140 18368 21146 18420
rect 21192 18380 23060 18408
rect 21192 18340 21220 18380
rect 20364 18312 21220 18340
rect 21358 18300 21364 18352
rect 21416 18340 21422 18352
rect 22281 18343 22339 18349
rect 22281 18340 22293 18343
rect 21416 18312 22293 18340
rect 21416 18300 21422 18312
rect 22281 18309 22293 18312
rect 22327 18309 22339 18343
rect 22833 18343 22891 18349
rect 22833 18340 22845 18343
rect 22281 18303 22339 18309
rect 22388 18312 22845 18340
rect 18248 18244 18736 18272
rect 17635 18176 18184 18204
rect 17635 18173 17647 18176
rect 17589 18167 17647 18173
rect 18506 18164 18512 18216
rect 18564 18164 18570 18216
rect 18708 18204 18736 18244
rect 18782 18232 18788 18284
rect 18840 18272 18846 18284
rect 19429 18275 19487 18281
rect 19429 18272 19441 18275
rect 18840 18244 19441 18272
rect 18840 18232 18846 18244
rect 19429 18241 19441 18244
rect 19475 18241 19487 18275
rect 21269 18275 21327 18281
rect 21269 18272 21281 18275
rect 19429 18235 19487 18241
rect 20456 18244 21281 18272
rect 19337 18207 19395 18213
rect 19337 18204 19349 18207
rect 18708 18176 19349 18204
rect 19337 18173 19349 18176
rect 19383 18173 19395 18207
rect 19337 18167 19395 18173
rect 19696 18207 19754 18213
rect 19696 18173 19708 18207
rect 19742 18204 19754 18207
rect 19978 18204 19984 18216
rect 19742 18176 19984 18204
rect 19742 18173 19754 18176
rect 19696 18167 19754 18173
rect 19978 18164 19984 18176
rect 20036 18164 20042 18216
rect 20070 18164 20076 18216
rect 20128 18204 20134 18216
rect 20456 18204 20484 18244
rect 21269 18241 21281 18244
rect 21315 18241 21327 18275
rect 21269 18235 21327 18241
rect 21450 18232 21456 18284
rect 21508 18272 21514 18284
rect 22388 18272 22416 18312
rect 22833 18309 22845 18312
rect 22879 18309 22891 18343
rect 22833 18303 22891 18309
rect 21508 18244 22416 18272
rect 22465 18275 22523 18281
rect 21508 18232 21514 18244
rect 22465 18241 22477 18275
rect 22511 18241 22523 18275
rect 22465 18235 22523 18241
rect 20128 18176 20484 18204
rect 20901 18207 20959 18213
rect 20128 18164 20134 18176
rect 20901 18173 20913 18207
rect 20947 18204 20959 18207
rect 22005 18207 22063 18213
rect 22005 18204 22017 18207
rect 20947 18176 22017 18204
rect 20947 18173 20959 18176
rect 20901 18167 20959 18173
rect 12222 18139 12280 18145
rect 12222 18136 12234 18139
rect 11227 18108 11836 18136
rect 11900 18108 12234 18136
rect 11227 18105 11239 18108
rect 11181 18099 11239 18105
rect 7248 18040 7972 18068
rect 7248 18028 7254 18040
rect 8018 18028 8024 18080
rect 8076 18068 8082 18080
rect 8389 18071 8447 18077
rect 8389 18068 8401 18071
rect 8076 18040 8401 18068
rect 8076 18028 8082 18040
rect 8389 18037 8401 18040
rect 8435 18037 8447 18071
rect 8389 18031 8447 18037
rect 8938 18028 8944 18080
rect 8996 18068 9002 18080
rect 9033 18071 9091 18077
rect 9033 18068 9045 18071
rect 8996 18040 9045 18068
rect 8996 18028 9002 18040
rect 9033 18037 9045 18040
rect 9079 18037 9091 18071
rect 9033 18031 9091 18037
rect 9122 18028 9128 18080
rect 9180 18068 9186 18080
rect 9401 18071 9459 18077
rect 9401 18068 9413 18071
rect 9180 18040 9413 18068
rect 9180 18028 9186 18040
rect 9401 18037 9413 18040
rect 9447 18037 9459 18071
rect 9401 18031 9459 18037
rect 9766 18028 9772 18080
rect 9824 18028 9830 18080
rect 11333 18071 11391 18077
rect 11333 18037 11345 18071
rect 11379 18068 11391 18071
rect 11514 18068 11520 18080
rect 11379 18040 11520 18068
rect 11379 18037 11391 18040
rect 11333 18031 11391 18037
rect 11514 18028 11520 18040
rect 11572 18028 11578 18080
rect 11900 18077 11928 18108
rect 12222 18105 12234 18108
rect 12268 18105 12280 18139
rect 12222 18099 12280 18105
rect 13709 18139 13767 18145
rect 13709 18105 13721 18139
rect 13755 18136 13767 18139
rect 13814 18136 13820 18148
rect 13755 18108 13820 18136
rect 13755 18105 13767 18108
rect 13709 18099 13767 18105
rect 13814 18096 13820 18108
rect 13872 18096 13878 18148
rect 13906 18096 13912 18148
rect 13964 18096 13970 18148
rect 14200 18136 14228 18164
rect 15194 18136 15200 18148
rect 14200 18108 15200 18136
rect 15194 18096 15200 18108
rect 15252 18096 15258 18148
rect 16945 18139 17003 18145
rect 16945 18105 16957 18139
rect 16991 18136 17003 18139
rect 17310 18136 17316 18148
rect 16991 18108 17316 18136
rect 16991 18105 17003 18108
rect 16945 18099 17003 18105
rect 17310 18096 17316 18108
rect 17368 18096 17374 18148
rect 17512 18136 17540 18164
rect 17954 18136 17960 18148
rect 17512 18108 17960 18136
rect 17954 18096 17960 18108
rect 18012 18096 18018 18148
rect 18049 18139 18107 18145
rect 18049 18105 18061 18139
rect 18095 18136 18107 18139
rect 18095 18108 18552 18136
rect 18095 18105 18107 18108
rect 18049 18099 18107 18105
rect 11885 18071 11943 18077
rect 11885 18037 11897 18071
rect 11931 18037 11943 18071
rect 11885 18031 11943 18037
rect 12986 18028 12992 18080
rect 13044 18068 13050 18080
rect 13924 18068 13952 18096
rect 13044 18040 13952 18068
rect 13044 18028 13050 18040
rect 14366 18028 14372 18080
rect 14424 18028 14430 18080
rect 14645 18071 14703 18077
rect 14645 18037 14657 18071
rect 14691 18068 14703 18071
rect 14826 18068 14832 18080
rect 14691 18040 14832 18068
rect 14691 18037 14703 18040
rect 14645 18031 14703 18037
rect 14826 18028 14832 18040
rect 14884 18068 14890 18080
rect 15746 18068 15752 18080
rect 14884 18040 15752 18068
rect 14884 18028 14890 18040
rect 15746 18028 15752 18040
rect 15804 18028 15810 18080
rect 15838 18028 15844 18080
rect 15896 18068 15902 18080
rect 18414 18068 18420 18080
rect 15896 18040 18420 18068
rect 15896 18028 15902 18040
rect 18414 18028 18420 18040
rect 18472 18028 18478 18080
rect 18524 18068 18552 18108
rect 18690 18096 18696 18148
rect 18748 18096 18754 18148
rect 18874 18096 18880 18148
rect 18932 18096 18938 18148
rect 19061 18071 19119 18077
rect 19061 18068 19073 18071
rect 18524 18040 19073 18068
rect 19061 18037 19073 18040
rect 19107 18037 19119 18071
rect 19061 18031 19119 18037
rect 19150 18028 19156 18080
rect 19208 18028 19214 18080
rect 20809 18071 20867 18077
rect 20809 18037 20821 18071
rect 20855 18068 20867 18071
rect 20898 18068 20904 18080
rect 20855 18040 20904 18068
rect 20855 18037 20867 18040
rect 20809 18031 20867 18037
rect 20898 18028 20904 18040
rect 20956 18028 20962 18080
rect 21450 18028 21456 18080
rect 21508 18028 21514 18080
rect 21542 18028 21548 18080
rect 21600 18028 21606 18080
rect 21928 18077 21956 18176
rect 22005 18173 22017 18176
rect 22051 18173 22063 18207
rect 22480 18204 22508 18235
rect 23032 18213 23060 18380
rect 22741 18207 22799 18213
rect 22741 18204 22753 18207
rect 22480 18176 22753 18204
rect 22005 18167 22063 18173
rect 22741 18173 22753 18176
rect 22787 18173 22799 18207
rect 22741 18167 22799 18173
rect 23017 18207 23075 18213
rect 23017 18173 23029 18207
rect 23063 18173 23075 18207
rect 23017 18167 23075 18173
rect 21913 18071 21971 18077
rect 21913 18037 21925 18071
rect 21959 18037 21971 18071
rect 21913 18031 21971 18037
rect 22557 18071 22615 18077
rect 22557 18037 22569 18071
rect 22603 18068 22615 18071
rect 23382 18068 23388 18080
rect 22603 18040 23388 18068
rect 22603 18037 22615 18040
rect 22557 18031 22615 18037
rect 23382 18028 23388 18040
rect 23440 18028 23446 18080
rect 552 17978 23368 18000
rect 552 17926 4366 17978
rect 4418 17926 4430 17978
rect 4482 17926 4494 17978
rect 4546 17926 4558 17978
rect 4610 17926 4622 17978
rect 4674 17926 4686 17978
rect 4738 17926 10366 17978
rect 10418 17926 10430 17978
rect 10482 17926 10494 17978
rect 10546 17926 10558 17978
rect 10610 17926 10622 17978
rect 10674 17926 10686 17978
rect 10738 17926 16366 17978
rect 16418 17926 16430 17978
rect 16482 17926 16494 17978
rect 16546 17926 16558 17978
rect 16610 17926 16622 17978
rect 16674 17926 16686 17978
rect 16738 17926 22366 17978
rect 22418 17926 22430 17978
rect 22482 17926 22494 17978
rect 22546 17926 22558 17978
rect 22610 17926 22622 17978
rect 22674 17926 22686 17978
rect 22738 17926 23368 17978
rect 552 17904 23368 17926
rect 2314 17824 2320 17876
rect 2372 17824 2378 17876
rect 2682 17824 2688 17876
rect 2740 17824 2746 17876
rect 4154 17824 4160 17876
rect 4212 17824 4218 17876
rect 4893 17867 4951 17873
rect 4893 17833 4905 17867
rect 4939 17864 4951 17867
rect 5442 17864 5448 17876
rect 4939 17836 5448 17864
rect 4939 17833 4951 17836
rect 4893 17827 4951 17833
rect 5442 17824 5448 17836
rect 5500 17824 5506 17876
rect 5718 17824 5724 17876
rect 5776 17864 5782 17876
rect 6178 17864 6184 17876
rect 5776 17836 6184 17864
rect 5776 17824 5782 17836
rect 6178 17824 6184 17836
rect 6236 17824 6242 17876
rect 6362 17824 6368 17876
rect 6420 17824 6426 17876
rect 6546 17824 6552 17876
rect 6604 17864 6610 17876
rect 7745 17867 7803 17873
rect 7745 17864 7757 17867
rect 6604 17836 7757 17864
rect 6604 17824 6610 17836
rect 7745 17833 7757 17836
rect 7791 17864 7803 17867
rect 7834 17864 7840 17876
rect 7791 17836 7840 17864
rect 7791 17833 7803 17836
rect 7745 17827 7803 17833
rect 7834 17824 7840 17836
rect 7892 17824 7898 17876
rect 7926 17824 7932 17876
rect 7984 17864 7990 17876
rect 8113 17867 8171 17873
rect 8113 17864 8125 17867
rect 7984 17836 8125 17864
rect 7984 17824 7990 17836
rect 8113 17833 8125 17836
rect 8159 17833 8171 17867
rect 8113 17827 8171 17833
rect 8754 17824 8760 17876
rect 8812 17824 8818 17876
rect 9030 17824 9036 17876
rect 9088 17864 9094 17876
rect 9088 17836 9260 17864
rect 9088 17824 9094 17836
rect 3878 17756 3884 17808
rect 3936 17756 3942 17808
rect 5258 17756 5264 17808
rect 5316 17756 5322 17808
rect 6196 17796 6224 17824
rect 6196 17768 6684 17796
rect 1210 17737 1216 17740
rect 1204 17691 1216 17737
rect 1210 17688 1216 17691
rect 1268 17688 1274 17740
rect 2409 17731 2467 17737
rect 2409 17697 2421 17731
rect 2455 17728 2467 17731
rect 2866 17728 2872 17740
rect 2455 17700 2872 17728
rect 2455 17697 2467 17700
rect 2409 17691 2467 17697
rect 2866 17688 2872 17700
rect 2924 17688 2930 17740
rect 3050 17737 3056 17740
rect 3044 17728 3056 17737
rect 3011 17700 3056 17728
rect 3044 17691 3056 17700
rect 3050 17688 3056 17691
rect 3108 17688 3114 17740
rect 3896 17728 3924 17756
rect 4617 17731 4675 17737
rect 4617 17728 4629 17731
rect 3896 17700 4629 17728
rect 4617 17697 4629 17700
rect 4663 17697 4675 17731
rect 4617 17691 4675 17697
rect 4709 17731 4767 17737
rect 4709 17697 4721 17731
rect 4755 17728 4767 17731
rect 4798 17728 4804 17740
rect 4755 17700 4804 17728
rect 4755 17697 4767 17700
rect 4709 17691 4767 17697
rect 842 17620 848 17672
rect 900 17660 906 17672
rect 937 17663 995 17669
rect 937 17660 949 17663
rect 900 17632 949 17660
rect 900 17620 906 17632
rect 937 17629 949 17632
rect 983 17629 995 17663
rect 937 17623 995 17629
rect 2682 17620 2688 17672
rect 2740 17620 2746 17672
rect 2777 17663 2835 17669
rect 2777 17629 2789 17663
rect 2823 17629 2835 17663
rect 2777 17623 2835 17629
rect 2498 17484 2504 17536
rect 2556 17484 2562 17536
rect 2792 17524 2820 17623
rect 3878 17620 3884 17672
rect 3936 17660 3942 17672
rect 4249 17663 4307 17669
rect 4249 17660 4261 17663
rect 3936 17632 4261 17660
rect 3936 17620 3942 17632
rect 4249 17629 4261 17632
rect 4295 17629 4307 17663
rect 4632 17660 4660 17691
rect 4798 17688 4804 17700
rect 4856 17688 4862 17740
rect 5997 17731 6055 17737
rect 5997 17697 6009 17731
rect 6043 17697 6055 17731
rect 5997 17691 6055 17697
rect 5350 17660 5356 17672
rect 4632 17632 5356 17660
rect 4249 17623 4307 17629
rect 5350 17620 5356 17632
rect 5408 17620 5414 17672
rect 5813 17663 5871 17669
rect 5813 17660 5825 17663
rect 5552 17632 5825 17660
rect 3694 17524 3700 17536
rect 2792 17496 3700 17524
rect 3694 17484 3700 17496
rect 3752 17484 3758 17536
rect 3786 17484 3792 17536
rect 3844 17524 3850 17536
rect 5077 17527 5135 17533
rect 5077 17524 5089 17527
rect 3844 17496 5089 17524
rect 3844 17484 3850 17496
rect 5077 17493 5089 17496
rect 5123 17493 5135 17527
rect 5077 17487 5135 17493
rect 5261 17527 5319 17533
rect 5261 17493 5273 17527
rect 5307 17524 5319 17527
rect 5552 17524 5580 17632
rect 5813 17629 5825 17632
rect 5859 17629 5871 17663
rect 6012 17660 6040 17691
rect 6086 17688 6092 17740
rect 6144 17728 6150 17740
rect 6656 17737 6684 17768
rect 6822 17756 6828 17808
rect 6880 17796 6886 17808
rect 7285 17799 7343 17805
rect 7285 17796 7297 17799
rect 6880 17768 7297 17796
rect 6880 17756 6886 17768
rect 7285 17765 7297 17768
rect 7331 17765 7343 17799
rect 7285 17759 7343 17765
rect 7374 17756 7380 17808
rect 7432 17756 7438 17808
rect 8018 17796 8024 17808
rect 7484 17768 8024 17796
rect 6273 17731 6331 17737
rect 6273 17728 6285 17731
rect 6144 17700 6285 17728
rect 6144 17688 6150 17700
rect 6273 17697 6285 17700
rect 6319 17728 6331 17731
rect 6549 17731 6607 17737
rect 6549 17728 6561 17731
rect 6319 17700 6561 17728
rect 6319 17697 6331 17700
rect 6273 17691 6331 17697
rect 6549 17697 6561 17700
rect 6595 17697 6607 17731
rect 6549 17691 6607 17697
rect 6641 17731 6699 17737
rect 6641 17697 6653 17731
rect 6687 17728 6699 17731
rect 6917 17731 6975 17737
rect 6917 17728 6929 17731
rect 6687 17700 6929 17728
rect 6687 17697 6699 17700
rect 6641 17691 6699 17697
rect 6917 17697 6929 17700
rect 6963 17697 6975 17731
rect 6917 17691 6975 17697
rect 7009 17731 7067 17737
rect 7009 17697 7021 17731
rect 7055 17697 7067 17731
rect 7009 17691 7067 17697
rect 7101 17731 7159 17737
rect 7101 17697 7113 17731
rect 7147 17728 7159 17731
rect 7484 17728 7512 17768
rect 8018 17756 8024 17768
rect 8076 17756 8082 17808
rect 8202 17756 8208 17808
rect 8260 17796 8266 17808
rect 8260 17768 9168 17796
rect 8260 17756 8266 17768
rect 8297 17731 8355 17737
rect 8297 17728 8309 17731
rect 7147 17700 7512 17728
rect 7944 17700 8309 17728
rect 7147 17697 7159 17700
rect 7101 17691 7159 17697
rect 6012 17632 6224 17660
rect 5813 17623 5871 17629
rect 5629 17595 5687 17601
rect 5629 17561 5641 17595
rect 5675 17592 5687 17595
rect 6196 17592 6224 17632
rect 6362 17620 6368 17672
rect 6420 17620 6426 17672
rect 6564 17660 6592 17691
rect 6564 17632 6960 17660
rect 6730 17592 6736 17604
rect 5675 17564 5880 17592
rect 6196 17564 6736 17592
rect 5675 17561 5687 17564
rect 5629 17555 5687 17561
rect 5307 17496 5580 17524
rect 5852 17524 5880 17564
rect 6730 17552 6736 17564
rect 6788 17552 6794 17604
rect 6086 17524 6092 17536
rect 5852 17496 6092 17524
rect 5307 17493 5319 17496
rect 5261 17487 5319 17493
rect 6086 17484 6092 17496
rect 6144 17484 6150 17536
rect 6932 17524 6960 17632
rect 7024 17592 7052 17691
rect 7944 17672 7972 17700
rect 8297 17697 8309 17700
rect 8343 17697 8355 17731
rect 8297 17691 8355 17697
rect 8386 17688 8392 17740
rect 8444 17688 8450 17740
rect 8478 17688 8484 17740
rect 8536 17688 8542 17740
rect 8938 17688 8944 17740
rect 8996 17688 9002 17740
rect 9140 17737 9168 17768
rect 9232 17737 9260 17836
rect 9306 17824 9312 17876
rect 9364 17864 9370 17876
rect 10781 17867 10839 17873
rect 10781 17864 10793 17867
rect 9364 17836 10793 17864
rect 9364 17824 9370 17836
rect 10781 17833 10793 17836
rect 10827 17864 10839 17867
rect 13725 17867 13783 17873
rect 10827 17836 12434 17864
rect 10827 17833 10839 17836
rect 10781 17827 10839 17833
rect 12406 17796 12434 17836
rect 13725 17833 13737 17867
rect 13771 17864 13783 17867
rect 13814 17864 13820 17876
rect 13771 17836 13820 17864
rect 13771 17833 13783 17836
rect 13725 17827 13783 17833
rect 13814 17824 13820 17836
rect 13872 17864 13878 17876
rect 13872 17836 14780 17864
rect 13872 17824 13878 17836
rect 13170 17796 13176 17808
rect 9416 17768 11008 17796
rect 12406 17768 13176 17796
rect 9416 17737 9444 17768
rect 10980 17740 11008 17768
rect 13170 17756 13176 17768
rect 13228 17756 13234 17808
rect 13265 17799 13323 17805
rect 13265 17765 13277 17799
rect 13311 17796 13323 17799
rect 14458 17796 14464 17808
rect 13311 17768 14464 17796
rect 13311 17765 13323 17768
rect 13265 17759 13323 17765
rect 14458 17756 14464 17768
rect 14516 17756 14522 17808
rect 9674 17737 9680 17740
rect 9125 17731 9183 17737
rect 9125 17697 9137 17731
rect 9171 17697 9183 17731
rect 9125 17691 9183 17697
rect 9217 17731 9275 17737
rect 9217 17697 9229 17731
rect 9263 17697 9275 17731
rect 9217 17691 9275 17697
rect 9401 17731 9459 17737
rect 9401 17697 9413 17731
rect 9447 17697 9459 17731
rect 9668 17728 9680 17737
rect 9635 17700 9680 17728
rect 9401 17691 9459 17697
rect 9668 17691 9680 17700
rect 9674 17688 9680 17691
rect 9732 17688 9738 17740
rect 10962 17688 10968 17740
rect 11020 17688 11026 17740
rect 11054 17688 11060 17740
rect 11112 17728 11118 17740
rect 11221 17731 11279 17737
rect 11221 17728 11233 17731
rect 11112 17700 11233 17728
rect 11112 17688 11118 17700
rect 11221 17697 11233 17700
rect 11267 17697 11279 17731
rect 11221 17691 11279 17697
rect 12621 17731 12679 17737
rect 12621 17697 12633 17731
rect 12667 17728 12679 17731
rect 12710 17728 12716 17740
rect 12667 17700 12716 17728
rect 12667 17697 12679 17700
rect 12621 17691 12679 17697
rect 12710 17688 12716 17700
rect 12768 17688 12774 17740
rect 12894 17688 12900 17740
rect 12952 17688 12958 17740
rect 12986 17688 12992 17740
rect 13044 17728 13050 17740
rect 13081 17731 13139 17737
rect 13081 17728 13093 17731
rect 13044 17700 13093 17728
rect 13044 17688 13050 17700
rect 13081 17697 13093 17700
rect 13127 17697 13139 17731
rect 13081 17691 13139 17697
rect 13817 17731 13875 17737
rect 13817 17697 13829 17731
rect 13863 17697 13875 17731
rect 13817 17691 13875 17697
rect 14093 17731 14151 17737
rect 14093 17697 14105 17731
rect 14139 17697 14151 17731
rect 14093 17691 14151 17697
rect 7558 17620 7564 17672
rect 7616 17620 7622 17672
rect 7653 17663 7711 17669
rect 7653 17629 7665 17663
rect 7699 17629 7711 17663
rect 7653 17623 7711 17629
rect 7668 17592 7696 17623
rect 7926 17620 7932 17672
rect 7984 17620 7990 17672
rect 8018 17620 8024 17672
rect 8076 17620 8082 17672
rect 9033 17663 9091 17669
rect 9033 17660 9045 17663
rect 8680 17632 9045 17660
rect 7834 17592 7840 17604
rect 7024 17564 7840 17592
rect 7834 17552 7840 17564
rect 7892 17552 7898 17604
rect 8680 17601 8708 17632
rect 9033 17629 9045 17632
rect 9079 17629 9091 17663
rect 9033 17623 9091 17629
rect 12802 17620 12808 17672
rect 12860 17620 12866 17672
rect 13357 17663 13415 17669
rect 13357 17629 13369 17663
rect 13403 17660 13415 17663
rect 13832 17660 13860 17691
rect 14001 17663 14059 17669
rect 14001 17660 14013 17663
rect 13403 17632 13768 17660
rect 13832 17632 14013 17660
rect 13403 17629 13415 17632
rect 13357 17623 13415 17629
rect 8665 17595 8723 17601
rect 8665 17561 8677 17595
rect 8711 17561 8723 17595
rect 8665 17555 8723 17561
rect 7190 17524 7196 17536
rect 6932 17496 7196 17524
rect 7190 17484 7196 17496
rect 7248 17484 7254 17536
rect 7282 17484 7288 17536
rect 7340 17524 7346 17536
rect 8680 17524 8708 17555
rect 11974 17552 11980 17604
rect 12032 17592 12038 17604
rect 13541 17595 13599 17601
rect 13541 17592 13553 17595
rect 12032 17564 13553 17592
rect 12032 17552 12038 17564
rect 13541 17561 13553 17564
rect 13587 17561 13599 17595
rect 13740 17592 13768 17632
rect 14001 17629 14013 17632
rect 14047 17629 14059 17663
rect 14108 17660 14136 17691
rect 14182 17688 14188 17740
rect 14240 17728 14246 17740
rect 14752 17737 14780 17836
rect 16942 17824 16948 17876
rect 17000 17864 17006 17876
rect 17954 17873 17960 17876
rect 17773 17867 17831 17873
rect 17773 17864 17785 17867
rect 17000 17836 17785 17864
rect 17000 17824 17006 17836
rect 17773 17833 17785 17836
rect 17819 17833 17831 17867
rect 17773 17827 17831 17833
rect 17941 17867 17960 17873
rect 17941 17833 17953 17867
rect 18012 17864 18018 17876
rect 18690 17864 18696 17876
rect 18012 17836 18696 17864
rect 17941 17827 17960 17833
rect 17954 17824 17960 17827
rect 18012 17824 18018 17836
rect 18690 17824 18696 17836
rect 18748 17824 18754 17876
rect 21085 17867 21143 17873
rect 21085 17833 21097 17867
rect 21131 17864 21143 17867
rect 21453 17867 21511 17873
rect 21131 17836 21312 17864
rect 21131 17833 21143 17836
rect 21085 17827 21143 17833
rect 15105 17799 15163 17805
rect 15105 17765 15117 17799
rect 15151 17796 15163 17799
rect 17034 17796 17040 17808
rect 15151 17768 16344 17796
rect 15151 17765 15163 17768
rect 15105 17759 15163 17765
rect 14553 17731 14611 17737
rect 14553 17728 14565 17731
rect 14240 17700 14565 17728
rect 14240 17688 14246 17700
rect 14553 17697 14565 17700
rect 14599 17697 14611 17731
rect 14553 17691 14611 17697
rect 14737 17731 14795 17737
rect 14737 17697 14749 17731
rect 14783 17697 14795 17731
rect 14737 17691 14795 17697
rect 15013 17731 15071 17737
rect 15013 17697 15025 17731
rect 15059 17697 15071 17731
rect 15013 17691 15071 17697
rect 15197 17731 15255 17737
rect 15197 17697 15209 17731
rect 15243 17697 15255 17731
rect 15197 17691 15255 17697
rect 14645 17663 14703 17669
rect 14645 17660 14657 17663
rect 14108 17632 14657 17660
rect 14001 17623 14059 17629
rect 14645 17629 14657 17632
rect 14691 17629 14703 17663
rect 14645 17623 14703 17629
rect 13906 17592 13912 17604
rect 13740 17564 13912 17592
rect 13541 17555 13599 17561
rect 13906 17552 13912 17564
rect 13964 17552 13970 17604
rect 14016 17592 14044 17623
rect 14016 17564 14504 17592
rect 7340 17496 8708 17524
rect 7340 17484 7346 17496
rect 12342 17484 12348 17536
rect 12400 17484 12406 17536
rect 12434 17484 12440 17536
rect 12492 17484 12498 17536
rect 12618 17484 12624 17536
rect 12676 17524 12682 17536
rect 12986 17524 12992 17536
rect 12676 17496 12992 17524
rect 12676 17484 12682 17496
rect 12986 17484 12992 17496
rect 13044 17484 13050 17536
rect 14274 17484 14280 17536
rect 14332 17524 14338 17536
rect 14369 17527 14427 17533
rect 14369 17524 14381 17527
rect 14332 17496 14381 17524
rect 14332 17484 14338 17496
rect 14369 17493 14381 17496
rect 14415 17493 14427 17527
rect 14476 17524 14504 17564
rect 14550 17552 14556 17604
rect 14608 17592 14614 17604
rect 15028 17592 15056 17691
rect 15212 17660 15240 17691
rect 15562 17688 15568 17740
rect 15620 17688 15626 17740
rect 15657 17731 15715 17737
rect 15657 17697 15669 17731
rect 15703 17728 15715 17731
rect 15746 17728 15752 17740
rect 15703 17700 15752 17728
rect 15703 17697 15715 17700
rect 15657 17691 15715 17697
rect 15746 17688 15752 17700
rect 15804 17688 15810 17740
rect 15838 17688 15844 17740
rect 15896 17688 15902 17740
rect 16316 17737 16344 17768
rect 16776 17768 17040 17796
rect 16776 17737 16804 17768
rect 17034 17756 17040 17768
rect 17092 17756 17098 17808
rect 18138 17756 18144 17808
rect 18196 17756 18202 17808
rect 19052 17799 19110 17805
rect 19052 17765 19064 17799
rect 19098 17796 19110 17799
rect 19150 17796 19156 17808
rect 19098 17768 19156 17796
rect 19098 17765 19110 17768
rect 19052 17759 19110 17765
rect 19150 17756 19156 17768
rect 19208 17756 19214 17808
rect 19242 17756 19248 17808
rect 19300 17796 19306 17808
rect 19300 17768 20944 17796
rect 19300 17756 19306 17768
rect 16301 17731 16359 17737
rect 16301 17697 16313 17731
rect 16347 17697 16359 17731
rect 16301 17691 16359 17697
rect 16761 17731 16819 17737
rect 16761 17697 16773 17731
rect 16807 17697 16819 17731
rect 16761 17691 16819 17697
rect 16942 17688 16948 17740
rect 17000 17688 17006 17740
rect 18782 17688 18788 17740
rect 18840 17688 18846 17740
rect 20714 17688 20720 17740
rect 20772 17688 20778 17740
rect 15289 17663 15347 17669
rect 15289 17660 15301 17663
rect 15212 17632 15301 17660
rect 15289 17629 15301 17632
rect 15335 17629 15347 17663
rect 15289 17623 15347 17629
rect 15473 17663 15531 17669
rect 15473 17629 15485 17663
rect 15519 17660 15531 17663
rect 16393 17663 16451 17669
rect 16393 17660 16405 17663
rect 15519 17632 16405 17660
rect 15519 17629 15531 17632
rect 15473 17623 15531 17629
rect 16393 17629 16405 17632
rect 16439 17660 16451 17663
rect 16853 17663 16911 17669
rect 16853 17660 16865 17663
rect 16439 17632 16865 17660
rect 16439 17629 16451 17632
rect 16393 17623 16451 17629
rect 16853 17629 16865 17632
rect 16899 17629 16911 17663
rect 16853 17623 16911 17629
rect 14608 17564 15056 17592
rect 15304 17592 15332 17623
rect 20070 17620 20076 17672
rect 20128 17660 20134 17672
rect 20441 17663 20499 17669
rect 20441 17660 20453 17663
rect 20128 17632 20453 17660
rect 20128 17620 20134 17632
rect 20441 17629 20453 17632
rect 20487 17629 20499 17663
rect 20441 17623 20499 17629
rect 20625 17663 20683 17669
rect 20625 17629 20637 17663
rect 20671 17660 20683 17663
rect 20806 17660 20812 17672
rect 20671 17632 20812 17660
rect 20671 17629 20683 17632
rect 20625 17623 20683 17629
rect 20806 17620 20812 17632
rect 20864 17620 20870 17672
rect 15749 17595 15807 17601
rect 15749 17592 15761 17595
rect 15304 17564 15761 17592
rect 14608 17552 14614 17564
rect 15749 17561 15761 17564
rect 15795 17561 15807 17595
rect 15749 17555 15807 17561
rect 16669 17595 16727 17601
rect 16669 17561 16681 17595
rect 16715 17592 16727 17595
rect 17770 17592 17776 17604
rect 16715 17564 17776 17592
rect 16715 17561 16727 17564
rect 16669 17555 16727 17561
rect 17770 17552 17776 17564
rect 17828 17552 17834 17604
rect 17880 17564 18828 17592
rect 15381 17527 15439 17533
rect 15381 17524 15393 17527
rect 14476 17496 15393 17524
rect 14369 17487 14427 17493
rect 15381 17493 15393 17496
rect 15427 17493 15439 17527
rect 15381 17487 15439 17493
rect 16022 17484 16028 17536
rect 16080 17524 16086 17536
rect 17880 17524 17908 17564
rect 16080 17496 17908 17524
rect 16080 17484 16086 17496
rect 17954 17484 17960 17536
rect 18012 17524 18018 17536
rect 18506 17524 18512 17536
rect 18012 17496 18512 17524
rect 18012 17484 18018 17496
rect 18506 17484 18512 17496
rect 18564 17484 18570 17536
rect 18800 17524 18828 17564
rect 19978 17524 19984 17536
rect 18800 17496 19984 17524
rect 19978 17484 19984 17496
rect 20036 17484 20042 17536
rect 20070 17484 20076 17536
rect 20128 17524 20134 17536
rect 20165 17527 20223 17533
rect 20165 17524 20177 17527
rect 20128 17496 20177 17524
rect 20128 17484 20134 17496
rect 20165 17493 20177 17496
rect 20211 17493 20223 17527
rect 20916 17524 20944 17768
rect 21284 17737 21312 17836
rect 21453 17833 21465 17867
rect 21499 17864 21511 17867
rect 22186 17864 22192 17876
rect 21499 17836 22192 17864
rect 21499 17833 21511 17836
rect 21453 17827 21511 17833
rect 22186 17824 22192 17836
rect 22244 17864 22250 17876
rect 23290 17864 23296 17876
rect 22244 17836 23296 17864
rect 22244 17824 22250 17836
rect 23290 17824 23296 17836
rect 23348 17824 23354 17876
rect 21893 17799 21951 17805
rect 21893 17765 21905 17799
rect 21939 17796 21951 17799
rect 22002 17796 22008 17808
rect 21939 17768 22008 17796
rect 21939 17765 21951 17768
rect 21893 17759 21951 17765
rect 22002 17756 22008 17768
rect 22060 17756 22066 17808
rect 21269 17731 21327 17737
rect 21269 17697 21281 17731
rect 21315 17728 21327 17731
rect 21358 17728 21364 17740
rect 21315 17700 21364 17728
rect 21315 17697 21327 17700
rect 21269 17691 21327 17697
rect 21358 17688 21364 17700
rect 21416 17688 21422 17740
rect 21637 17731 21695 17737
rect 21637 17697 21649 17731
rect 21683 17728 21695 17731
rect 21726 17728 21732 17740
rect 21683 17700 21732 17728
rect 21683 17697 21695 17700
rect 21637 17691 21695 17697
rect 21726 17688 21732 17700
rect 21784 17688 21790 17740
rect 23017 17527 23075 17533
rect 23017 17524 23029 17527
rect 20916 17496 23029 17524
rect 20165 17487 20223 17493
rect 23017 17493 23029 17496
rect 23063 17493 23075 17527
rect 23017 17487 23075 17493
rect 552 17434 23368 17456
rect 552 17382 1366 17434
rect 1418 17382 1430 17434
rect 1482 17382 1494 17434
rect 1546 17382 1558 17434
rect 1610 17382 1622 17434
rect 1674 17382 1686 17434
rect 1738 17382 7366 17434
rect 7418 17382 7430 17434
rect 7482 17382 7494 17434
rect 7546 17382 7558 17434
rect 7610 17382 7622 17434
rect 7674 17382 7686 17434
rect 7738 17382 13366 17434
rect 13418 17382 13430 17434
rect 13482 17382 13494 17434
rect 13546 17382 13558 17434
rect 13610 17382 13622 17434
rect 13674 17382 13686 17434
rect 13738 17382 19366 17434
rect 19418 17382 19430 17434
rect 19482 17382 19494 17434
rect 19546 17382 19558 17434
rect 19610 17382 19622 17434
rect 19674 17382 19686 17434
rect 19738 17382 23368 17434
rect 552 17360 23368 17382
rect 1210 17280 1216 17332
rect 1268 17320 1274 17332
rect 1581 17323 1639 17329
rect 1581 17320 1593 17323
rect 1268 17292 1593 17320
rect 1268 17280 1274 17292
rect 1581 17289 1593 17292
rect 1627 17289 1639 17323
rect 1581 17283 1639 17289
rect 2225 17323 2283 17329
rect 2225 17289 2237 17323
rect 2271 17320 2283 17323
rect 2498 17320 2504 17332
rect 2271 17292 2504 17320
rect 2271 17289 2283 17292
rect 2225 17283 2283 17289
rect 2498 17280 2504 17292
rect 2556 17280 2562 17332
rect 2685 17323 2743 17329
rect 2685 17289 2697 17323
rect 2731 17320 2743 17323
rect 2774 17320 2780 17332
rect 2731 17292 2780 17320
rect 2731 17289 2743 17292
rect 2685 17283 2743 17289
rect 2774 17280 2780 17292
rect 2832 17280 2838 17332
rect 2866 17280 2872 17332
rect 2924 17320 2930 17332
rect 3050 17320 3056 17332
rect 2924 17292 3056 17320
rect 2924 17280 2930 17292
rect 3050 17280 3056 17292
rect 3108 17280 3114 17332
rect 6178 17280 6184 17332
rect 6236 17280 6242 17332
rect 6362 17280 6368 17332
rect 6420 17320 6426 17332
rect 6641 17323 6699 17329
rect 6641 17320 6653 17323
rect 6420 17292 6653 17320
rect 6420 17280 6426 17292
rect 6641 17289 6653 17292
rect 6687 17289 6699 17323
rect 7098 17320 7104 17332
rect 6641 17283 6699 17289
rect 6748 17292 7104 17320
rect 5261 17255 5319 17261
rect 5261 17221 5273 17255
rect 5307 17252 5319 17255
rect 5626 17252 5632 17264
rect 5307 17224 5632 17252
rect 5307 17221 5319 17224
rect 5261 17215 5319 17221
rect 5626 17212 5632 17224
rect 5684 17212 5690 17264
rect 6089 17255 6147 17261
rect 6089 17221 6101 17255
rect 6135 17252 6147 17255
rect 6748 17252 6776 17292
rect 7098 17280 7104 17292
rect 7156 17280 7162 17332
rect 7190 17280 7196 17332
rect 7248 17320 7254 17332
rect 7469 17323 7527 17329
rect 7248 17292 7420 17320
rect 7248 17280 7254 17292
rect 6135 17224 6776 17252
rect 6135 17221 6147 17224
rect 6089 17215 6147 17221
rect 3602 17184 3608 17196
rect 1320 17156 3608 17184
rect 1320 17125 1348 17156
rect 3602 17144 3608 17156
rect 3660 17144 3666 17196
rect 5534 17184 5540 17196
rect 5000 17156 5540 17184
rect 1305 17119 1363 17125
rect 1305 17085 1317 17119
rect 1351 17085 1363 17119
rect 1305 17079 1363 17085
rect 1581 17119 1639 17125
rect 1581 17085 1593 17119
rect 1627 17116 1639 17119
rect 1670 17116 1676 17128
rect 1627 17088 1676 17116
rect 1627 17085 1639 17088
rect 1581 17079 1639 17085
rect 1670 17076 1676 17088
rect 1728 17076 1734 17128
rect 1765 17119 1823 17125
rect 1765 17085 1777 17119
rect 1811 17085 1823 17119
rect 1765 17079 1823 17085
rect 1780 17048 1808 17079
rect 1946 17076 1952 17128
rect 2004 17076 2010 17128
rect 2038 17076 2044 17128
rect 2096 17116 2102 17128
rect 2866 17116 2872 17128
rect 2096 17088 2872 17116
rect 2096 17076 2102 17088
rect 2866 17076 2872 17088
rect 2924 17076 2930 17128
rect 2958 17076 2964 17128
rect 3016 17116 3022 17128
rect 5000 17125 5028 17156
rect 5534 17144 5540 17156
rect 5592 17144 5598 17196
rect 6104 17184 6132 17215
rect 6822 17212 6828 17264
rect 6880 17252 6886 17264
rect 7285 17255 7343 17261
rect 7285 17252 7297 17255
rect 6880 17224 7297 17252
rect 6880 17212 6886 17224
rect 7285 17221 7297 17224
rect 7331 17221 7343 17255
rect 7392 17252 7420 17292
rect 7469 17289 7481 17323
rect 7515 17320 7527 17323
rect 7926 17320 7932 17332
rect 7515 17292 7932 17320
rect 7515 17289 7527 17292
rect 7469 17283 7527 17289
rect 7926 17280 7932 17292
rect 7984 17280 7990 17332
rect 8662 17280 8668 17332
rect 8720 17320 8726 17332
rect 8757 17323 8815 17329
rect 8757 17320 8769 17323
rect 8720 17292 8769 17320
rect 8720 17280 8726 17292
rect 8757 17289 8769 17292
rect 8803 17289 8815 17323
rect 8757 17283 8815 17289
rect 9582 17280 9588 17332
rect 9640 17280 9646 17332
rect 10781 17323 10839 17329
rect 10781 17289 10793 17323
rect 10827 17320 10839 17323
rect 11054 17320 11060 17332
rect 10827 17292 11060 17320
rect 10827 17289 10839 17292
rect 10781 17283 10839 17289
rect 11054 17280 11060 17292
rect 11112 17280 11118 17332
rect 11333 17323 11391 17329
rect 11333 17289 11345 17323
rect 11379 17320 11391 17323
rect 11422 17320 11428 17332
rect 11379 17292 11428 17320
rect 11379 17289 11391 17292
rect 11333 17283 11391 17289
rect 11422 17280 11428 17292
rect 11480 17280 11486 17332
rect 11517 17323 11575 17329
rect 11517 17289 11529 17323
rect 11563 17320 11575 17323
rect 11698 17320 11704 17332
rect 11563 17292 11704 17320
rect 11563 17289 11575 17292
rect 11517 17283 11575 17289
rect 11698 17280 11704 17292
rect 11756 17280 11762 17332
rect 13633 17323 13691 17329
rect 13633 17289 13645 17323
rect 13679 17320 13691 17323
rect 13814 17320 13820 17332
rect 13679 17292 13820 17320
rect 13679 17289 13691 17292
rect 13633 17283 13691 17289
rect 13814 17280 13820 17292
rect 13872 17280 13878 17332
rect 13906 17280 13912 17332
rect 13964 17320 13970 17332
rect 14185 17323 14243 17329
rect 14185 17320 14197 17323
rect 13964 17292 14197 17320
rect 13964 17280 13970 17292
rect 14185 17289 14197 17292
rect 14231 17289 14243 17323
rect 14185 17283 14243 17289
rect 15562 17280 15568 17332
rect 15620 17320 15626 17332
rect 15841 17323 15899 17329
rect 15841 17320 15853 17323
rect 15620 17292 15853 17320
rect 15620 17280 15626 17292
rect 15841 17289 15853 17292
rect 15887 17289 15899 17323
rect 15841 17283 15899 17289
rect 16666 17280 16672 17332
rect 16724 17320 16730 17332
rect 16853 17323 16911 17329
rect 16853 17320 16865 17323
rect 16724 17292 16865 17320
rect 16724 17280 16730 17292
rect 16853 17289 16865 17292
rect 16899 17320 16911 17323
rect 16942 17320 16948 17332
rect 16899 17292 16948 17320
rect 16899 17289 16911 17292
rect 16853 17283 16911 17289
rect 16942 17280 16948 17292
rect 17000 17280 17006 17332
rect 18046 17280 18052 17332
rect 18104 17320 18110 17332
rect 19886 17320 19892 17332
rect 18104 17292 19892 17320
rect 18104 17280 18110 17292
rect 19886 17280 19892 17292
rect 19944 17280 19950 17332
rect 21266 17280 21272 17332
rect 21324 17320 21330 17332
rect 23382 17320 23388 17332
rect 21324 17292 23388 17320
rect 21324 17280 21330 17292
rect 23382 17280 23388 17292
rect 23440 17280 23446 17332
rect 7561 17255 7619 17261
rect 7561 17252 7573 17255
rect 7392 17224 7573 17252
rect 7285 17215 7343 17221
rect 7561 17221 7573 17224
rect 7607 17252 7619 17255
rect 8389 17255 8447 17261
rect 8389 17252 8401 17255
rect 7607 17224 8401 17252
rect 7607 17221 7619 17224
rect 7561 17215 7619 17221
rect 8389 17221 8401 17224
rect 8435 17221 8447 17255
rect 9766 17252 9772 17264
rect 8389 17215 8447 17221
rect 8496 17224 9772 17252
rect 5644 17156 6132 17184
rect 4985 17119 5043 17125
rect 3016 17088 3924 17116
rect 3016 17076 3022 17088
rect 2498 17048 2504 17060
rect 1780 17020 2504 17048
rect 2498 17008 2504 17020
rect 2556 17008 2562 17060
rect 3068 17057 3096 17088
rect 3053 17051 3111 17057
rect 3053 17017 3065 17051
rect 3099 17017 3111 17051
rect 3896 17048 3924 17088
rect 4985 17085 4997 17119
rect 5031 17085 5043 17119
rect 4985 17079 5043 17085
rect 5074 17076 5080 17128
rect 5132 17076 5138 17128
rect 5644 17116 5672 17156
rect 5184 17088 5672 17116
rect 5184 17048 5212 17088
rect 5810 17076 5816 17128
rect 5868 17116 5874 17128
rect 5905 17119 5963 17125
rect 5905 17116 5917 17119
rect 5868 17088 5917 17116
rect 5868 17076 5874 17088
rect 5905 17085 5917 17088
rect 5951 17085 5963 17119
rect 5905 17079 5963 17085
rect 6362 17076 6368 17128
rect 6420 17076 6426 17128
rect 7745 17119 7803 17125
rect 7745 17116 7757 17119
rect 6640 17091 7757 17116
rect 6595 17088 7757 17091
rect 6595 17085 6668 17088
rect 3053 17011 3111 17017
rect 3620 17020 3832 17048
rect 3896 17020 5212 17048
rect 1118 16940 1124 16992
rect 1176 16940 1182 16992
rect 2866 16989 2872 16992
rect 2853 16983 2872 16989
rect 2853 16949 2865 16983
rect 2924 16980 2930 16992
rect 3620 16980 3648 17020
rect 2924 16952 3648 16980
rect 2853 16943 2872 16949
rect 2866 16940 2872 16943
rect 2924 16940 2930 16952
rect 3694 16940 3700 16992
rect 3752 16940 3758 16992
rect 3804 16980 3832 17020
rect 5442 17008 5448 17060
rect 5500 17008 5506 17060
rect 5629 17051 5687 17057
rect 5629 17017 5641 17051
rect 5675 17048 5687 17051
rect 6270 17048 6276 17060
rect 5675 17020 6276 17048
rect 5675 17017 5687 17020
rect 5629 17011 5687 17017
rect 6270 17008 6276 17020
rect 6328 17008 6334 17060
rect 6595 17051 6607 17085
rect 6641 17054 6668 17085
rect 7745 17085 7757 17088
rect 7791 17116 7803 17119
rect 8496 17116 8524 17224
rect 9766 17212 9772 17224
rect 9824 17212 9830 17264
rect 10229 17255 10287 17261
rect 10229 17221 10241 17255
rect 10275 17221 10287 17255
rect 16758 17252 16764 17264
rect 10229 17215 10287 17221
rect 11624 17224 16764 17252
rect 9306 17144 9312 17196
rect 9364 17184 9370 17196
rect 9493 17187 9551 17193
rect 9493 17184 9505 17187
rect 9364 17156 9505 17184
rect 9364 17144 9370 17156
rect 9493 17153 9505 17156
rect 9539 17184 9551 17187
rect 10244 17184 10272 17215
rect 9539 17156 10272 17184
rect 10413 17187 10471 17193
rect 9539 17153 9551 17156
rect 9493 17147 9551 17153
rect 10413 17153 10425 17187
rect 10459 17184 10471 17187
rect 10459 17156 10640 17184
rect 10459 17153 10471 17156
rect 10413 17147 10471 17153
rect 9033 17119 9091 17125
rect 9033 17116 9045 17119
rect 7791 17088 8524 17116
rect 8956 17088 9045 17116
rect 7791 17085 7803 17088
rect 7745 17079 7803 17085
rect 6641 17051 6653 17054
rect 6595 17045 6653 17051
rect 6825 17051 6883 17057
rect 6825 17017 6837 17051
rect 6871 17017 6883 17051
rect 6825 17011 6883 17017
rect 6086 16980 6092 16992
rect 3804 16952 6092 16980
rect 6086 16940 6092 16952
rect 6144 16980 6150 16992
rect 6457 16983 6515 16989
rect 6457 16980 6469 16983
rect 6144 16952 6469 16980
rect 6144 16940 6150 16952
rect 6457 16949 6469 16952
rect 6503 16949 6515 16983
rect 6457 16943 6515 16949
rect 6730 16940 6736 16992
rect 6788 16980 6794 16992
rect 6840 16980 6868 17011
rect 7006 17008 7012 17060
rect 7064 17008 7070 17060
rect 8570 16980 8576 16992
rect 6788 16952 8576 16980
rect 6788 16940 6794 16952
rect 8570 16940 8576 16952
rect 8628 16940 8634 16992
rect 8754 16940 8760 16992
rect 8812 16940 8818 16992
rect 8956 16989 8984 17088
rect 9033 17085 9045 17088
rect 9079 17085 9091 17119
rect 9033 17079 9091 17085
rect 9582 17076 9588 17128
rect 9640 17116 9646 17128
rect 10612 17125 10640 17156
rect 10870 17144 10876 17196
rect 10928 17184 10934 17196
rect 11624 17193 11652 17224
rect 16758 17212 16764 17224
rect 16816 17212 16822 17264
rect 18414 17212 18420 17264
rect 18472 17252 18478 17264
rect 21358 17252 21364 17264
rect 18472 17224 21364 17252
rect 18472 17212 18478 17224
rect 21358 17212 21364 17224
rect 21416 17212 21422 17264
rect 11609 17187 11667 17193
rect 11609 17184 11621 17187
rect 10928 17156 11621 17184
rect 10928 17144 10934 17156
rect 11609 17153 11621 17156
rect 11655 17153 11667 17187
rect 12434 17184 12440 17196
rect 11609 17147 11667 17153
rect 12406 17144 12440 17184
rect 12492 17144 12498 17196
rect 13170 17144 13176 17196
rect 13228 17184 13234 17196
rect 13228 17156 14688 17184
rect 13228 17144 13234 17156
rect 9677 17119 9735 17125
rect 9677 17116 9689 17119
rect 9640 17088 9689 17116
rect 9640 17076 9646 17088
rect 9677 17085 9689 17088
rect 9723 17085 9735 17119
rect 9677 17079 9735 17085
rect 9769 17119 9827 17125
rect 9769 17085 9781 17119
rect 9815 17085 9827 17119
rect 9769 17079 9827 17085
rect 10597 17119 10655 17125
rect 10597 17085 10609 17119
rect 10643 17085 10655 17119
rect 12406 17116 12434 17144
rect 10597 17079 10655 17085
rect 10704 17088 12434 17116
rect 9122 17008 9128 17060
rect 9180 17048 9186 17060
rect 9784 17048 9812 17079
rect 9180 17020 9812 17048
rect 9180 17008 9186 17020
rect 9950 17008 9956 17060
rect 10008 17008 10014 17060
rect 8941 16983 8999 16989
rect 8941 16949 8953 16983
rect 8987 16949 8999 16983
rect 8941 16943 8999 16949
rect 9217 16983 9275 16989
rect 9217 16949 9229 16983
rect 9263 16980 9275 16983
rect 9306 16980 9312 16992
rect 9263 16952 9312 16980
rect 9263 16949 9275 16952
rect 9217 16943 9275 16949
rect 9306 16940 9312 16952
rect 9364 16940 9370 16992
rect 9582 16940 9588 16992
rect 9640 16980 9646 16992
rect 10704 16980 10732 17088
rect 13262 17076 13268 17128
rect 13320 17116 13326 17128
rect 13357 17119 13415 17125
rect 13357 17116 13369 17119
rect 13320 17088 13369 17116
rect 13320 17076 13326 17088
rect 13357 17085 13369 17088
rect 13403 17085 13415 17119
rect 13357 17079 13415 17085
rect 13906 17076 13912 17128
rect 13964 17116 13970 17128
rect 14093 17119 14151 17125
rect 14093 17116 14105 17119
rect 13964 17088 14105 17116
rect 13964 17076 13970 17088
rect 14093 17085 14105 17088
rect 14139 17085 14151 17119
rect 14093 17079 14151 17085
rect 14277 17119 14335 17125
rect 14277 17085 14289 17119
rect 14323 17116 14335 17119
rect 14366 17116 14372 17128
rect 14323 17088 14372 17116
rect 14323 17085 14335 17088
rect 14277 17079 14335 17085
rect 14366 17076 14372 17088
rect 14424 17076 14430 17128
rect 14660 17125 14688 17156
rect 14918 17144 14924 17196
rect 14976 17184 14982 17196
rect 16666 17184 16672 17196
rect 14976 17156 16672 17184
rect 14976 17144 14982 17156
rect 16666 17144 16672 17156
rect 16724 17144 16730 17196
rect 16776 17184 16804 17212
rect 16776 17156 19472 17184
rect 14553 17119 14611 17125
rect 14553 17085 14565 17119
rect 14599 17085 14611 17119
rect 14553 17079 14611 17085
rect 14645 17119 14703 17125
rect 14645 17085 14657 17119
rect 14691 17116 14703 17119
rect 15105 17119 15163 17125
rect 15105 17116 15117 17119
rect 14691 17088 15117 17116
rect 14691 17085 14703 17088
rect 14645 17079 14703 17085
rect 15105 17085 15117 17088
rect 15151 17085 15163 17119
rect 15105 17079 15163 17085
rect 15381 17119 15439 17125
rect 15381 17085 15393 17119
rect 15427 17085 15439 17119
rect 15381 17079 15439 17085
rect 10778 17008 10784 17060
rect 10836 17048 10842 17060
rect 11149 17051 11207 17057
rect 11149 17048 11161 17051
rect 10836 17020 11161 17048
rect 10836 17008 10842 17020
rect 11149 17017 11161 17020
rect 11195 17017 11207 17051
rect 11149 17011 11207 17017
rect 11330 17008 11336 17060
rect 11388 17057 11394 17060
rect 11388 17051 11407 17057
rect 11395 17017 11407 17051
rect 11388 17011 11407 17017
rect 11388 17008 11394 17011
rect 12710 17008 12716 17060
rect 12768 17048 12774 17060
rect 12986 17048 12992 17060
rect 12768 17020 12992 17048
rect 12768 17008 12774 17020
rect 12986 17008 12992 17020
rect 13044 17008 13050 17060
rect 13078 17008 13084 17060
rect 13136 17048 13142 17060
rect 13630 17048 13636 17060
rect 13136 17020 13636 17048
rect 13136 17008 13142 17020
rect 13630 17008 13636 17020
rect 13688 17048 13694 17060
rect 13817 17051 13875 17057
rect 13817 17048 13829 17051
rect 13688 17020 13829 17048
rect 13688 17008 13694 17020
rect 13817 17017 13829 17020
rect 13863 17017 13875 17051
rect 13817 17011 13875 17017
rect 9640 16952 10732 16980
rect 13832 16980 13860 17011
rect 13998 17008 14004 17060
rect 14056 17008 14062 17060
rect 14568 17048 14596 17079
rect 14200 17020 14596 17048
rect 14200 16980 14228 17020
rect 14734 17008 14740 17060
rect 14792 17048 14798 17060
rect 14829 17051 14887 17057
rect 14829 17048 14841 17051
rect 14792 17020 14841 17048
rect 14792 17008 14798 17020
rect 14829 17017 14841 17020
rect 14875 17017 14887 17051
rect 14829 17011 14887 17017
rect 15013 17051 15071 17057
rect 15013 17017 15025 17051
rect 15059 17048 15071 17051
rect 15396 17048 15424 17079
rect 15470 17076 15476 17128
rect 15528 17116 15534 17128
rect 15565 17119 15623 17125
rect 15565 17116 15577 17119
rect 15528 17088 15577 17116
rect 15528 17076 15534 17088
rect 15565 17085 15577 17088
rect 15611 17085 15623 17119
rect 15565 17079 15623 17085
rect 15657 17119 15715 17125
rect 15657 17085 15669 17119
rect 15703 17116 15715 17119
rect 15746 17116 15752 17128
rect 15703 17088 15752 17116
rect 15703 17085 15715 17088
rect 15657 17079 15715 17085
rect 15746 17076 15752 17088
rect 15804 17076 15810 17128
rect 15841 17119 15899 17125
rect 15841 17085 15853 17119
rect 15887 17116 15899 17119
rect 15933 17119 15991 17125
rect 15933 17116 15945 17119
rect 15887 17088 15945 17116
rect 15887 17085 15899 17088
rect 15841 17079 15899 17085
rect 15933 17085 15945 17088
rect 15979 17116 15991 17119
rect 17497 17119 17555 17125
rect 17497 17116 17509 17119
rect 15979 17088 17509 17116
rect 15979 17085 15991 17088
rect 15933 17079 15991 17085
rect 17497 17085 17509 17088
rect 17543 17116 17555 17119
rect 17543 17088 17816 17116
rect 17543 17085 17555 17088
rect 17497 17079 17555 17085
rect 17037 17051 17095 17057
rect 15059 17020 15424 17048
rect 15488 17020 16988 17048
rect 15059 17017 15071 17020
rect 15013 17011 15071 17017
rect 13832 16952 14228 16980
rect 9640 16940 9646 16952
rect 14366 16940 14372 16992
rect 14424 16940 14430 16992
rect 14550 16940 14556 16992
rect 14608 16980 14614 16992
rect 15289 16983 15347 16989
rect 15289 16980 15301 16983
rect 14608 16952 15301 16980
rect 14608 16940 14614 16952
rect 15289 16949 15301 16952
rect 15335 16980 15347 16983
rect 15488 16980 15516 17020
rect 15335 16952 15516 16980
rect 15335 16949 15347 16952
rect 15289 16943 15347 16949
rect 15562 16940 15568 16992
rect 15620 16940 15626 16992
rect 15930 16940 15936 16992
rect 15988 16980 15994 16992
rect 16117 16983 16175 16989
rect 16117 16980 16129 16983
rect 15988 16952 16129 16980
rect 15988 16940 15994 16952
rect 16117 16949 16129 16952
rect 16163 16949 16175 16983
rect 16117 16943 16175 16949
rect 16666 16940 16672 16992
rect 16724 16940 16730 16992
rect 16850 16989 16856 16992
rect 16837 16983 16856 16989
rect 16837 16949 16849 16983
rect 16837 16943 16856 16949
rect 16850 16940 16856 16943
rect 16908 16940 16914 16992
rect 16960 16980 16988 17020
rect 17037 17017 17049 17051
rect 17083 17048 17095 17051
rect 17402 17048 17408 17060
rect 17083 17020 17408 17048
rect 17083 17017 17095 17020
rect 17037 17011 17095 17017
rect 17402 17008 17408 17020
rect 17460 17048 17466 17060
rect 17678 17048 17684 17060
rect 17460 17020 17684 17048
rect 17460 17008 17466 17020
rect 17678 17008 17684 17020
rect 17736 17008 17742 17060
rect 17218 16980 17224 16992
rect 16960 16952 17224 16980
rect 17218 16940 17224 16952
rect 17276 16940 17282 16992
rect 17788 16980 17816 17088
rect 18046 17076 18052 17128
rect 18104 17116 18110 17128
rect 18141 17119 18199 17125
rect 18141 17116 18153 17119
rect 18104 17088 18153 17116
rect 18104 17076 18110 17088
rect 18141 17085 18153 17088
rect 18187 17085 18199 17119
rect 18141 17079 18199 17085
rect 18233 17119 18291 17125
rect 18233 17085 18245 17119
rect 18279 17116 18291 17119
rect 18322 17116 18328 17128
rect 18279 17088 18328 17116
rect 18279 17085 18291 17088
rect 18233 17079 18291 17085
rect 18322 17076 18328 17088
rect 18380 17076 18386 17128
rect 18414 17076 18420 17128
rect 18472 17076 18478 17128
rect 19444 17125 19472 17156
rect 20806 17144 20812 17196
rect 20864 17184 20870 17196
rect 21269 17187 21327 17193
rect 21269 17184 21281 17187
rect 20864 17156 21281 17184
rect 20864 17144 20870 17156
rect 21269 17153 21281 17156
rect 21315 17153 21327 17187
rect 21269 17147 21327 17153
rect 18693 17119 18751 17125
rect 18693 17085 18705 17119
rect 18739 17085 18751 17119
rect 18877 17119 18935 17125
rect 18877 17116 18889 17119
rect 18693 17079 18751 17085
rect 18800 17088 18889 17116
rect 17865 17051 17923 17057
rect 17865 17017 17877 17051
rect 17911 17048 17923 17051
rect 18708 17048 18736 17079
rect 17911 17020 18736 17048
rect 17911 17017 17923 17020
rect 17865 17011 17923 17017
rect 18800 16992 18828 17088
rect 18877 17085 18889 17088
rect 18923 17085 18935 17119
rect 18877 17079 18935 17085
rect 19429 17119 19487 17125
rect 19429 17085 19441 17119
rect 19475 17085 19487 17119
rect 19429 17079 19487 17085
rect 21177 17119 21235 17125
rect 21177 17085 21189 17119
rect 21223 17116 21235 17119
rect 21637 17119 21695 17125
rect 21637 17116 21649 17119
rect 21223 17088 21649 17116
rect 21223 17085 21235 17088
rect 21177 17079 21235 17085
rect 21637 17085 21649 17088
rect 21683 17116 21695 17119
rect 21726 17116 21732 17128
rect 21683 17088 21732 17116
rect 21683 17085 21695 17088
rect 21637 17079 21695 17085
rect 21726 17076 21732 17088
rect 21784 17076 21790 17128
rect 21904 17119 21962 17125
rect 21904 17085 21916 17119
rect 21950 17116 21962 17119
rect 22186 17116 22192 17128
rect 21950 17088 22192 17116
rect 21950 17085 21962 17088
rect 21904 17079 21962 17085
rect 22186 17076 22192 17088
rect 22244 17076 22250 17128
rect 19150 17008 19156 17060
rect 19208 17008 19214 17060
rect 19334 17008 19340 17060
rect 19392 17008 19398 17060
rect 19978 17008 19984 17060
rect 20036 17048 20042 17060
rect 21453 17051 21511 17057
rect 21453 17048 21465 17051
rect 20036 17020 21465 17048
rect 20036 17008 20042 17020
rect 21453 17017 21465 17020
rect 21499 17048 21511 17051
rect 21499 17020 22094 17048
rect 21499 17017 21511 17020
rect 21453 17011 21511 17017
rect 17957 16983 18015 16989
rect 17957 16980 17969 16983
rect 17788 16952 17969 16980
rect 17957 16949 17969 16952
rect 18003 16980 18015 16983
rect 18322 16980 18328 16992
rect 18003 16952 18328 16980
rect 18003 16949 18015 16952
rect 17957 16943 18015 16949
rect 18322 16940 18328 16952
rect 18380 16940 18386 16992
rect 18417 16983 18475 16989
rect 18417 16949 18429 16983
rect 18463 16980 18475 16983
rect 18782 16980 18788 16992
rect 18463 16952 18788 16980
rect 18463 16949 18475 16952
rect 18417 16943 18475 16949
rect 18782 16940 18788 16952
rect 18840 16940 18846 16992
rect 18874 16940 18880 16992
rect 18932 16940 18938 16992
rect 22066 16980 22094 17020
rect 23017 16983 23075 16989
rect 23017 16980 23029 16983
rect 22066 16952 23029 16980
rect 23017 16949 23029 16952
rect 23063 16949 23075 16983
rect 23017 16943 23075 16949
rect 552 16890 23368 16912
rect 552 16838 4366 16890
rect 4418 16838 4430 16890
rect 4482 16838 4494 16890
rect 4546 16838 4558 16890
rect 4610 16838 4622 16890
rect 4674 16838 4686 16890
rect 4738 16838 10366 16890
rect 10418 16838 10430 16890
rect 10482 16838 10494 16890
rect 10546 16838 10558 16890
rect 10610 16838 10622 16890
rect 10674 16838 10686 16890
rect 10738 16838 16366 16890
rect 16418 16838 16430 16890
rect 16482 16838 16494 16890
rect 16546 16838 16558 16890
rect 16610 16838 16622 16890
rect 16674 16838 16686 16890
rect 16738 16838 22366 16890
rect 22418 16838 22430 16890
rect 22482 16838 22494 16890
rect 22546 16838 22558 16890
rect 22610 16838 22622 16890
rect 22674 16838 22686 16890
rect 22738 16838 23368 16890
rect 552 16816 23368 16838
rect 952 16748 3740 16776
rect 842 16600 848 16652
rect 900 16640 906 16652
rect 952 16649 980 16748
rect 3712 16720 3740 16748
rect 3878 16736 3884 16788
rect 3936 16736 3942 16788
rect 3970 16736 3976 16788
rect 4028 16776 4034 16788
rect 4249 16779 4307 16785
rect 4249 16776 4261 16779
rect 4028 16748 4261 16776
rect 4028 16736 4034 16748
rect 4249 16745 4261 16748
rect 4295 16745 4307 16779
rect 4249 16739 4307 16745
rect 4338 16736 4344 16788
rect 4396 16776 4402 16788
rect 4433 16779 4491 16785
rect 4433 16776 4445 16779
rect 4396 16748 4445 16776
rect 4396 16736 4402 16748
rect 4433 16745 4445 16748
rect 4479 16745 4491 16779
rect 4433 16739 4491 16745
rect 4522 16736 4528 16788
rect 4580 16776 4586 16788
rect 5074 16776 5080 16788
rect 4580 16748 5080 16776
rect 4580 16736 4586 16748
rect 5074 16736 5080 16748
rect 5132 16736 5138 16788
rect 5258 16736 5264 16788
rect 5316 16776 5322 16788
rect 5399 16779 5457 16785
rect 5399 16776 5411 16779
rect 5316 16748 5411 16776
rect 5316 16736 5322 16748
rect 5399 16745 5411 16748
rect 5445 16776 5457 16779
rect 6638 16776 6644 16788
rect 5445 16748 6644 16776
rect 5445 16745 5457 16748
rect 5399 16739 5457 16745
rect 6638 16736 6644 16748
rect 6696 16736 6702 16788
rect 7282 16736 7288 16788
rect 7340 16776 7346 16788
rect 7653 16779 7711 16785
rect 7653 16776 7665 16779
rect 7340 16748 7665 16776
rect 7340 16736 7346 16748
rect 7653 16745 7665 16748
rect 7699 16745 7711 16779
rect 7653 16739 7711 16745
rect 7834 16736 7840 16788
rect 7892 16736 7898 16788
rect 8113 16779 8171 16785
rect 8113 16745 8125 16779
rect 8159 16776 8171 16779
rect 8478 16776 8484 16788
rect 8159 16748 8484 16776
rect 8159 16745 8171 16748
rect 8113 16739 8171 16745
rect 8478 16736 8484 16748
rect 8536 16736 8542 16788
rect 9030 16776 9036 16788
rect 8772 16748 9036 16776
rect 1204 16711 1262 16717
rect 1204 16677 1216 16711
rect 1250 16708 1262 16711
rect 3145 16711 3203 16717
rect 3145 16708 3157 16711
rect 1250 16680 3157 16708
rect 1250 16677 1262 16680
rect 1204 16671 1262 16677
rect 3145 16677 3157 16680
rect 3191 16677 3203 16711
rect 3145 16671 3203 16677
rect 3694 16668 3700 16720
rect 3752 16708 3758 16720
rect 8297 16711 8355 16717
rect 3752 16680 8064 16708
rect 3752 16668 3758 16680
rect 937 16643 995 16649
rect 937 16640 949 16643
rect 900 16612 949 16640
rect 900 16600 906 16612
rect 937 16609 949 16612
rect 983 16609 995 16643
rect 937 16603 995 16609
rect 2406 16600 2412 16652
rect 2464 16600 2470 16652
rect 2498 16600 2504 16652
rect 2556 16640 2562 16652
rect 2593 16643 2651 16649
rect 2593 16640 2605 16643
rect 2556 16612 2605 16640
rect 2556 16600 2562 16612
rect 2593 16609 2605 16612
rect 2639 16609 2651 16643
rect 2593 16603 2651 16609
rect 2682 16600 2688 16652
rect 2740 16600 2746 16652
rect 2777 16643 2835 16649
rect 2777 16609 2789 16643
rect 2823 16609 2835 16643
rect 2777 16603 2835 16609
rect 3421 16643 3479 16649
rect 3421 16609 3433 16643
rect 3467 16609 3479 16643
rect 3421 16603 3479 16609
rect 2314 16396 2320 16448
rect 2372 16396 2378 16448
rect 2682 16396 2688 16448
rect 2740 16436 2746 16448
rect 2792 16436 2820 16603
rect 3436 16572 3464 16603
rect 3510 16600 3516 16652
rect 3568 16600 3574 16652
rect 3602 16600 3608 16652
rect 3660 16600 3666 16652
rect 3786 16600 3792 16652
rect 3844 16600 3850 16652
rect 4062 16600 4068 16652
rect 4120 16600 4126 16652
rect 4157 16643 4215 16649
rect 4157 16609 4169 16643
rect 4203 16609 4215 16643
rect 4157 16603 4215 16609
rect 4172 16572 4200 16603
rect 4246 16600 4252 16652
rect 4304 16640 4310 16652
rect 4525 16643 4583 16649
rect 4525 16640 4537 16643
rect 4304 16612 4537 16640
rect 4304 16600 4310 16612
rect 4525 16609 4537 16612
rect 4571 16609 4583 16643
rect 5166 16640 5172 16652
rect 4525 16603 4583 16609
rect 4632 16612 5172 16640
rect 4632 16572 4660 16612
rect 5166 16600 5172 16612
rect 5224 16600 5230 16652
rect 5626 16600 5632 16652
rect 5684 16600 5690 16652
rect 5828 16649 5856 16680
rect 5813 16643 5871 16649
rect 5813 16609 5825 16643
rect 5859 16609 5871 16643
rect 5813 16603 5871 16609
rect 5902 16600 5908 16652
rect 5960 16640 5966 16652
rect 6069 16643 6127 16649
rect 6069 16640 6081 16643
rect 5960 16612 6081 16640
rect 5960 16600 5966 16612
rect 6069 16609 6081 16612
rect 6115 16609 6127 16643
rect 6069 16603 6127 16609
rect 7006 16600 7012 16652
rect 7064 16640 7070 16652
rect 7285 16643 7343 16649
rect 7285 16640 7297 16643
rect 7064 16612 7297 16640
rect 7064 16600 7070 16612
rect 7285 16609 7297 16612
rect 7331 16609 7343 16643
rect 7285 16603 7343 16609
rect 7466 16600 7472 16652
rect 7524 16600 7530 16652
rect 7742 16600 7748 16652
rect 7800 16600 7806 16652
rect 7929 16643 7987 16649
rect 7929 16609 7941 16643
rect 7975 16609 7987 16643
rect 8036 16640 8064 16680
rect 8297 16677 8309 16711
rect 8343 16708 8355 16711
rect 8772 16708 8800 16748
rect 9030 16736 9036 16748
rect 9088 16736 9094 16788
rect 9950 16736 9956 16788
rect 10008 16776 10014 16788
rect 10689 16779 10747 16785
rect 10008 16748 10088 16776
rect 10008 16736 10014 16748
rect 8343 16680 8800 16708
rect 8849 16711 8907 16717
rect 8343 16677 8355 16680
rect 8297 16671 8355 16677
rect 8849 16677 8861 16711
rect 8895 16708 8907 16711
rect 8938 16708 8944 16720
rect 8895 16680 8944 16708
rect 8895 16677 8907 16680
rect 8849 16671 8907 16677
rect 8938 16668 8944 16680
rect 8996 16668 9002 16720
rect 9306 16649 9312 16652
rect 9033 16643 9091 16649
rect 9033 16640 9045 16643
rect 8036 16612 9045 16640
rect 7929 16603 7987 16609
rect 9033 16609 9045 16612
rect 9079 16609 9091 16643
rect 9300 16640 9312 16649
rect 9267 16612 9312 16640
rect 9033 16603 9091 16609
rect 9300 16603 9312 16612
rect 3436 16544 3536 16572
rect 4172 16544 4660 16572
rect 7484 16572 7512 16600
rect 7944 16572 7972 16603
rect 9306 16600 9312 16603
rect 9364 16600 9370 16652
rect 7484 16544 7972 16572
rect 8389 16575 8447 16581
rect 3053 16507 3111 16513
rect 3053 16473 3065 16507
rect 3099 16504 3111 16507
rect 3326 16504 3332 16516
rect 3099 16476 3332 16504
rect 3099 16473 3111 16476
rect 3053 16467 3111 16473
rect 3326 16464 3332 16476
rect 3384 16464 3390 16516
rect 3508 16504 3536 16544
rect 8389 16541 8401 16575
rect 8435 16572 8447 16575
rect 8478 16572 8484 16584
rect 8435 16544 8484 16572
rect 8435 16541 8447 16544
rect 8389 16535 8447 16541
rect 8478 16532 8484 16544
rect 8536 16532 8542 16584
rect 4798 16504 4804 16516
rect 3508 16476 4804 16504
rect 4798 16464 4804 16476
rect 4856 16464 4862 16516
rect 7742 16504 7748 16516
rect 6748 16476 7748 16504
rect 2740 16408 2820 16436
rect 2740 16396 2746 16408
rect 3786 16396 3792 16448
rect 3844 16436 3850 16448
rect 6454 16436 6460 16448
rect 3844 16408 6460 16436
rect 3844 16396 3850 16408
rect 6454 16396 6460 16408
rect 6512 16396 6518 16448
rect 6546 16396 6552 16448
rect 6604 16436 6610 16448
rect 6748 16436 6776 16476
rect 7742 16464 7748 16476
rect 7800 16464 7806 16516
rect 8849 16507 8907 16513
rect 8849 16473 8861 16507
rect 8895 16473 8907 16507
rect 8849 16467 8907 16473
rect 10060 16504 10088 16748
rect 10689 16745 10701 16779
rect 10735 16745 10747 16779
rect 10689 16739 10747 16745
rect 10704 16708 10732 16739
rect 12342 16736 12348 16788
rect 12400 16776 12406 16788
rect 12400 16748 13400 16776
rect 12400 16736 12406 16748
rect 10704 16680 12112 16708
rect 10594 16600 10600 16652
rect 10652 16600 10658 16652
rect 10778 16600 10784 16652
rect 10836 16600 10842 16652
rect 11072 16640 11100 16680
rect 11149 16643 11207 16649
rect 11149 16640 11161 16643
rect 11072 16612 11161 16640
rect 11149 16609 11161 16612
rect 11195 16609 11207 16643
rect 11149 16603 11207 16609
rect 11330 16600 11336 16652
rect 11388 16640 11394 16652
rect 11793 16643 11851 16649
rect 11793 16640 11805 16643
rect 11388 16612 11805 16640
rect 11388 16600 11394 16612
rect 11793 16609 11805 16612
rect 11839 16609 11851 16643
rect 11793 16603 11851 16609
rect 11974 16600 11980 16652
rect 12032 16600 12038 16652
rect 12084 16649 12112 16680
rect 12250 16668 12256 16720
rect 12308 16708 12314 16720
rect 13372 16708 13400 16748
rect 13722 16736 13728 16788
rect 13780 16776 13786 16788
rect 14366 16776 14372 16788
rect 13780 16748 14372 16776
rect 13780 16736 13786 16748
rect 14366 16736 14372 16748
rect 14424 16736 14430 16788
rect 14737 16779 14795 16785
rect 14737 16745 14749 16779
rect 14783 16776 14795 16779
rect 15470 16776 15476 16788
rect 14783 16748 15476 16776
rect 14783 16745 14795 16748
rect 14737 16739 14795 16745
rect 14918 16708 14924 16720
rect 12308 16680 12848 16708
rect 12308 16668 12314 16680
rect 12069 16643 12127 16649
rect 12069 16609 12081 16643
rect 12115 16609 12127 16643
rect 12069 16603 12127 16609
rect 12158 16600 12164 16652
rect 12216 16600 12222 16652
rect 12342 16600 12348 16652
rect 12400 16640 12406 16652
rect 12820 16649 12848 16680
rect 13372 16680 14924 16708
rect 12529 16643 12587 16649
rect 12400 16600 12434 16640
rect 12529 16609 12541 16643
rect 12575 16640 12587 16643
rect 12621 16643 12679 16649
rect 12621 16640 12633 16643
rect 12575 16612 12633 16640
rect 12575 16609 12587 16612
rect 12529 16603 12587 16609
rect 12621 16609 12633 16612
rect 12667 16609 12679 16643
rect 12621 16603 12679 16609
rect 12805 16643 12863 16649
rect 12805 16609 12817 16643
rect 12851 16609 12863 16643
rect 12805 16603 12863 16609
rect 12986 16600 12992 16652
rect 13044 16640 13050 16652
rect 13372 16649 13400 16680
rect 14918 16668 14924 16680
rect 14976 16668 14982 16720
rect 13081 16643 13139 16649
rect 13081 16640 13093 16643
rect 13044 16612 13093 16640
rect 13044 16600 13050 16612
rect 13081 16609 13093 16612
rect 13127 16609 13139 16643
rect 13081 16603 13139 16609
rect 13357 16643 13415 16649
rect 13357 16609 13369 16643
rect 13403 16609 13415 16643
rect 13357 16603 13415 16609
rect 13630 16600 13636 16652
rect 13688 16600 13694 16652
rect 13998 16600 14004 16652
rect 14056 16640 14062 16652
rect 14550 16640 14556 16652
rect 14056 16612 14556 16640
rect 14056 16600 14062 16612
rect 14550 16600 14556 16612
rect 14608 16600 14614 16652
rect 14737 16643 14795 16649
rect 14737 16609 14749 16643
rect 14783 16640 14795 16643
rect 14826 16640 14832 16652
rect 14783 16612 14832 16640
rect 14783 16609 14795 16612
rect 14737 16603 14795 16609
rect 14826 16600 14832 16612
rect 14884 16600 14890 16652
rect 15028 16649 15056 16748
rect 15470 16736 15476 16748
rect 15528 16736 15534 16788
rect 16294 16779 16352 16785
rect 16294 16776 16306 16779
rect 15764 16748 16306 16776
rect 15764 16708 15792 16748
rect 16294 16745 16306 16748
rect 16340 16745 16352 16779
rect 16294 16739 16352 16745
rect 17957 16779 18015 16785
rect 17957 16745 17969 16779
rect 18003 16776 18015 16779
rect 18414 16776 18420 16788
rect 18003 16748 18420 16776
rect 18003 16745 18015 16748
rect 17957 16739 18015 16745
rect 15212 16680 15792 16708
rect 16393 16711 16451 16717
rect 15212 16649 15240 16680
rect 15013 16643 15071 16649
rect 15013 16609 15025 16643
rect 15059 16609 15071 16643
rect 15013 16603 15071 16609
rect 15197 16643 15255 16649
rect 15197 16609 15209 16643
rect 15243 16609 15255 16643
rect 15197 16603 15255 16609
rect 15289 16643 15347 16649
rect 15289 16609 15301 16643
rect 15335 16640 15347 16643
rect 15562 16640 15568 16652
rect 15335 16612 15568 16640
rect 15335 16609 15347 16612
rect 15289 16603 15347 16609
rect 15562 16600 15568 16612
rect 15620 16600 15626 16652
rect 10134 16532 10140 16584
rect 10192 16572 10198 16584
rect 10686 16572 10692 16584
rect 10192 16544 10692 16572
rect 10192 16532 10198 16544
rect 10686 16532 10692 16544
rect 10744 16532 10750 16584
rect 11057 16575 11115 16581
rect 11057 16541 11069 16575
rect 11103 16572 11115 16575
rect 11992 16572 12020 16600
rect 11103 16544 12020 16572
rect 12406 16572 12434 16600
rect 13262 16572 13268 16584
rect 12406 16544 13268 16572
rect 11103 16541 11115 16544
rect 11057 16535 11115 16541
rect 13262 16532 13268 16544
rect 13320 16572 13326 16584
rect 13722 16572 13728 16584
rect 13320 16544 13728 16572
rect 13320 16532 13326 16544
rect 13722 16532 13728 16544
rect 13780 16532 13786 16584
rect 15672 16581 15700 16680
rect 16393 16677 16405 16711
rect 16439 16708 16451 16711
rect 16758 16708 16764 16720
rect 16439 16680 16764 16708
rect 16439 16677 16451 16680
rect 16393 16671 16451 16677
rect 16758 16668 16764 16680
rect 16816 16708 16822 16720
rect 17126 16708 17132 16720
rect 16816 16680 17132 16708
rect 16816 16668 16822 16680
rect 17126 16668 17132 16680
rect 17184 16668 17190 16720
rect 17420 16680 17816 16708
rect 17420 16652 17448 16680
rect 15930 16600 15936 16652
rect 15988 16640 15994 16652
rect 16117 16643 16175 16649
rect 16117 16640 16129 16643
rect 15988 16612 16129 16640
rect 15988 16600 15994 16612
rect 16117 16609 16129 16612
rect 16163 16609 16175 16643
rect 16117 16603 16175 16609
rect 16206 16600 16212 16652
rect 16264 16600 16270 16652
rect 17034 16600 17040 16652
rect 17092 16600 17098 16652
rect 17218 16600 17224 16652
rect 17276 16640 17282 16652
rect 17276 16612 17356 16640
rect 17276 16600 17282 16612
rect 15657 16575 15715 16581
rect 15657 16541 15669 16575
rect 15703 16541 15715 16575
rect 17328 16572 17356 16612
rect 17402 16600 17408 16652
rect 17460 16600 17466 16652
rect 17788 16649 17816 16680
rect 17497 16643 17555 16649
rect 17497 16609 17509 16643
rect 17543 16609 17555 16643
rect 17497 16603 17555 16609
rect 17681 16643 17739 16649
rect 17681 16609 17693 16643
rect 17727 16609 17739 16643
rect 17681 16603 17739 16609
rect 17773 16643 17831 16649
rect 17773 16609 17785 16643
rect 17819 16609 17831 16643
rect 17773 16603 17831 16609
rect 17512 16572 17540 16603
rect 17328 16544 17540 16572
rect 17696 16572 17724 16603
rect 17972 16572 18000 16739
rect 18414 16736 18420 16748
rect 18472 16736 18478 16788
rect 20717 16779 20775 16785
rect 20717 16776 20729 16779
rect 18616 16748 20729 16776
rect 18616 16581 18644 16748
rect 18874 16708 18880 16720
rect 18708 16680 18880 16708
rect 18708 16649 18736 16680
rect 18874 16668 18880 16680
rect 18932 16708 18938 16720
rect 18932 16680 19196 16708
rect 18932 16668 18938 16680
rect 18693 16643 18751 16649
rect 18693 16609 18705 16643
rect 18739 16609 18751 16643
rect 18693 16603 18751 16609
rect 18782 16600 18788 16652
rect 18840 16640 18846 16652
rect 19168 16649 19196 16680
rect 19352 16649 19380 16748
rect 20717 16745 20729 16748
rect 20763 16745 20775 16779
rect 20717 16739 20775 16745
rect 21082 16736 21088 16788
rect 21140 16736 21146 16788
rect 21174 16736 21180 16788
rect 21232 16776 21238 16788
rect 21453 16779 21511 16785
rect 21453 16776 21465 16779
rect 21232 16748 21465 16776
rect 21232 16736 21238 16748
rect 21453 16745 21465 16748
rect 21499 16745 21511 16779
rect 21453 16739 21511 16745
rect 22186 16736 22192 16788
rect 22244 16776 22250 16788
rect 22738 16776 22744 16788
rect 22244 16748 22744 16776
rect 22244 16736 22250 16748
rect 22738 16736 22744 16748
rect 22796 16736 22802 16788
rect 23017 16779 23075 16785
rect 23017 16745 23029 16779
rect 23063 16776 23075 16779
rect 23198 16776 23204 16788
rect 23063 16748 23204 16776
rect 23063 16745 23075 16748
rect 23017 16739 23075 16745
rect 23198 16736 23204 16748
rect 23256 16736 23262 16788
rect 19886 16668 19892 16720
rect 19944 16668 19950 16720
rect 20070 16668 20076 16720
rect 20128 16708 20134 16720
rect 21100 16708 21128 16736
rect 20128 16680 20944 16708
rect 21100 16680 21947 16708
rect 20128 16668 20134 16680
rect 18969 16643 19027 16649
rect 18969 16640 18981 16643
rect 18840 16612 18981 16640
rect 18840 16600 18846 16612
rect 18969 16609 18981 16612
rect 19015 16609 19027 16643
rect 18969 16603 19027 16609
rect 19153 16643 19211 16649
rect 19153 16609 19165 16643
rect 19199 16609 19211 16643
rect 19153 16603 19211 16609
rect 19337 16643 19395 16649
rect 19337 16609 19349 16643
rect 19383 16609 19395 16643
rect 19904 16640 19932 16668
rect 20349 16643 20407 16649
rect 20349 16640 20361 16643
rect 19904 16612 20361 16640
rect 19337 16603 19395 16609
rect 20349 16609 20361 16612
rect 20395 16609 20407 16643
rect 20349 16603 20407 16609
rect 20533 16643 20591 16649
rect 20533 16609 20545 16643
rect 20579 16609 20591 16643
rect 20533 16603 20591 16609
rect 20625 16643 20683 16649
rect 20625 16609 20637 16643
rect 20671 16640 20683 16643
rect 20714 16640 20720 16652
rect 20671 16612 20720 16640
rect 20671 16609 20683 16612
rect 20625 16603 20683 16609
rect 17696 16544 18000 16572
rect 18601 16575 18659 16581
rect 15657 16535 15715 16541
rect 18601 16541 18613 16575
rect 18647 16541 18659 16575
rect 18601 16535 18659 16541
rect 12802 16504 12808 16516
rect 10060 16476 12434 16504
rect 6604 16408 6776 16436
rect 6604 16396 6610 16408
rect 7098 16396 7104 16448
rect 7156 16436 7162 16448
rect 7193 16439 7251 16445
rect 7193 16436 7205 16439
rect 7156 16408 7205 16436
rect 7156 16396 7162 16408
rect 7193 16405 7205 16408
rect 7239 16405 7251 16439
rect 8864 16436 8892 16467
rect 9674 16436 9680 16448
rect 8864 16408 9680 16436
rect 7193 16399 7251 16405
rect 9674 16396 9680 16408
rect 9732 16436 9738 16448
rect 10060 16436 10088 16476
rect 9732 16408 10088 16436
rect 9732 16396 9738 16408
rect 10410 16396 10416 16448
rect 10468 16436 10474 16448
rect 10962 16436 10968 16448
rect 10468 16408 10968 16436
rect 10468 16396 10474 16408
rect 10962 16396 10968 16408
rect 11020 16396 11026 16448
rect 11514 16396 11520 16448
rect 11572 16396 11578 16448
rect 11606 16396 11612 16448
rect 11664 16396 11670 16448
rect 11974 16396 11980 16448
rect 12032 16436 12038 16448
rect 12158 16436 12164 16448
rect 12032 16408 12164 16436
rect 12032 16396 12038 16408
rect 12158 16396 12164 16408
rect 12216 16396 12222 16448
rect 12406 16436 12434 16476
rect 12636 16476 12808 16504
rect 12636 16436 12664 16476
rect 12802 16464 12808 16476
rect 12860 16464 12866 16516
rect 12894 16464 12900 16516
rect 12952 16464 12958 16516
rect 12986 16464 12992 16516
rect 13044 16504 13050 16516
rect 14829 16507 14887 16513
rect 14829 16504 14841 16507
rect 13044 16476 14841 16504
rect 13044 16464 13050 16476
rect 14829 16473 14841 16476
rect 14875 16473 14887 16507
rect 14829 16467 14887 16473
rect 18322 16464 18328 16516
rect 18380 16464 18386 16516
rect 18506 16464 18512 16516
rect 18564 16504 18570 16516
rect 19150 16504 19156 16516
rect 18564 16476 19156 16504
rect 18564 16464 18570 16476
rect 19150 16464 19156 16476
rect 19208 16464 19214 16516
rect 20556 16504 20584 16603
rect 20714 16600 20720 16612
rect 20772 16600 20778 16652
rect 20916 16649 20944 16680
rect 20809 16643 20867 16649
rect 20809 16609 20821 16643
rect 20855 16609 20867 16643
rect 20809 16603 20867 16609
rect 20901 16643 20959 16649
rect 20901 16609 20913 16643
rect 20947 16609 20959 16643
rect 20901 16603 20959 16609
rect 20824 16572 20852 16603
rect 21082 16600 21088 16652
rect 21140 16640 21146 16652
rect 21269 16643 21327 16649
rect 21269 16640 21281 16643
rect 21140 16612 21281 16640
rect 21140 16600 21146 16612
rect 21269 16609 21281 16612
rect 21315 16609 21327 16643
rect 21269 16603 21327 16609
rect 21637 16643 21695 16649
rect 21637 16609 21649 16643
rect 21683 16640 21695 16643
rect 21726 16640 21732 16652
rect 21683 16612 21732 16640
rect 21683 16609 21695 16612
rect 21637 16603 21695 16609
rect 21726 16600 21732 16612
rect 21784 16600 21790 16652
rect 21919 16649 21947 16680
rect 21904 16643 21962 16649
rect 21904 16609 21916 16643
rect 21950 16640 21962 16643
rect 22370 16640 22376 16652
rect 21950 16612 22376 16640
rect 21950 16609 21962 16612
rect 21904 16603 21962 16609
rect 22370 16600 22376 16612
rect 22428 16600 22434 16652
rect 21100 16572 21128 16600
rect 20824 16544 21128 16572
rect 20824 16504 20852 16544
rect 20556 16476 20852 16504
rect 12406 16408 12664 16436
rect 12710 16396 12716 16448
rect 12768 16396 12774 16448
rect 13078 16396 13084 16448
rect 13136 16436 13142 16448
rect 13173 16439 13231 16445
rect 13173 16436 13185 16439
rect 13136 16408 13185 16436
rect 13136 16396 13142 16408
rect 13173 16405 13185 16408
rect 13219 16405 13231 16439
rect 13173 16399 13231 16405
rect 13354 16396 13360 16448
rect 13412 16436 13418 16448
rect 13449 16439 13507 16445
rect 13449 16436 13461 16439
rect 13412 16408 13461 16436
rect 13412 16396 13418 16408
rect 13449 16405 13461 16408
rect 13495 16405 13507 16439
rect 13449 16399 13507 16405
rect 15930 16396 15936 16448
rect 15988 16396 15994 16448
rect 17494 16396 17500 16448
rect 17552 16396 17558 16448
rect 19058 16396 19064 16448
rect 19116 16396 19122 16448
rect 20070 16396 20076 16448
rect 20128 16436 20134 16448
rect 20257 16439 20315 16445
rect 20257 16436 20269 16439
rect 20128 16408 20269 16436
rect 20128 16396 20134 16408
rect 20257 16405 20269 16408
rect 20303 16405 20315 16439
rect 20257 16399 20315 16405
rect 20438 16396 20444 16448
rect 20496 16396 20502 16448
rect 21082 16396 21088 16448
rect 21140 16396 21146 16448
rect 552 16346 23368 16368
rect 552 16294 1366 16346
rect 1418 16294 1430 16346
rect 1482 16294 1494 16346
rect 1546 16294 1558 16346
rect 1610 16294 1622 16346
rect 1674 16294 1686 16346
rect 1738 16294 7366 16346
rect 7418 16294 7430 16346
rect 7482 16294 7494 16346
rect 7546 16294 7558 16346
rect 7610 16294 7622 16346
rect 7674 16294 7686 16346
rect 7738 16294 13366 16346
rect 13418 16294 13430 16346
rect 13482 16294 13494 16346
rect 13546 16294 13558 16346
rect 13610 16294 13622 16346
rect 13674 16294 13686 16346
rect 13738 16294 19366 16346
rect 19418 16294 19430 16346
rect 19482 16294 19494 16346
rect 19546 16294 19558 16346
rect 19610 16294 19622 16346
rect 19674 16294 19686 16346
rect 19738 16294 23368 16346
rect 552 16272 23368 16294
rect 2314 16192 2320 16244
rect 2372 16232 2378 16244
rect 4982 16232 4988 16244
rect 2372 16204 4988 16232
rect 2372 16192 2378 16204
rect 4982 16192 4988 16204
rect 5040 16192 5046 16244
rect 5442 16192 5448 16244
rect 5500 16232 5506 16244
rect 6181 16235 6239 16241
rect 6181 16232 6193 16235
rect 5500 16204 6193 16232
rect 5500 16192 5506 16204
rect 6181 16201 6193 16204
rect 6227 16201 6239 16235
rect 6181 16195 6239 16201
rect 7745 16235 7803 16241
rect 7745 16201 7757 16235
rect 7791 16232 7803 16235
rect 8202 16232 8208 16244
rect 7791 16204 8208 16232
rect 7791 16201 7803 16204
rect 7745 16195 7803 16201
rect 8202 16192 8208 16204
rect 8260 16192 8266 16244
rect 8389 16235 8447 16241
rect 8389 16201 8401 16235
rect 8435 16232 8447 16235
rect 8478 16232 8484 16244
rect 8435 16204 8484 16232
rect 8435 16201 8447 16204
rect 8389 16195 8447 16201
rect 8478 16192 8484 16204
rect 8536 16192 8542 16244
rect 8754 16192 8760 16244
rect 8812 16192 8818 16244
rect 9674 16232 9680 16244
rect 9416 16204 9680 16232
rect 2225 16167 2283 16173
rect 2225 16133 2237 16167
rect 2271 16164 2283 16167
rect 2866 16164 2872 16176
rect 2271 16136 2872 16164
rect 2271 16133 2283 16136
rect 2225 16127 2283 16133
rect 2866 16124 2872 16136
rect 2924 16124 2930 16176
rect 5626 16124 5632 16176
rect 5684 16164 5690 16176
rect 6457 16167 6515 16173
rect 6457 16164 6469 16167
rect 5684 16136 6469 16164
rect 5684 16124 5690 16136
rect 6457 16133 6469 16136
rect 6503 16164 6515 16167
rect 6822 16164 6828 16176
rect 6503 16136 6828 16164
rect 6503 16133 6515 16136
rect 6457 16127 6515 16133
rect 6822 16124 6828 16136
rect 6880 16164 6886 16176
rect 6880 16136 7144 16164
rect 6880 16124 6886 16136
rect 842 16056 848 16108
rect 900 16056 906 16108
rect 2682 16056 2688 16108
rect 2740 16096 2746 16108
rect 3050 16096 3056 16108
rect 2740 16068 3056 16096
rect 2740 16056 2746 16068
rect 3050 16056 3056 16068
rect 3108 16056 3114 16108
rect 4890 16056 4896 16108
rect 4948 16056 4954 16108
rect 5718 16056 5724 16108
rect 5776 16056 5782 16108
rect 5813 16099 5871 16105
rect 5813 16065 5825 16099
rect 5859 16096 5871 16099
rect 6089 16099 6147 16105
rect 5859 16068 6040 16096
rect 5859 16065 5871 16068
rect 5813 16059 5871 16065
rect 1118 16037 1124 16040
rect 1112 16028 1124 16037
rect 1079 16000 1124 16028
rect 1112 15991 1124 16000
rect 1118 15988 1124 15991
rect 1176 15988 1182 16040
rect 2409 16031 2467 16037
rect 2409 15997 2421 16031
rect 2455 15997 2467 16031
rect 2409 15991 2467 15997
rect 2424 15960 2452 15991
rect 2774 15988 2780 16040
rect 2832 16028 2838 16040
rect 2869 16031 2927 16037
rect 2869 16028 2881 16031
rect 2832 16000 2881 16028
rect 2832 15988 2838 16000
rect 2869 15997 2881 16000
rect 2915 15997 2927 16031
rect 2869 15991 2927 15997
rect 3234 15988 3240 16040
rect 3292 15988 3298 16040
rect 3326 15988 3332 16040
rect 3384 16028 3390 16040
rect 3493 16031 3551 16037
rect 3493 16028 3505 16031
rect 3384 16000 3505 16028
rect 3384 15988 3390 16000
rect 3493 15997 3505 16000
rect 3539 15997 3551 16031
rect 3493 15991 3551 15997
rect 4982 15988 4988 16040
rect 5040 16028 5046 16040
rect 5629 16031 5687 16037
rect 5629 16028 5641 16031
rect 5040 16000 5641 16028
rect 5040 15988 5046 16000
rect 5629 15997 5641 16000
rect 5675 15997 5687 16031
rect 5629 15991 5687 15997
rect 5905 16031 5963 16037
rect 5905 15997 5917 16031
rect 5951 15997 5963 16031
rect 6012 16028 6040 16068
rect 6089 16065 6101 16099
rect 6135 16096 6147 16099
rect 6135 16068 6684 16096
rect 6135 16065 6147 16068
rect 6089 16059 6147 16065
rect 6178 16028 6184 16040
rect 6012 16000 6184 16028
rect 5905 15991 5963 15997
rect 2424 15932 4660 15960
rect 2498 15852 2504 15904
rect 2556 15892 2562 15904
rect 2593 15895 2651 15901
rect 2593 15892 2605 15895
rect 2556 15864 2605 15892
rect 2556 15852 2562 15864
rect 2593 15861 2605 15864
rect 2639 15861 2651 15895
rect 2593 15855 2651 15861
rect 2685 15895 2743 15901
rect 2685 15861 2697 15895
rect 2731 15892 2743 15895
rect 2774 15892 2780 15904
rect 2731 15864 2780 15892
rect 2731 15861 2743 15864
rect 2685 15855 2743 15861
rect 2774 15852 2780 15864
rect 2832 15852 2838 15904
rect 4632 15901 4660 15932
rect 4798 15920 4804 15972
rect 4856 15960 4862 15972
rect 5920 15960 5948 15991
rect 6178 15988 6184 16000
rect 6236 15988 6242 16040
rect 6365 16031 6423 16037
rect 6365 16028 6377 16031
rect 6288 16000 6377 16028
rect 4856 15932 5948 15960
rect 4856 15920 4862 15932
rect 4617 15895 4675 15901
rect 4617 15861 4629 15895
rect 4663 15892 4675 15895
rect 4982 15892 4988 15904
rect 4663 15864 4988 15892
rect 4663 15861 4675 15864
rect 4617 15855 4675 15861
rect 4982 15852 4988 15864
rect 5040 15852 5046 15904
rect 5077 15895 5135 15901
rect 5077 15861 5089 15895
rect 5123 15892 5135 15895
rect 5258 15892 5264 15904
rect 5123 15864 5264 15892
rect 5123 15861 5135 15864
rect 5077 15855 5135 15861
rect 5258 15852 5264 15864
rect 5316 15852 5322 15904
rect 5442 15852 5448 15904
rect 5500 15852 5506 15904
rect 5718 15852 5724 15904
rect 5776 15892 5782 15904
rect 6288 15892 6316 16000
rect 6365 15997 6377 16000
rect 6411 15997 6423 16031
rect 6365 15991 6423 15997
rect 6546 15988 6552 16040
rect 6604 15988 6610 16040
rect 6656 16037 6684 16068
rect 6730 16056 6736 16108
rect 6788 16096 6794 16108
rect 7116 16105 7144 16136
rect 7101 16099 7159 16105
rect 6788 16068 7052 16096
rect 6788 16056 6794 16068
rect 6641 16031 6699 16037
rect 6641 15997 6653 16031
rect 6687 15997 6699 16031
rect 6641 15991 6699 15997
rect 6825 16031 6883 16037
rect 6825 15997 6837 16031
rect 6871 16028 6883 16031
rect 6914 16028 6920 16040
rect 6871 16000 6920 16028
rect 6871 15997 6883 16000
rect 6825 15991 6883 15997
rect 6454 15920 6460 15972
rect 6512 15960 6518 15972
rect 6840 15960 6868 15991
rect 6914 15988 6920 16000
rect 6972 15988 6978 16040
rect 7024 16037 7052 16068
rect 7101 16065 7113 16099
rect 7147 16065 7159 16099
rect 7101 16059 7159 16065
rect 7190 16056 7196 16108
rect 7248 16096 7254 16108
rect 7377 16099 7435 16105
rect 7377 16096 7389 16099
rect 7248 16068 7389 16096
rect 7248 16056 7254 16068
rect 7377 16065 7389 16068
rect 7423 16065 7435 16099
rect 7377 16059 7435 16065
rect 9125 16099 9183 16105
rect 9125 16065 9137 16099
rect 9171 16096 9183 16099
rect 9416 16096 9444 16204
rect 9674 16192 9680 16204
rect 9732 16192 9738 16244
rect 9861 16235 9919 16241
rect 9861 16201 9873 16235
rect 9907 16232 9919 16235
rect 9950 16232 9956 16244
rect 9907 16204 9956 16232
rect 9907 16201 9919 16204
rect 9861 16195 9919 16201
rect 9950 16192 9956 16204
rect 10008 16192 10014 16244
rect 10594 16192 10600 16244
rect 10652 16232 10658 16244
rect 10689 16235 10747 16241
rect 10689 16232 10701 16235
rect 10652 16204 10701 16232
rect 10652 16192 10658 16204
rect 10689 16201 10701 16204
rect 10735 16201 10747 16235
rect 10689 16195 10747 16201
rect 10778 16192 10784 16244
rect 10836 16232 10842 16244
rect 10873 16235 10931 16241
rect 10873 16232 10885 16235
rect 10836 16204 10885 16232
rect 10836 16192 10842 16204
rect 10873 16201 10885 16204
rect 10919 16201 10931 16235
rect 10873 16195 10931 16201
rect 11885 16235 11943 16241
rect 11885 16201 11897 16235
rect 11931 16232 11943 16235
rect 12250 16232 12256 16244
rect 11931 16204 12256 16232
rect 11931 16201 11943 16204
rect 11885 16195 11943 16201
rect 12250 16192 12256 16204
rect 12308 16192 12314 16244
rect 15654 16192 15660 16244
rect 15712 16232 15718 16244
rect 16206 16232 16212 16244
rect 15712 16204 16212 16232
rect 15712 16192 15718 16204
rect 16206 16192 16212 16204
rect 16264 16232 16270 16244
rect 16485 16235 16543 16241
rect 16485 16232 16497 16235
rect 16264 16204 16497 16232
rect 16264 16192 16270 16204
rect 16485 16201 16497 16204
rect 16531 16232 16543 16235
rect 18230 16232 18236 16244
rect 16531 16204 18236 16232
rect 16531 16201 16543 16204
rect 16485 16195 16543 16201
rect 18230 16192 18236 16204
rect 18288 16192 18294 16244
rect 21174 16232 21180 16244
rect 18340 16204 21180 16232
rect 9766 16164 9772 16176
rect 9508 16136 9772 16164
rect 9508 16105 9536 16136
rect 9766 16124 9772 16136
rect 9824 16164 9830 16176
rect 14093 16167 14151 16173
rect 14093 16164 14105 16167
rect 9824 16136 14105 16164
rect 9824 16124 9830 16136
rect 14093 16133 14105 16136
rect 14139 16133 14151 16167
rect 14093 16127 14151 16133
rect 17954 16124 17960 16176
rect 18012 16164 18018 16176
rect 18340 16164 18368 16204
rect 21174 16192 21180 16204
rect 21232 16192 21238 16244
rect 22097 16235 22155 16241
rect 22097 16201 22109 16235
rect 22143 16232 22155 16235
rect 22278 16232 22284 16244
rect 22143 16204 22284 16232
rect 22143 16201 22155 16204
rect 22097 16195 22155 16201
rect 22278 16192 22284 16204
rect 22336 16192 22342 16244
rect 22833 16235 22891 16241
rect 22833 16201 22845 16235
rect 22879 16232 22891 16235
rect 22922 16232 22928 16244
rect 22879 16204 22928 16232
rect 22879 16201 22891 16204
rect 22833 16195 22891 16201
rect 22922 16192 22928 16204
rect 22980 16192 22986 16244
rect 18012 16136 18368 16164
rect 18012 16124 18018 16136
rect 20254 16124 20260 16176
rect 20312 16164 20318 16176
rect 20990 16164 20996 16176
rect 20312 16136 20996 16164
rect 20312 16124 20318 16136
rect 20990 16124 20996 16136
rect 21048 16124 21054 16176
rect 21266 16124 21272 16176
rect 21324 16164 21330 16176
rect 21821 16167 21879 16173
rect 21821 16164 21833 16167
rect 21324 16136 21833 16164
rect 21324 16124 21330 16136
rect 21821 16133 21833 16136
rect 21867 16133 21879 16167
rect 21821 16127 21879 16133
rect 9171 16068 9444 16096
rect 9493 16099 9551 16105
rect 9171 16065 9183 16068
rect 9125 16059 9183 16065
rect 9493 16065 9505 16099
rect 9539 16065 9551 16099
rect 10137 16099 10195 16105
rect 10137 16096 10149 16099
rect 9493 16059 9551 16065
rect 9600 16068 10149 16096
rect 7009 16031 7067 16037
rect 7009 15997 7021 16031
rect 7055 15997 7067 16031
rect 7009 15991 7067 15997
rect 7834 15988 7840 16040
rect 7892 16028 7898 16040
rect 8021 16031 8079 16037
rect 8021 16028 8033 16031
rect 7892 16000 8033 16028
rect 7892 15988 7898 16000
rect 8021 15997 8033 16000
rect 8067 15997 8079 16031
rect 8021 15991 8079 15997
rect 8202 15988 8208 16040
rect 8260 15988 8266 16040
rect 8573 16031 8631 16037
rect 8573 15997 8585 16031
rect 8619 15997 8631 16031
rect 8573 15991 8631 15997
rect 8941 16031 8999 16037
rect 8941 15997 8953 16031
rect 8987 15997 8999 16031
rect 8941 15991 8999 15997
rect 6512 15932 6868 15960
rect 6512 15920 6518 15932
rect 7190 15920 7196 15972
rect 7248 15960 7254 15972
rect 7469 15963 7527 15969
rect 7469 15960 7481 15963
rect 7248 15932 7481 15960
rect 7248 15920 7254 15932
rect 7469 15929 7481 15932
rect 7515 15929 7527 15963
rect 7469 15923 7527 15929
rect 7586 15963 7644 15969
rect 7586 15929 7598 15963
rect 7632 15929 7644 15963
rect 8588 15960 8616 15991
rect 7586 15923 7644 15929
rect 7852 15932 8616 15960
rect 8956 15960 8984 15991
rect 9030 15988 9036 16040
rect 9088 15988 9094 16040
rect 9600 16037 9628 16068
rect 10137 16065 10149 16068
rect 10183 16065 10195 16099
rect 10410 16096 10416 16108
rect 10137 16059 10195 16065
rect 10336 16068 10416 16096
rect 9217 16031 9275 16037
rect 9217 15997 9229 16031
rect 9263 15997 9275 16031
rect 9217 15991 9275 15997
rect 9585 16031 9643 16037
rect 9585 15997 9597 16031
rect 9631 16028 9643 16031
rect 9674 16028 9680 16040
rect 9631 16000 9680 16028
rect 9631 15997 9643 16000
rect 9585 15991 9643 15997
rect 9122 15960 9128 15972
rect 8956 15932 9128 15960
rect 5776 15864 6316 15892
rect 6917 15895 6975 15901
rect 5776 15852 5782 15864
rect 6917 15861 6929 15895
rect 6963 15892 6975 15895
rect 7282 15892 7288 15904
rect 6963 15864 7288 15892
rect 6963 15861 6975 15864
rect 6917 15855 6975 15861
rect 7282 15852 7288 15864
rect 7340 15852 7346 15904
rect 7601 15892 7629 15923
rect 7852 15904 7880 15932
rect 9122 15920 9128 15932
rect 9180 15920 9186 15972
rect 9232 15960 9260 15991
rect 9674 15988 9680 16000
rect 9732 15988 9738 16040
rect 10042 15988 10048 16040
rect 10100 15988 10106 16040
rect 10226 15988 10232 16040
rect 10284 15988 10290 16040
rect 10336 16037 10364 16068
rect 10410 16056 10416 16068
rect 10468 16056 10474 16108
rect 12250 16096 12256 16108
rect 10612 16068 11100 16096
rect 10612 16037 10640 16068
rect 11072 16037 11100 16068
rect 11164 16068 11836 16096
rect 10321 16031 10379 16037
rect 10321 15997 10333 16031
rect 10367 15997 10379 16031
rect 10597 16031 10655 16037
rect 10597 16028 10609 16031
rect 10321 15991 10379 15997
rect 10428 16000 10609 16028
rect 10134 15960 10140 15972
rect 9232 15932 10140 15960
rect 10134 15920 10140 15932
rect 10192 15920 10198 15972
rect 7834 15892 7840 15904
rect 7601 15864 7840 15892
rect 7834 15852 7840 15864
rect 7892 15852 7898 15904
rect 8018 15852 8024 15904
rect 8076 15852 8082 15904
rect 8662 15852 8668 15904
rect 8720 15892 8726 15904
rect 9398 15892 9404 15904
rect 8720 15864 9404 15892
rect 8720 15852 8726 15864
rect 9398 15852 9404 15864
rect 9456 15892 9462 15904
rect 10428 15892 10456 16000
rect 10597 15997 10609 16000
rect 10643 15997 10655 16031
rect 10597 15991 10655 15997
rect 10774 16031 10832 16037
rect 10774 15997 10786 16031
rect 10820 15997 10832 16031
rect 10774 15991 10832 15997
rect 11057 16031 11115 16037
rect 11057 15997 11069 16031
rect 11103 15997 11115 16031
rect 11057 15991 11115 15997
rect 10796 15960 10824 15991
rect 11164 15960 11192 16068
rect 11808 16040 11836 16068
rect 11900 16068 12256 16096
rect 11241 16031 11299 16037
rect 11241 15997 11253 16031
rect 11287 16028 11299 16031
rect 11517 16031 11575 16037
rect 11517 16028 11529 16031
rect 11287 16000 11529 16028
rect 11287 15997 11299 16000
rect 11241 15991 11299 15997
rect 11517 15997 11529 16000
rect 11563 15997 11575 16031
rect 11517 15991 11575 15997
rect 10796 15932 11192 15960
rect 9456 15864 10456 15892
rect 10505 15895 10563 15901
rect 9456 15852 9462 15864
rect 10505 15861 10517 15895
rect 10551 15892 10563 15895
rect 11256 15892 11284 15991
rect 10551 15864 11284 15892
rect 10551 15861 10563 15864
rect 10505 15855 10563 15861
rect 11330 15852 11336 15904
rect 11388 15852 11394 15904
rect 11532 15892 11560 15991
rect 11790 15988 11796 16040
rect 11848 15988 11854 16040
rect 11900 15960 11928 16068
rect 12250 16056 12256 16068
rect 12308 16056 12314 16108
rect 12621 16099 12679 16105
rect 12621 16065 12633 16099
rect 12667 16096 12679 16099
rect 12710 16096 12716 16108
rect 12667 16068 12716 16096
rect 12667 16065 12679 16068
rect 12621 16059 12679 16065
rect 12710 16056 12716 16068
rect 12768 16096 12774 16108
rect 12768 16068 12940 16096
rect 12768 16056 12774 16068
rect 11977 16031 12035 16037
rect 11977 15997 11989 16031
rect 12023 16028 12035 16031
rect 12342 16028 12348 16040
rect 12023 16000 12348 16028
rect 12023 15997 12035 16000
rect 11977 15991 12035 15997
rect 12342 15988 12348 16000
rect 12400 15988 12406 16040
rect 12912 16037 12940 16068
rect 12986 16056 12992 16108
rect 13044 16056 13050 16108
rect 13078 16056 13084 16108
rect 13136 16096 13142 16108
rect 13265 16099 13323 16105
rect 13265 16096 13277 16099
rect 13136 16068 13277 16096
rect 13136 16056 13142 16068
rect 13265 16065 13277 16068
rect 13311 16065 13323 16099
rect 14461 16099 14519 16105
rect 13265 16059 13323 16065
rect 13556 16068 14412 16096
rect 12437 16031 12495 16037
rect 12437 15997 12449 16031
rect 12483 15997 12495 16031
rect 12437 15991 12495 15997
rect 12897 16031 12955 16037
rect 12897 15997 12909 16031
rect 12943 15997 12955 16031
rect 12897 15991 12955 15997
rect 12069 15963 12127 15969
rect 12069 15960 12081 15963
rect 11900 15932 12081 15960
rect 12069 15929 12081 15932
rect 12115 15929 12127 15963
rect 12069 15923 12127 15929
rect 12161 15963 12219 15969
rect 12161 15929 12173 15963
rect 12207 15960 12219 15963
rect 12250 15960 12256 15972
rect 12207 15932 12256 15960
rect 12207 15929 12219 15932
rect 12161 15923 12219 15929
rect 12250 15920 12256 15932
rect 12308 15920 12314 15972
rect 12452 15960 12480 15991
rect 13004 15960 13032 16056
rect 13556 16040 13584 16068
rect 13538 15988 13544 16040
rect 13596 15988 13602 16040
rect 14384 16037 14412 16068
rect 14461 16065 14473 16099
rect 14507 16096 14519 16099
rect 14921 16099 14979 16105
rect 14921 16096 14933 16099
rect 14507 16068 14933 16096
rect 14507 16065 14519 16068
rect 14461 16059 14519 16065
rect 14921 16065 14933 16068
rect 14967 16096 14979 16099
rect 19058 16096 19064 16108
rect 14967 16068 19064 16096
rect 14967 16065 14979 16068
rect 14921 16059 14979 16065
rect 19058 16056 19064 16068
rect 19116 16056 19122 16108
rect 21836 16096 21864 16127
rect 22002 16124 22008 16176
rect 22060 16164 22066 16176
rect 22465 16167 22523 16173
rect 22465 16164 22477 16167
rect 22060 16136 22477 16164
rect 22060 16124 22066 16136
rect 22465 16133 22477 16136
rect 22511 16133 22523 16167
rect 22465 16127 22523 16133
rect 22094 16096 22100 16108
rect 21376 16068 21680 16096
rect 21836 16068 22100 16096
rect 21376 16040 21404 16068
rect 13725 16031 13783 16037
rect 13725 15997 13737 16031
rect 13771 15997 13783 16031
rect 13725 15991 13783 15997
rect 14369 16031 14427 16037
rect 14369 15997 14381 16031
rect 14415 15997 14427 16031
rect 14369 15991 14427 15997
rect 14829 16031 14887 16037
rect 14829 15997 14841 16031
rect 14875 15997 14887 16031
rect 14829 15991 14887 15997
rect 16393 16031 16451 16037
rect 16393 15997 16405 16031
rect 16439 16028 16451 16031
rect 16669 16031 16727 16037
rect 16669 16028 16681 16031
rect 16439 16000 16681 16028
rect 16439 15997 16451 16000
rect 16393 15991 16451 15997
rect 16669 15997 16681 16000
rect 16715 16028 16727 16031
rect 16942 16028 16948 16040
rect 16715 16000 16948 16028
rect 16715 15997 16727 16000
rect 16669 15991 16727 15997
rect 12452 15932 13032 15960
rect 13740 15960 13768 15991
rect 13814 15960 13820 15972
rect 13740 15932 13820 15960
rect 13814 15920 13820 15932
rect 13872 15920 13878 15972
rect 14844 15960 14872 15991
rect 16942 15988 16948 16000
rect 17000 15988 17006 16040
rect 17037 16031 17095 16037
rect 17037 15997 17049 16031
rect 17083 15997 17095 16031
rect 19702 16028 19708 16040
rect 17037 15991 17095 15997
rect 17880 16000 19708 16028
rect 14016 15932 14872 15960
rect 11974 15892 11980 15904
rect 11532 15864 11980 15892
rect 11974 15852 11980 15864
rect 12032 15852 12038 15904
rect 13725 15895 13783 15901
rect 13725 15861 13737 15895
rect 13771 15892 13783 15895
rect 14016 15892 14044 15932
rect 15378 15920 15384 15972
rect 15436 15960 15442 15972
rect 16114 15960 16120 15972
rect 15436 15932 16120 15960
rect 15436 15920 15442 15932
rect 16114 15920 16120 15932
rect 16172 15960 16178 15972
rect 17052 15960 17080 15991
rect 17402 15960 17408 15972
rect 16172 15932 17080 15960
rect 17144 15932 17408 15960
rect 16172 15920 16178 15932
rect 13771 15864 14044 15892
rect 13771 15861 13783 15864
rect 13725 15855 13783 15861
rect 14642 15852 14648 15904
rect 14700 15892 14706 15904
rect 15197 15895 15255 15901
rect 15197 15892 15209 15895
rect 14700 15864 15209 15892
rect 14700 15852 14706 15864
rect 15197 15861 15209 15864
rect 15243 15861 15255 15895
rect 15197 15855 15255 15861
rect 16206 15852 16212 15904
rect 16264 15892 16270 15904
rect 17144 15892 17172 15932
rect 17402 15920 17408 15932
rect 17460 15920 17466 15972
rect 17880 15904 17908 16000
rect 19702 15988 19708 16000
rect 19760 16028 19766 16040
rect 19797 16031 19855 16037
rect 19797 16028 19809 16031
rect 19760 16000 19809 16028
rect 19760 15988 19766 16000
rect 19797 15997 19809 16000
rect 19843 15997 19855 16031
rect 19797 15991 19855 15997
rect 20070 15988 20076 16040
rect 20128 15988 20134 16040
rect 20257 16031 20315 16037
rect 20257 15997 20269 16031
rect 20303 16028 20315 16031
rect 20438 16028 20444 16040
rect 20303 16000 20444 16028
rect 20303 15997 20315 16000
rect 20257 15991 20315 15997
rect 20438 15988 20444 16000
rect 20496 15988 20502 16040
rect 21358 15988 21364 16040
rect 21416 15988 21422 16040
rect 21652 16037 21680 16068
rect 22094 16056 22100 16068
rect 22152 16056 22158 16108
rect 22186 16056 22192 16108
rect 22244 16096 22250 16108
rect 22649 16099 22707 16105
rect 22649 16096 22661 16099
rect 22244 16068 22661 16096
rect 22244 16056 22250 16068
rect 22649 16065 22661 16068
rect 22695 16065 22707 16099
rect 22649 16059 22707 16065
rect 21545 16031 21603 16037
rect 21545 15997 21557 16031
rect 21591 15997 21603 16031
rect 21545 15991 21603 15997
rect 21637 16031 21695 16037
rect 21637 15997 21649 16031
rect 21683 15997 21695 16031
rect 21637 15991 21695 15997
rect 21560 15960 21588 15991
rect 21910 15988 21916 16040
rect 21968 15988 21974 16040
rect 22281 16031 22339 16037
rect 22281 15997 22293 16031
rect 22327 15997 22339 16031
rect 22281 15991 22339 15997
rect 22002 15960 22008 15972
rect 19996 15932 22008 15960
rect 16264 15864 17172 15892
rect 17221 15895 17279 15901
rect 16264 15852 16270 15864
rect 17221 15861 17233 15895
rect 17267 15892 17279 15895
rect 17862 15892 17868 15904
rect 17267 15864 17868 15892
rect 17267 15861 17279 15864
rect 17221 15855 17279 15861
rect 17862 15852 17868 15864
rect 17920 15852 17926 15904
rect 19426 15852 19432 15904
rect 19484 15892 19490 15904
rect 19996 15901 20024 15932
rect 22002 15920 22008 15932
rect 22060 15920 22066 15972
rect 22296 15960 22324 15991
rect 22370 15988 22376 16040
rect 22428 16028 22434 16040
rect 22557 16031 22615 16037
rect 22557 16028 22569 16031
rect 22428 16000 22569 16028
rect 22428 15988 22434 16000
rect 22557 15997 22569 16000
rect 22603 15997 22615 16031
rect 22557 15991 22615 15997
rect 22738 15988 22744 16040
rect 22796 15988 22802 16040
rect 23017 16031 23075 16037
rect 23017 15997 23029 16031
rect 23063 16028 23075 16031
rect 23106 16028 23112 16040
rect 23063 16000 23112 16028
rect 23063 15997 23075 16000
rect 23017 15991 23075 15997
rect 23106 15988 23112 16000
rect 23164 15988 23170 16040
rect 23474 15960 23480 15972
rect 22296 15932 23480 15960
rect 23474 15920 23480 15932
rect 23532 15920 23538 15972
rect 19981 15895 20039 15901
rect 19981 15892 19993 15895
rect 19484 15864 19993 15892
rect 19484 15852 19490 15864
rect 19981 15861 19993 15864
rect 20027 15861 20039 15895
rect 19981 15855 20039 15861
rect 20257 15895 20315 15901
rect 20257 15861 20269 15895
rect 20303 15892 20315 15895
rect 20346 15892 20352 15904
rect 20303 15864 20352 15892
rect 20303 15861 20315 15864
rect 20257 15855 20315 15861
rect 20346 15852 20352 15864
rect 20404 15852 20410 15904
rect 21453 15895 21511 15901
rect 21453 15861 21465 15895
rect 21499 15892 21511 15895
rect 21818 15892 21824 15904
rect 21499 15864 21824 15892
rect 21499 15861 21511 15864
rect 21453 15855 21511 15861
rect 21818 15852 21824 15864
rect 21876 15852 21882 15904
rect 552 15802 23368 15824
rect 552 15750 4366 15802
rect 4418 15750 4430 15802
rect 4482 15750 4494 15802
rect 4546 15750 4558 15802
rect 4610 15750 4622 15802
rect 4674 15750 4686 15802
rect 4738 15750 10366 15802
rect 10418 15750 10430 15802
rect 10482 15750 10494 15802
rect 10546 15750 10558 15802
rect 10610 15750 10622 15802
rect 10674 15750 10686 15802
rect 10738 15750 16366 15802
rect 16418 15750 16430 15802
rect 16482 15750 16494 15802
rect 16546 15750 16558 15802
rect 16610 15750 16622 15802
rect 16674 15750 16686 15802
rect 16738 15750 22366 15802
rect 22418 15750 22430 15802
rect 22482 15750 22494 15802
rect 22546 15750 22558 15802
rect 22610 15750 22622 15802
rect 22674 15750 22686 15802
rect 22738 15750 23368 15802
rect 552 15728 23368 15750
rect 2958 15648 2964 15700
rect 3016 15648 3022 15700
rect 3786 15648 3792 15700
rect 3844 15648 3850 15700
rect 5442 15648 5448 15700
rect 5500 15688 5506 15700
rect 6457 15691 6515 15697
rect 6457 15688 6469 15691
rect 5500 15660 6469 15688
rect 5500 15648 5506 15660
rect 6457 15657 6469 15660
rect 6503 15657 6515 15691
rect 6457 15651 6515 15657
rect 6638 15648 6644 15700
rect 6696 15688 6702 15700
rect 6917 15691 6975 15697
rect 6917 15688 6929 15691
rect 6696 15660 6929 15688
rect 6696 15648 6702 15660
rect 6917 15657 6929 15660
rect 6963 15657 6975 15691
rect 7374 15688 7380 15700
rect 6917 15651 6975 15657
rect 7208 15660 7380 15688
rect 934 15580 940 15632
rect 992 15620 998 15632
rect 1210 15620 1216 15632
rect 992 15592 1216 15620
rect 992 15580 998 15592
rect 1210 15580 1216 15592
rect 1268 15580 1274 15632
rect 1429 15623 1487 15629
rect 1429 15589 1441 15623
rect 1475 15620 1487 15623
rect 1765 15623 1823 15629
rect 1765 15620 1777 15623
rect 1475 15592 1777 15620
rect 1475 15589 1487 15592
rect 1429 15583 1487 15589
rect 1765 15589 1777 15592
rect 1811 15589 1823 15623
rect 1765 15583 1823 15589
rect 2409 15623 2467 15629
rect 2409 15589 2421 15623
rect 2455 15620 2467 15623
rect 2774 15620 2780 15632
rect 2455 15592 2780 15620
rect 2455 15589 2467 15592
rect 2409 15583 2467 15589
rect 2746 15580 2780 15592
rect 2832 15580 2838 15632
rect 3234 15580 3240 15632
rect 3292 15620 3298 15632
rect 3881 15623 3939 15629
rect 3881 15620 3893 15623
rect 3292 15592 3893 15620
rect 3292 15580 3298 15592
rect 3881 15589 3893 15592
rect 3927 15589 3939 15623
rect 3881 15583 3939 15589
rect 5534 15580 5540 15632
rect 5592 15620 5598 15632
rect 5629 15623 5687 15629
rect 5629 15620 5641 15623
rect 5592 15592 5641 15620
rect 5592 15580 5598 15592
rect 5629 15589 5641 15592
rect 5675 15589 5687 15623
rect 5629 15583 5687 15589
rect 1670 15512 1676 15564
rect 1728 15512 1734 15564
rect 1857 15555 1915 15561
rect 1857 15521 1869 15555
rect 1903 15552 1915 15555
rect 1946 15552 1952 15564
rect 1903 15524 1952 15552
rect 1903 15521 1915 15524
rect 1857 15515 1915 15521
rect 1946 15512 1952 15524
rect 2004 15512 2010 15564
rect 2314 15512 2320 15564
rect 2372 15552 2378 15564
rect 2593 15555 2651 15561
rect 2593 15552 2605 15555
rect 2372 15524 2605 15552
rect 2372 15512 2378 15524
rect 2593 15521 2605 15524
rect 2639 15521 2651 15555
rect 2746 15552 2774 15580
rect 2869 15555 2927 15561
rect 2869 15552 2881 15555
rect 2746 15524 2881 15552
rect 2593 15515 2651 15521
rect 2869 15521 2881 15524
rect 2915 15521 2927 15555
rect 3602 15552 3608 15564
rect 2869 15515 2927 15521
rect 3160 15524 3608 15552
rect 2777 15487 2835 15493
rect 2777 15453 2789 15487
rect 2823 15484 2835 15487
rect 3160 15484 3188 15524
rect 3602 15512 3608 15524
rect 3660 15512 3666 15564
rect 5997 15555 6055 15561
rect 5997 15521 6009 15555
rect 6043 15552 6055 15555
rect 6546 15552 6552 15564
rect 6043 15524 6552 15552
rect 6043 15521 6055 15524
rect 5997 15515 6055 15521
rect 6546 15512 6552 15524
rect 6604 15512 6610 15564
rect 7098 15512 7104 15564
rect 7156 15512 7162 15564
rect 7208 15561 7236 15660
rect 7374 15648 7380 15660
rect 7432 15648 7438 15700
rect 9490 15648 9496 15700
rect 9548 15688 9554 15700
rect 11149 15691 11207 15697
rect 11149 15688 11161 15691
rect 9548 15660 10640 15688
rect 9548 15648 9554 15660
rect 8294 15580 8300 15632
rect 8352 15580 8358 15632
rect 8389 15623 8447 15629
rect 8389 15589 8401 15623
rect 8435 15620 8447 15623
rect 8478 15620 8484 15632
rect 8435 15592 8484 15620
rect 8435 15589 8447 15592
rect 8389 15583 8447 15589
rect 8478 15580 8484 15592
rect 8536 15580 8542 15632
rect 8605 15623 8663 15629
rect 8605 15589 8617 15623
rect 8651 15620 8663 15623
rect 9582 15620 9588 15632
rect 8651 15592 9588 15620
rect 8651 15589 8663 15592
rect 8605 15583 8663 15589
rect 9582 15580 9588 15592
rect 9640 15580 9646 15632
rect 9950 15580 9956 15632
rect 10008 15620 10014 15632
rect 10505 15623 10563 15629
rect 10505 15620 10517 15623
rect 10008 15592 10517 15620
rect 10008 15580 10014 15592
rect 10505 15589 10517 15592
rect 10551 15589 10563 15623
rect 10505 15583 10563 15589
rect 7193 15555 7251 15561
rect 7193 15521 7205 15555
rect 7239 15521 7251 15555
rect 7193 15515 7251 15521
rect 7374 15512 7380 15564
rect 7432 15512 7438 15564
rect 7653 15555 7711 15561
rect 7653 15521 7665 15555
rect 7699 15552 7711 15555
rect 7926 15552 7932 15564
rect 7699 15524 7932 15552
rect 7699 15521 7711 15524
rect 7653 15515 7711 15521
rect 7926 15512 7932 15524
rect 7984 15512 7990 15564
rect 8312 15545 8340 15580
rect 8297 15539 8355 15545
rect 8297 15505 8309 15539
rect 8343 15505 8355 15539
rect 9030 15512 9036 15564
rect 9088 15552 9094 15564
rect 9088 15524 9444 15552
rect 9088 15512 9094 15524
rect 8297 15499 8355 15505
rect 9416 15496 9444 15524
rect 9674 15512 9680 15564
rect 9732 15512 9738 15564
rect 9766 15512 9772 15564
rect 9824 15552 9830 15564
rect 9861 15555 9919 15561
rect 9861 15552 9873 15555
rect 9824 15524 9873 15552
rect 9824 15512 9830 15524
rect 9861 15521 9873 15524
rect 9907 15521 9919 15555
rect 9861 15515 9919 15521
rect 10042 15512 10048 15564
rect 10100 15552 10106 15564
rect 10229 15555 10287 15561
rect 10229 15552 10241 15555
rect 10100 15524 10241 15552
rect 10100 15512 10106 15524
rect 10229 15521 10241 15524
rect 10275 15552 10287 15555
rect 10318 15552 10324 15564
rect 10275 15524 10324 15552
rect 10275 15521 10287 15524
rect 10229 15515 10287 15521
rect 10318 15512 10324 15524
rect 10376 15512 10382 15564
rect 2823 15456 3188 15484
rect 2823 15453 2835 15456
rect 2777 15447 2835 15453
rect 3326 15444 3332 15496
rect 3384 15444 3390 15496
rect 5442 15484 5448 15496
rect 3620 15456 5448 15484
rect 1854 15416 1860 15428
rect 1412 15388 1860 15416
rect 1412 15357 1440 15388
rect 1854 15376 1860 15388
rect 1912 15376 1918 15428
rect 3142 15416 3148 15428
rect 2746 15388 3148 15416
rect 1397 15351 1455 15357
rect 1397 15317 1409 15351
rect 1443 15317 1455 15351
rect 1397 15311 1455 15317
rect 1581 15351 1639 15357
rect 1581 15317 1593 15351
rect 1627 15348 1639 15351
rect 2746 15348 2774 15388
rect 3142 15376 3148 15388
rect 3200 15376 3206 15428
rect 3620 15425 3648 15456
rect 5442 15444 5448 15456
rect 5500 15444 5506 15496
rect 6270 15444 6276 15496
rect 6328 15444 6334 15496
rect 6365 15487 6423 15493
rect 6365 15453 6377 15487
rect 6411 15484 6423 15487
rect 7285 15487 7343 15493
rect 7285 15484 7297 15487
rect 6411 15456 7297 15484
rect 6411 15453 6423 15456
rect 6365 15447 6423 15453
rect 7285 15453 7297 15456
rect 7331 15453 7343 15487
rect 7285 15447 7343 15453
rect 9214 15444 9220 15496
rect 9272 15444 9278 15496
rect 9306 15444 9312 15496
rect 9364 15444 9370 15496
rect 9398 15444 9404 15496
rect 9456 15444 9462 15496
rect 9493 15487 9551 15493
rect 9493 15453 9505 15487
rect 9539 15484 9551 15487
rect 10134 15484 10140 15496
rect 9539 15456 10140 15484
rect 9539 15453 9551 15456
rect 9493 15447 9551 15453
rect 10134 15444 10140 15456
rect 10192 15484 10198 15496
rect 10410 15484 10416 15496
rect 10192 15456 10416 15484
rect 10192 15444 10198 15456
rect 10410 15444 10416 15456
rect 10468 15444 10474 15496
rect 3605 15419 3663 15425
rect 3605 15385 3617 15419
rect 3651 15385 3663 15419
rect 5813 15419 5871 15425
rect 5813 15416 5825 15419
rect 3605 15379 3663 15385
rect 4816 15388 5825 15416
rect 1627 15320 2774 15348
rect 1627 15317 1639 15320
rect 1581 15311 1639 15317
rect 3050 15308 3056 15360
rect 3108 15348 3114 15360
rect 4816 15348 4844 15388
rect 5813 15385 5825 15388
rect 5859 15416 5871 15419
rect 6454 15416 6460 15428
rect 5859 15388 6460 15416
rect 5859 15385 5871 15388
rect 5813 15379 5871 15385
rect 6454 15376 6460 15388
rect 6512 15376 6518 15428
rect 6914 15376 6920 15428
rect 6972 15416 6978 15428
rect 7469 15419 7527 15425
rect 7469 15416 7481 15419
rect 6972 15388 7481 15416
rect 6972 15376 6978 15388
rect 7469 15385 7481 15388
rect 7515 15416 7527 15419
rect 8202 15416 8208 15428
rect 7515 15388 8208 15416
rect 7515 15385 7527 15388
rect 7469 15379 7527 15385
rect 8202 15376 8208 15388
rect 8260 15376 8266 15428
rect 9582 15376 9588 15428
rect 9640 15416 9646 15428
rect 9861 15419 9919 15425
rect 9861 15416 9873 15419
rect 9640 15388 9873 15416
rect 9640 15376 9646 15388
rect 9861 15385 9873 15388
rect 9907 15385 9919 15419
rect 9861 15379 9919 15385
rect 10226 15376 10232 15428
rect 10284 15416 10290 15428
rect 10321 15419 10379 15425
rect 10321 15416 10333 15419
rect 10284 15388 10333 15416
rect 10284 15376 10290 15388
rect 10321 15385 10333 15388
rect 10367 15385 10379 15419
rect 10321 15379 10379 15385
rect 3108 15320 4844 15348
rect 3108 15308 3114 15320
rect 6362 15308 6368 15360
rect 6420 15348 6426 15360
rect 6825 15351 6883 15357
rect 6825 15348 6837 15351
rect 6420 15320 6837 15348
rect 6420 15308 6426 15320
rect 6825 15317 6837 15320
rect 6871 15317 6883 15351
rect 6825 15311 6883 15317
rect 8110 15308 8116 15360
rect 8168 15308 8174 15360
rect 8294 15308 8300 15360
rect 8352 15348 8358 15360
rect 8573 15351 8631 15357
rect 8573 15348 8585 15351
rect 8352 15320 8585 15348
rect 8352 15308 8358 15320
rect 8573 15317 8585 15320
rect 8619 15317 8631 15351
rect 8573 15311 8631 15317
rect 8757 15351 8815 15357
rect 8757 15317 8769 15351
rect 8803 15348 8815 15351
rect 8846 15348 8852 15360
rect 8803 15320 8852 15348
rect 8803 15317 8815 15320
rect 8757 15311 8815 15317
rect 8846 15308 8852 15320
rect 8904 15308 8910 15360
rect 9033 15351 9091 15357
rect 9033 15317 9045 15351
rect 9079 15348 9091 15351
rect 9398 15348 9404 15360
rect 9079 15320 9404 15348
rect 9079 15317 9091 15320
rect 9033 15311 9091 15317
rect 9398 15308 9404 15320
rect 9456 15308 9462 15360
rect 10520 15348 10548 15583
rect 10612 15552 10640 15660
rect 10704 15660 11161 15688
rect 10704 15629 10732 15660
rect 11149 15657 11161 15660
rect 11195 15688 11207 15691
rect 11790 15688 11796 15700
rect 11195 15660 11796 15688
rect 11195 15657 11207 15660
rect 11149 15651 11207 15657
rect 11790 15648 11796 15660
rect 11848 15688 11854 15700
rect 11848 15660 12756 15688
rect 11848 15648 11854 15660
rect 10689 15623 10747 15629
rect 10689 15589 10701 15623
rect 10735 15589 10747 15623
rect 10689 15583 10747 15589
rect 10796 15592 11100 15620
rect 10796 15552 10824 15592
rect 10612 15524 10824 15552
rect 10962 15512 10968 15564
rect 11020 15512 11026 15564
rect 11072 15552 11100 15592
rect 12158 15580 12164 15632
rect 12216 15620 12222 15632
rect 12253 15623 12311 15629
rect 12253 15620 12265 15623
rect 12216 15592 12265 15620
rect 12216 15580 12222 15592
rect 12253 15589 12265 15592
rect 12299 15589 12311 15623
rect 12253 15583 12311 15589
rect 12360 15592 12664 15620
rect 12360 15552 12388 15592
rect 11072 15524 12388 15552
rect 12434 15512 12440 15564
rect 12492 15512 12498 15564
rect 10686 15444 10692 15496
rect 10744 15484 10750 15496
rect 11330 15484 11336 15496
rect 10744 15456 11336 15484
rect 10744 15444 10750 15456
rect 11330 15444 11336 15456
rect 11388 15484 11394 15496
rect 11790 15484 11796 15496
rect 11388 15456 11796 15484
rect 11388 15444 11394 15456
rect 11790 15444 11796 15456
rect 11848 15444 11854 15496
rect 12636 15484 12664 15592
rect 12728 15561 12756 15660
rect 13538 15648 13544 15700
rect 13596 15688 13602 15700
rect 13725 15691 13783 15697
rect 13725 15688 13737 15691
rect 13596 15660 13737 15688
rect 13596 15648 13602 15660
rect 13725 15657 13737 15660
rect 13771 15657 13783 15691
rect 13725 15651 13783 15657
rect 13814 15648 13820 15700
rect 13872 15688 13878 15700
rect 13909 15691 13967 15697
rect 13909 15688 13921 15691
rect 13872 15660 13921 15688
rect 13872 15648 13878 15660
rect 13909 15657 13921 15660
rect 13955 15657 13967 15691
rect 13909 15651 13967 15657
rect 15194 15648 15200 15700
rect 15252 15688 15258 15700
rect 15381 15691 15439 15697
rect 15381 15688 15393 15691
rect 15252 15660 15393 15688
rect 15252 15648 15258 15660
rect 15381 15657 15393 15660
rect 15427 15688 15439 15691
rect 17586 15688 17592 15700
rect 15427 15660 17592 15688
rect 15427 15657 15439 15660
rect 15381 15651 15439 15657
rect 17586 15648 17592 15660
rect 17644 15648 17650 15700
rect 18046 15648 18052 15700
rect 18104 15688 18110 15700
rect 19521 15691 19579 15697
rect 19521 15688 19533 15691
rect 18104 15660 19533 15688
rect 18104 15648 18110 15660
rect 19521 15657 19533 15660
rect 19567 15688 19579 15691
rect 22462 15688 22468 15700
rect 19567 15660 20024 15688
rect 19567 15657 19579 15660
rect 19521 15651 19579 15657
rect 16206 15620 16212 15632
rect 12912 15592 16212 15620
rect 12912 15561 12940 15592
rect 13556 15561 13584 15592
rect 16206 15580 16212 15592
rect 16264 15580 16270 15632
rect 17402 15580 17408 15632
rect 17460 15620 17466 15632
rect 17460 15592 18920 15620
rect 17460 15580 17466 15592
rect 12713 15555 12771 15561
rect 12713 15521 12725 15555
rect 12759 15521 12771 15555
rect 12713 15515 12771 15521
rect 12897 15555 12955 15561
rect 12897 15521 12909 15555
rect 12943 15521 12955 15555
rect 12897 15515 12955 15521
rect 13357 15555 13415 15561
rect 13357 15521 13369 15555
rect 13403 15521 13415 15555
rect 13357 15515 13415 15521
rect 13541 15555 13599 15561
rect 13541 15521 13553 15555
rect 13587 15521 13599 15555
rect 13541 15515 13599 15521
rect 13372 15484 13400 15515
rect 13814 15512 13820 15564
rect 13872 15512 13878 15564
rect 14001 15555 14059 15561
rect 14001 15521 14013 15555
rect 14047 15521 14059 15555
rect 14001 15515 14059 15521
rect 14645 15555 14703 15561
rect 14645 15521 14657 15555
rect 14691 15552 14703 15555
rect 14826 15552 14832 15564
rect 14691 15524 14832 15552
rect 14691 15521 14703 15524
rect 14645 15515 14703 15521
rect 13906 15484 13912 15496
rect 12636 15456 13912 15484
rect 13906 15444 13912 15456
rect 13964 15444 13970 15496
rect 14016 15484 14044 15515
rect 14826 15512 14832 15524
rect 14884 15512 14890 15564
rect 15010 15512 15016 15564
rect 15068 15552 15074 15564
rect 15105 15555 15163 15561
rect 15105 15552 15117 15555
rect 15068 15524 15117 15552
rect 15068 15512 15074 15524
rect 15105 15521 15117 15524
rect 15151 15521 15163 15555
rect 15105 15515 15163 15521
rect 15565 15555 15623 15561
rect 15565 15521 15577 15555
rect 15611 15521 15623 15555
rect 15565 15515 15623 15521
rect 15580 15484 15608 15515
rect 15654 15512 15660 15564
rect 15712 15512 15718 15564
rect 15746 15512 15752 15564
rect 15804 15552 15810 15564
rect 16577 15555 16635 15561
rect 16577 15552 16589 15555
rect 15804 15524 16589 15552
rect 15804 15512 15810 15524
rect 16577 15521 16589 15524
rect 16623 15552 16635 15555
rect 16623 15524 17816 15552
rect 16623 15521 16635 15524
rect 16577 15515 16635 15521
rect 14016 15456 15884 15484
rect 15120 15428 15148 15456
rect 10870 15376 10876 15428
rect 10928 15416 10934 15428
rect 12250 15416 12256 15428
rect 10928 15388 12256 15416
rect 10928 15376 10934 15388
rect 12250 15376 12256 15388
rect 12308 15376 12314 15428
rect 14090 15416 14096 15428
rect 12544 15388 14096 15416
rect 12544 15348 12572 15388
rect 14090 15376 14096 15388
rect 14148 15416 14154 15428
rect 14461 15419 14519 15425
rect 14461 15416 14473 15419
rect 14148 15388 14473 15416
rect 14148 15376 14154 15388
rect 14461 15385 14473 15388
rect 14507 15416 14519 15419
rect 14918 15416 14924 15428
rect 14507 15388 14924 15416
rect 14507 15385 14519 15388
rect 14461 15379 14519 15385
rect 14918 15376 14924 15388
rect 14976 15376 14982 15428
rect 15102 15376 15108 15428
rect 15160 15376 15166 15428
rect 15289 15419 15347 15425
rect 15289 15385 15301 15419
rect 15335 15416 15347 15419
rect 15470 15416 15476 15428
rect 15335 15388 15476 15416
rect 15335 15385 15347 15388
rect 15289 15379 15347 15385
rect 15470 15376 15476 15388
rect 15528 15376 15534 15428
rect 15856 15425 15884 15456
rect 16114 15444 16120 15496
rect 16172 15484 16178 15496
rect 16669 15487 16727 15493
rect 16669 15484 16681 15487
rect 16172 15456 16681 15484
rect 16172 15444 16178 15456
rect 16669 15453 16681 15456
rect 16715 15453 16727 15487
rect 16669 15447 16727 15453
rect 16945 15487 17003 15493
rect 16945 15453 16957 15487
rect 16991 15484 17003 15487
rect 17126 15484 17132 15496
rect 16991 15456 17132 15484
rect 16991 15453 17003 15456
rect 16945 15447 17003 15453
rect 17126 15444 17132 15456
rect 17184 15484 17190 15496
rect 17221 15487 17279 15493
rect 17221 15484 17233 15487
rect 17184 15456 17233 15484
rect 17184 15444 17190 15456
rect 17221 15453 17233 15456
rect 17267 15453 17279 15487
rect 17221 15447 17279 15453
rect 17313 15487 17371 15493
rect 17313 15453 17325 15487
rect 17359 15453 17371 15487
rect 17313 15447 17371 15453
rect 15841 15419 15899 15425
rect 15841 15385 15853 15419
rect 15887 15385 15899 15419
rect 15841 15379 15899 15385
rect 10520 15320 12572 15348
rect 12621 15351 12679 15357
rect 12621 15317 12633 15351
rect 12667 15348 12679 15351
rect 12710 15348 12716 15360
rect 12667 15320 12716 15348
rect 12667 15317 12679 15320
rect 12621 15311 12679 15317
rect 12710 15308 12716 15320
rect 12768 15308 12774 15360
rect 12805 15351 12863 15357
rect 12805 15317 12817 15351
rect 12851 15348 12863 15351
rect 12986 15348 12992 15360
rect 12851 15320 12992 15348
rect 12851 15317 12863 15320
rect 12805 15311 12863 15317
rect 12986 15308 12992 15320
rect 13044 15308 13050 15360
rect 14829 15351 14887 15357
rect 14829 15317 14841 15351
rect 14875 15348 14887 15351
rect 15010 15348 15016 15360
rect 14875 15320 15016 15348
rect 14875 15317 14887 15320
rect 14829 15311 14887 15317
rect 15010 15308 15016 15320
rect 15068 15308 15074 15360
rect 15488 15348 15516 15376
rect 16482 15348 16488 15360
rect 15488 15320 16488 15348
rect 16482 15308 16488 15320
rect 16540 15308 16546 15360
rect 16758 15308 16764 15360
rect 16816 15348 16822 15360
rect 17037 15351 17095 15357
rect 17037 15348 17049 15351
rect 16816 15320 17049 15348
rect 16816 15308 16822 15320
rect 17037 15317 17049 15320
rect 17083 15317 17095 15351
rect 17328 15348 17356 15447
rect 17402 15444 17408 15496
rect 17460 15444 17466 15496
rect 17497 15487 17555 15493
rect 17497 15453 17509 15487
rect 17543 15484 17555 15487
rect 17681 15487 17739 15493
rect 17681 15484 17693 15487
rect 17543 15456 17693 15484
rect 17543 15453 17555 15456
rect 17497 15447 17555 15453
rect 17681 15453 17693 15456
rect 17727 15453 17739 15487
rect 17788 15484 17816 15524
rect 17862 15512 17868 15564
rect 17920 15552 17926 15564
rect 18892 15561 18920 15592
rect 18325 15555 18383 15561
rect 18325 15552 18337 15555
rect 17920 15524 18337 15552
rect 17920 15512 17926 15524
rect 18325 15521 18337 15524
rect 18371 15521 18383 15555
rect 18325 15515 18383 15521
rect 18601 15555 18659 15561
rect 18601 15521 18613 15555
rect 18647 15521 18659 15555
rect 18601 15515 18659 15521
rect 18785 15555 18843 15561
rect 18785 15521 18797 15555
rect 18831 15521 18843 15555
rect 18785 15515 18843 15521
rect 18877 15555 18935 15561
rect 18877 15521 18889 15555
rect 18923 15521 18935 15555
rect 18877 15515 18935 15521
rect 19061 15555 19119 15561
rect 19061 15521 19073 15555
rect 19107 15552 19119 15555
rect 19426 15552 19432 15564
rect 19107 15524 19432 15552
rect 19107 15521 19119 15524
rect 19061 15515 19119 15521
rect 18049 15487 18107 15493
rect 18049 15484 18061 15487
rect 17788 15456 18061 15484
rect 17681 15447 17739 15453
rect 18049 15453 18061 15456
rect 18095 15453 18107 15487
rect 18049 15447 18107 15453
rect 18141 15487 18199 15493
rect 18141 15453 18153 15487
rect 18187 15484 18199 15487
rect 18230 15484 18236 15496
rect 18187 15456 18236 15484
rect 18187 15453 18199 15456
rect 18141 15447 18199 15453
rect 18230 15444 18236 15456
rect 18288 15444 18294 15496
rect 18509 15419 18567 15425
rect 18509 15385 18521 15419
rect 18555 15416 18567 15419
rect 18616 15416 18644 15515
rect 18690 15444 18696 15496
rect 18748 15444 18754 15496
rect 18800 15484 18828 15515
rect 19426 15512 19432 15524
rect 19484 15512 19490 15564
rect 19702 15512 19708 15564
rect 19760 15552 19766 15564
rect 19889 15555 19947 15561
rect 19889 15552 19901 15555
rect 19760 15524 19901 15552
rect 19760 15512 19766 15524
rect 19889 15521 19901 15524
rect 19935 15521 19947 15555
rect 19996 15552 20024 15660
rect 22066 15660 22468 15688
rect 20162 15580 20168 15632
rect 20220 15620 20226 15632
rect 20625 15623 20683 15629
rect 20625 15620 20637 15623
rect 20220 15592 20637 15620
rect 20220 15580 20226 15592
rect 20625 15589 20637 15592
rect 20671 15589 20683 15623
rect 20625 15583 20683 15589
rect 20993 15623 21051 15629
rect 20993 15589 21005 15623
rect 21039 15620 21051 15623
rect 22066 15620 22094 15660
rect 22462 15648 22468 15660
rect 22520 15648 22526 15700
rect 22830 15648 22836 15700
rect 22888 15648 22894 15700
rect 21039 15592 22094 15620
rect 22373 15623 22431 15629
rect 21039 15589 21051 15592
rect 20993 15583 21051 15589
rect 20349 15555 20407 15561
rect 20349 15552 20361 15555
rect 19996 15524 20361 15552
rect 19889 15515 19947 15521
rect 20349 15521 20361 15524
rect 20395 15521 20407 15555
rect 20349 15515 20407 15521
rect 20806 15512 20812 15564
rect 20864 15552 20870 15564
rect 20901 15555 20959 15561
rect 20901 15552 20913 15555
rect 20864 15524 20913 15552
rect 20864 15512 20870 15524
rect 20901 15521 20913 15524
rect 20947 15521 20959 15555
rect 20901 15515 20959 15521
rect 21082 15512 21088 15564
rect 21140 15512 21146 15564
rect 21637 15555 21695 15561
rect 21637 15521 21649 15555
rect 21683 15521 21695 15555
rect 21637 15515 21695 15521
rect 18969 15487 19027 15493
rect 18969 15484 18981 15487
rect 18800 15456 18981 15484
rect 18969 15453 18981 15456
rect 19015 15453 19027 15487
rect 18969 15447 19027 15453
rect 19981 15487 20039 15493
rect 19981 15453 19993 15487
rect 20027 15484 20039 15487
rect 20027 15456 20392 15484
rect 20027 15453 20039 15456
rect 19981 15447 20039 15453
rect 19150 15416 19156 15428
rect 18555 15388 19156 15416
rect 18555 15385 18567 15388
rect 18509 15379 18567 15385
rect 19150 15376 19156 15388
rect 19208 15376 19214 15428
rect 20364 15360 20392 15456
rect 20438 15444 20444 15496
rect 20496 15484 20502 15496
rect 20625 15487 20683 15493
rect 20625 15484 20637 15487
rect 20496 15456 20637 15484
rect 20496 15444 20502 15456
rect 20625 15453 20637 15456
rect 20671 15453 20683 15487
rect 20625 15447 20683 15453
rect 20530 15376 20536 15428
rect 20588 15416 20594 15428
rect 21082 15416 21088 15428
rect 20588 15388 21088 15416
rect 20588 15376 20594 15388
rect 21082 15376 21088 15388
rect 21140 15376 21146 15428
rect 21652 15416 21680 15515
rect 21818 15512 21824 15564
rect 21876 15512 21882 15564
rect 21928 15561 21956 15592
rect 22373 15589 22385 15623
rect 22419 15620 22431 15623
rect 22419 15592 22784 15620
rect 22419 15589 22431 15592
rect 22373 15583 22431 15589
rect 21913 15555 21971 15561
rect 21913 15521 21925 15555
rect 21959 15521 21971 15555
rect 21913 15515 21971 15521
rect 22002 15512 22008 15564
rect 22060 15512 22066 15564
rect 22094 15512 22100 15564
rect 22152 15552 22158 15564
rect 22189 15555 22247 15561
rect 22189 15552 22201 15555
rect 22152 15524 22201 15552
rect 22152 15512 22158 15524
rect 22189 15521 22201 15524
rect 22235 15521 22247 15555
rect 22189 15515 22247 15521
rect 22278 15512 22284 15564
rect 22336 15512 22342 15564
rect 22756 15561 22784 15592
rect 22557 15555 22615 15561
rect 22557 15521 22569 15555
rect 22603 15521 22615 15555
rect 22557 15515 22615 15521
rect 22741 15555 22799 15561
rect 22741 15521 22753 15555
rect 22787 15521 22799 15555
rect 22741 15515 22799 15521
rect 21836 15484 21864 15512
rect 22572 15484 22600 15515
rect 23014 15512 23020 15564
rect 23072 15512 23078 15564
rect 21836 15456 22600 15484
rect 22097 15419 22155 15425
rect 22097 15416 22109 15419
rect 21652 15388 22109 15416
rect 22097 15385 22109 15388
rect 22143 15416 22155 15419
rect 22278 15416 22284 15428
rect 22143 15388 22284 15416
rect 22143 15385 22155 15388
rect 22097 15379 22155 15385
rect 22278 15376 22284 15388
rect 22336 15376 22342 15428
rect 19242 15348 19248 15360
rect 17328 15320 19248 15348
rect 17037 15311 17095 15317
rect 19242 15308 19248 15320
rect 19300 15308 19306 15360
rect 20254 15308 20260 15360
rect 20312 15308 20318 15360
rect 20346 15308 20352 15360
rect 20404 15348 20410 15360
rect 20441 15351 20499 15357
rect 20441 15348 20453 15351
rect 20404 15320 20453 15348
rect 20404 15308 20410 15320
rect 20441 15317 20453 15320
rect 20487 15317 20499 15351
rect 20441 15311 20499 15317
rect 20714 15308 20720 15360
rect 20772 15348 20778 15360
rect 21453 15351 21511 15357
rect 21453 15348 21465 15351
rect 20772 15320 21465 15348
rect 20772 15308 20778 15320
rect 21453 15317 21465 15320
rect 21499 15317 21511 15351
rect 21453 15311 21511 15317
rect 22554 15308 22560 15360
rect 22612 15308 22618 15360
rect 552 15258 23368 15280
rect 552 15206 1366 15258
rect 1418 15206 1430 15258
rect 1482 15206 1494 15258
rect 1546 15206 1558 15258
rect 1610 15206 1622 15258
rect 1674 15206 1686 15258
rect 1738 15206 7366 15258
rect 7418 15206 7430 15258
rect 7482 15206 7494 15258
rect 7546 15206 7558 15258
rect 7610 15206 7622 15258
rect 7674 15206 7686 15258
rect 7738 15206 13366 15258
rect 13418 15206 13430 15258
rect 13482 15206 13494 15258
rect 13546 15206 13558 15258
rect 13610 15206 13622 15258
rect 13674 15206 13686 15258
rect 13738 15206 19366 15258
rect 19418 15206 19430 15258
rect 19482 15206 19494 15258
rect 19546 15206 19558 15258
rect 19610 15206 19622 15258
rect 19674 15206 19686 15258
rect 19738 15206 23368 15258
rect 552 15184 23368 15206
rect 2498 15104 2504 15156
rect 2556 15144 2562 15156
rect 4433 15147 4491 15153
rect 2556 15116 3648 15144
rect 2556 15104 2562 15116
rect 3234 15076 3240 15088
rect 2332 15048 3240 15076
rect 1210 14900 1216 14952
rect 1268 14940 1274 14952
rect 2332 14949 2360 15048
rect 3234 15036 3240 15048
rect 3292 15036 3298 15088
rect 3620 15076 3648 15116
rect 4433 15113 4445 15147
rect 4479 15144 4491 15147
rect 4706 15144 4712 15156
rect 4479 15116 4712 15144
rect 4479 15113 4491 15116
rect 4433 15107 4491 15113
rect 4706 15104 4712 15116
rect 4764 15104 4770 15156
rect 6365 15147 6423 15153
rect 6365 15113 6377 15147
rect 6411 15144 6423 15147
rect 6546 15144 6552 15156
rect 6411 15116 6552 15144
rect 6411 15113 6423 15116
rect 6365 15107 6423 15113
rect 6546 15104 6552 15116
rect 6604 15104 6610 15156
rect 6825 15147 6883 15153
rect 6825 15113 6837 15147
rect 6871 15144 6883 15147
rect 7190 15144 7196 15156
rect 6871 15116 7196 15144
rect 6871 15113 6883 15116
rect 6825 15107 6883 15113
rect 7190 15104 7196 15116
rect 7248 15104 7254 15156
rect 8478 15144 8484 15156
rect 8404 15116 8484 15144
rect 3620 15048 4476 15076
rect 2498 14968 2504 15020
rect 2556 14968 2562 15020
rect 2866 14968 2872 15020
rect 2924 15008 2930 15020
rect 2961 15011 3019 15017
rect 2961 15008 2973 15011
rect 2924 14980 2973 15008
rect 2924 14968 2930 14980
rect 2961 14977 2973 14980
rect 3007 14977 3019 15011
rect 4154 15008 4160 15020
rect 2961 14971 3019 14977
rect 3804 14980 4160 15008
rect 2317 14943 2375 14949
rect 2317 14940 2329 14943
rect 1268 14912 2329 14940
rect 1268 14900 1274 14912
rect 2317 14909 2329 14912
rect 2363 14909 2375 14943
rect 2317 14903 2375 14909
rect 2590 14900 2596 14952
rect 2648 14900 2654 14952
rect 3804 14949 3832 14980
rect 4154 14968 4160 14980
rect 4212 14968 4218 15020
rect 3329 14943 3387 14949
rect 3329 14909 3341 14943
rect 3375 14940 3387 14943
rect 3789 14943 3847 14949
rect 3789 14940 3801 14943
rect 3375 14912 3801 14940
rect 3375 14909 3387 14912
rect 3329 14903 3387 14909
rect 3789 14909 3801 14912
rect 3835 14909 3847 14943
rect 3789 14903 3847 14909
rect 3973 14943 4031 14949
rect 3973 14909 3985 14943
rect 4019 14909 4031 14943
rect 3973 14903 4031 14909
rect 2072 14875 2130 14881
rect 2072 14841 2084 14875
rect 2118 14872 2130 14875
rect 3418 14872 3424 14884
rect 2118 14844 3424 14872
rect 2118 14841 2130 14844
rect 2072 14835 2130 14841
rect 3418 14832 3424 14844
rect 3476 14832 3482 14884
rect 3878 14872 3884 14884
rect 3528 14844 3884 14872
rect 937 14807 995 14813
rect 937 14773 949 14807
rect 983 14804 995 14807
rect 1578 14804 1584 14816
rect 983 14776 1584 14804
rect 983 14773 995 14776
rect 937 14767 995 14773
rect 1578 14764 1584 14776
rect 1636 14804 1642 14816
rect 1946 14804 1952 14816
rect 1636 14776 1952 14804
rect 1636 14764 1642 14776
rect 1946 14764 1952 14776
rect 2004 14764 2010 14816
rect 3528 14813 3556 14844
rect 3878 14832 3884 14844
rect 3936 14832 3942 14884
rect 3988 14872 4016 14903
rect 4062 14900 4068 14952
rect 4120 14940 4126 14952
rect 4249 14943 4307 14949
rect 4249 14940 4261 14943
rect 4120 14912 4261 14940
rect 4120 14900 4126 14912
rect 4249 14909 4261 14912
rect 4295 14940 4307 14943
rect 4338 14940 4344 14952
rect 4295 14912 4344 14940
rect 4295 14909 4307 14912
rect 4249 14903 4307 14909
rect 4338 14900 4344 14912
rect 4396 14900 4402 14952
rect 4448 14940 4476 15048
rect 6454 15036 6460 15088
rect 6512 15036 6518 15088
rect 4890 14968 4896 15020
rect 4948 14968 4954 15020
rect 6104 14980 6684 15008
rect 4798 14940 4804 14952
rect 4448 14912 4804 14940
rect 4798 14900 4804 14912
rect 4856 14940 4862 14952
rect 4985 14943 5043 14949
rect 4985 14940 4997 14943
rect 4856 14912 4997 14940
rect 4856 14900 4862 14912
rect 4985 14909 4997 14912
rect 5031 14909 5043 14943
rect 4985 14903 5043 14909
rect 5077 14943 5135 14949
rect 5077 14909 5089 14943
rect 5123 14940 5135 14943
rect 5534 14940 5540 14952
rect 5123 14912 5540 14940
rect 5123 14909 5135 14912
rect 5077 14903 5135 14909
rect 5534 14900 5540 14912
rect 5592 14940 5598 14952
rect 5837 14943 5895 14949
rect 5592 14912 5764 14940
rect 5592 14900 5598 14912
rect 4430 14872 4436 14884
rect 3988 14844 4436 14872
rect 4430 14832 4436 14844
rect 4488 14832 4494 14884
rect 4706 14832 4712 14884
rect 4764 14832 4770 14884
rect 4890 14832 4896 14884
rect 4948 14872 4954 14884
rect 5166 14872 5172 14884
rect 4948 14844 5172 14872
rect 4948 14832 4954 14844
rect 5166 14832 5172 14844
rect 5224 14832 5230 14884
rect 5445 14875 5503 14881
rect 5445 14841 5457 14875
rect 5491 14841 5503 14875
rect 5736 14872 5764 14912
rect 5837 14909 5849 14943
rect 5883 14940 5895 14943
rect 6104 14940 6132 14980
rect 5883 14912 6132 14940
rect 5883 14909 5895 14912
rect 5837 14903 5895 14909
rect 6178 14900 6184 14952
rect 6236 14900 6242 14952
rect 6656 14949 6684 14980
rect 6641 14943 6699 14949
rect 6641 14909 6653 14943
rect 6687 14909 6699 14943
rect 6641 14903 6699 14909
rect 6270 14872 6276 14884
rect 5736 14844 6276 14872
rect 5445 14835 5503 14841
rect 3513 14807 3571 14813
rect 3513 14773 3525 14807
rect 3559 14773 3571 14807
rect 3513 14767 3571 14773
rect 3694 14764 3700 14816
rect 3752 14764 3758 14816
rect 3786 14764 3792 14816
rect 3844 14804 3850 14816
rect 4065 14807 4123 14813
rect 4065 14804 4077 14807
rect 3844 14776 4077 14804
rect 3844 14764 3850 14776
rect 4065 14773 4077 14776
rect 4111 14804 4123 14807
rect 5460 14804 5488 14835
rect 6270 14832 6276 14844
rect 6328 14832 6334 14884
rect 6656 14872 6684 14903
rect 6914 14900 6920 14952
rect 6972 14900 6978 14952
rect 7009 14943 7067 14949
rect 7009 14909 7021 14943
rect 7055 14909 7067 14943
rect 7009 14903 7067 14909
rect 7285 14943 7343 14949
rect 7285 14909 7297 14943
rect 7331 14940 7343 14943
rect 7834 14940 7840 14952
rect 7331 14912 7840 14940
rect 7331 14909 7343 14912
rect 7285 14903 7343 14909
rect 7024 14872 7052 14903
rect 7834 14900 7840 14912
rect 7892 14900 7898 14952
rect 8205 14943 8263 14949
rect 8205 14909 8217 14943
rect 8251 14940 8263 14943
rect 8404 14940 8432 15116
rect 8478 15104 8484 15116
rect 8536 15104 8542 15156
rect 9125 15147 9183 15153
rect 9125 15113 9137 15147
rect 9171 15144 9183 15147
rect 9214 15144 9220 15156
rect 9171 15116 9220 15144
rect 9171 15113 9183 15116
rect 9125 15107 9183 15113
rect 9214 15104 9220 15116
rect 9272 15104 9278 15156
rect 10318 15104 10324 15156
rect 10376 15104 10382 15156
rect 12158 15144 12164 15156
rect 11532 15116 12164 15144
rect 10226 15076 10232 15088
rect 8620 15048 10232 15076
rect 8620 15017 8648 15048
rect 10226 15036 10232 15048
rect 10284 15036 10290 15088
rect 11532 15085 11560 15116
rect 12158 15104 12164 15116
rect 12216 15104 12222 15156
rect 12434 15104 12440 15156
rect 12492 15144 12498 15156
rect 12618 15144 12624 15156
rect 12492 15116 12624 15144
rect 12492 15104 12498 15116
rect 12618 15104 12624 15116
rect 12676 15104 12682 15156
rect 14645 15147 14703 15153
rect 14645 15113 14657 15147
rect 14691 15144 14703 15147
rect 15286 15144 15292 15156
rect 14691 15116 15292 15144
rect 14691 15113 14703 15116
rect 14645 15107 14703 15113
rect 15286 15104 15292 15116
rect 15344 15104 15350 15156
rect 16393 15147 16451 15153
rect 16393 15113 16405 15147
rect 16439 15144 16451 15147
rect 20714 15144 20720 15156
rect 16439 15116 20720 15144
rect 16439 15113 16451 15116
rect 16393 15107 16451 15113
rect 11517 15079 11575 15085
rect 11517 15045 11529 15079
rect 11563 15045 11575 15079
rect 11517 15039 11575 15045
rect 12710 15036 12716 15088
rect 12768 15076 12774 15088
rect 12894 15076 12900 15088
rect 12768 15048 12900 15076
rect 12768 15036 12774 15048
rect 12894 15036 12900 15048
rect 12952 15036 12958 15088
rect 13262 15036 13268 15088
rect 13320 15076 13326 15088
rect 13722 15076 13728 15088
rect 13320 15048 13728 15076
rect 13320 15036 13326 15048
rect 13722 15036 13728 15048
rect 13780 15036 13786 15088
rect 15473 15079 15531 15085
rect 15473 15045 15485 15079
rect 15519 15076 15531 15079
rect 15519 15048 15884 15076
rect 15519 15045 15531 15048
rect 15473 15039 15531 15045
rect 8573 15011 8648 15017
rect 8573 14977 8585 15011
rect 8619 14980 8648 15011
rect 8619 14977 8631 14980
rect 8573 14971 8631 14977
rect 9306 14968 9312 15020
rect 9364 14968 9370 15020
rect 10686 15008 10692 15020
rect 9416 14980 10692 15008
rect 9416 14940 9444 14980
rect 8251 14912 9444 14940
rect 9585 14943 9643 14949
rect 8251 14909 8263 14912
rect 8205 14903 8263 14909
rect 9585 14909 9597 14943
rect 9631 14909 9643 14943
rect 9585 14903 9643 14909
rect 6656 14844 7052 14872
rect 6932 14816 6960 14844
rect 7466 14832 7472 14884
rect 7524 14872 7530 14884
rect 7524 14844 8156 14872
rect 7524 14832 7530 14844
rect 4111 14776 5488 14804
rect 4111 14773 4123 14776
rect 4065 14767 4123 14773
rect 5902 14764 5908 14816
rect 5960 14804 5966 14816
rect 5997 14807 6055 14813
rect 5997 14804 6009 14807
rect 5960 14776 6009 14804
rect 5960 14764 5966 14776
rect 5997 14773 6009 14776
rect 6043 14773 6055 14807
rect 5997 14767 6055 14773
rect 6914 14764 6920 14816
rect 6972 14764 6978 14816
rect 7006 14764 7012 14816
rect 7064 14804 7070 14816
rect 7926 14804 7932 14816
rect 7064 14776 7932 14804
rect 7064 14764 7070 14776
rect 7926 14764 7932 14776
rect 7984 14804 7990 14816
rect 8021 14807 8079 14813
rect 8021 14804 8033 14807
rect 7984 14776 8033 14804
rect 7984 14764 7990 14776
rect 8021 14773 8033 14776
rect 8067 14773 8079 14807
rect 8128 14804 8156 14844
rect 9122 14832 9128 14884
rect 9180 14872 9186 14884
rect 9600 14872 9628 14903
rect 10134 14900 10140 14952
rect 10192 14940 10198 14952
rect 10428 14949 10456 14980
rect 10686 14968 10692 14980
rect 10744 14968 10750 15020
rect 11790 14968 11796 15020
rect 11848 14968 11854 15020
rect 11931 15011 11989 15017
rect 11931 14977 11943 15011
rect 11977 15008 11989 15011
rect 13814 15008 13820 15020
rect 11977 14980 13820 15008
rect 11977 14977 11989 14980
rect 11931 14971 11989 14977
rect 10229 14943 10287 14949
rect 10229 14940 10241 14943
rect 10192 14912 10241 14940
rect 10192 14900 10198 14912
rect 10229 14909 10241 14912
rect 10275 14909 10287 14943
rect 10229 14903 10287 14909
rect 10413 14943 10471 14949
rect 10413 14909 10425 14943
rect 10459 14909 10471 14943
rect 10413 14903 10471 14909
rect 10594 14900 10600 14952
rect 10652 14900 10658 14952
rect 10873 14943 10931 14949
rect 10873 14909 10885 14943
rect 10919 14940 10931 14943
rect 10962 14940 10968 14952
rect 10919 14912 10968 14940
rect 10919 14909 10931 14912
rect 10873 14903 10931 14909
rect 10962 14900 10968 14912
rect 11020 14900 11026 14952
rect 11054 14900 11060 14952
rect 11112 14900 11118 14952
rect 12066 14900 12072 14952
rect 12124 14900 12130 14952
rect 9180 14844 9628 14872
rect 9692 14844 11100 14872
rect 9180 14832 9186 14844
rect 8665 14807 8723 14813
rect 8665 14804 8677 14807
rect 8128 14776 8677 14804
rect 8021 14767 8079 14773
rect 8665 14773 8677 14776
rect 8711 14773 8723 14807
rect 8665 14767 8723 14773
rect 8754 14764 8760 14816
rect 8812 14764 8818 14816
rect 9030 14764 9036 14816
rect 9088 14804 9094 14816
rect 9692 14804 9720 14844
rect 9088 14776 9720 14804
rect 9088 14764 9094 14776
rect 10410 14764 10416 14816
rect 10468 14804 10474 14816
rect 10781 14807 10839 14813
rect 10781 14804 10793 14807
rect 10468 14776 10793 14804
rect 10468 14764 10474 14776
rect 10781 14773 10793 14776
rect 10827 14804 10839 14807
rect 10962 14804 10968 14816
rect 10827 14776 10968 14804
rect 10827 14773 10839 14776
rect 10781 14767 10839 14773
rect 10962 14764 10968 14776
rect 11020 14764 11026 14816
rect 11072 14804 11100 14844
rect 12636 14804 12664 14980
rect 13814 14968 13820 14980
rect 13872 14968 13878 15020
rect 15010 15008 15016 15020
rect 14660 14980 15016 15008
rect 12805 14943 12863 14949
rect 12805 14909 12817 14943
rect 12851 14940 12863 14943
rect 12894 14940 12900 14952
rect 12851 14912 12900 14940
rect 12851 14909 12863 14912
rect 12805 14903 12863 14909
rect 12894 14900 12900 14912
rect 12952 14900 12958 14952
rect 12986 14900 12992 14952
rect 13044 14900 13050 14952
rect 13081 14943 13139 14949
rect 13081 14909 13093 14943
rect 13127 14940 13139 14943
rect 13541 14943 13599 14949
rect 13127 14912 13492 14940
rect 13127 14909 13139 14912
rect 13081 14903 13139 14909
rect 11072 14776 12664 14804
rect 12713 14807 12771 14813
rect 12713 14773 12725 14807
rect 12759 14804 12771 14807
rect 12802 14804 12808 14816
rect 12759 14776 12808 14804
rect 12759 14773 12771 14776
rect 12713 14767 12771 14773
rect 12802 14764 12808 14776
rect 12860 14764 12866 14816
rect 12894 14764 12900 14816
rect 12952 14764 12958 14816
rect 13262 14764 13268 14816
rect 13320 14764 13326 14816
rect 13464 14804 13492 14912
rect 13541 14909 13553 14943
rect 13587 14940 13599 14943
rect 13998 14940 14004 14952
rect 13587 14912 14004 14940
rect 13587 14909 13599 14912
rect 13541 14903 13599 14909
rect 13998 14900 14004 14912
rect 14056 14900 14062 14952
rect 14185 14943 14243 14949
rect 14185 14909 14197 14943
rect 14231 14940 14243 14943
rect 14366 14940 14372 14952
rect 14231 14912 14372 14940
rect 14231 14909 14243 14912
rect 14185 14903 14243 14909
rect 14366 14900 14372 14912
rect 14424 14900 14430 14952
rect 13722 14832 13728 14884
rect 13780 14832 13786 14884
rect 13906 14832 13912 14884
rect 13964 14872 13970 14884
rect 14660 14872 14688 14980
rect 15010 14968 15016 14980
rect 15068 14968 15074 15020
rect 14737 14943 14795 14949
rect 14737 14909 14749 14943
rect 14783 14940 14795 14943
rect 14826 14940 14832 14952
rect 14783 14912 14832 14940
rect 14783 14909 14795 14912
rect 14737 14903 14795 14909
rect 14826 14900 14832 14912
rect 14884 14900 14890 14952
rect 15102 14900 15108 14952
rect 15160 14900 15166 14952
rect 15856 14949 15884 15048
rect 15933 15011 15991 15017
rect 15933 14977 15945 15011
rect 15979 15008 15991 15011
rect 16408 15008 16436 15107
rect 20714 15104 20720 15116
rect 20772 15104 20778 15156
rect 16482 15036 16488 15088
rect 16540 15076 16546 15088
rect 16540 15048 16896 15076
rect 16540 15036 16546 15048
rect 15979 14980 16436 15008
rect 16577 15011 16635 15017
rect 15979 14977 15991 14980
rect 15933 14971 15991 14977
rect 16577 14977 16589 15011
rect 16623 15008 16635 15011
rect 16761 15011 16819 15017
rect 16761 15008 16773 15011
rect 16623 14980 16773 15008
rect 16623 14977 16635 14980
rect 16577 14971 16635 14977
rect 16761 14977 16773 14980
rect 16807 14977 16819 15011
rect 16761 14971 16819 14977
rect 16868 14949 16896 15048
rect 18984 15048 19288 15076
rect 18984 15020 19012 15048
rect 17221 15011 17279 15017
rect 17221 14977 17233 15011
rect 17267 15008 17279 15011
rect 17678 15008 17684 15020
rect 17267 14980 17684 15008
rect 17267 14977 17279 14980
rect 17221 14971 17279 14977
rect 17678 14968 17684 14980
rect 17736 14968 17742 15020
rect 18690 14968 18696 15020
rect 18748 15008 18754 15020
rect 18877 15011 18935 15017
rect 18877 15008 18889 15011
rect 18748 14980 18889 15008
rect 18748 14968 18754 14980
rect 18877 14977 18889 14980
rect 18923 14977 18935 15011
rect 18877 14971 18935 14977
rect 18966 14968 18972 15020
rect 19024 14968 19030 15020
rect 19150 14968 19156 15020
rect 19208 14968 19214 15020
rect 19260 15008 19288 15048
rect 19334 15036 19340 15088
rect 19392 15036 19398 15088
rect 19794 15036 19800 15088
rect 19852 15076 19858 15088
rect 19889 15079 19947 15085
rect 19889 15076 19901 15079
rect 19852 15048 19901 15076
rect 19852 15036 19858 15048
rect 19889 15045 19901 15048
rect 19935 15045 19947 15079
rect 19889 15039 19947 15045
rect 19978 15036 19984 15088
rect 20036 15076 20042 15088
rect 20441 15079 20499 15085
rect 20441 15076 20453 15079
rect 20036 15048 20453 15076
rect 20036 15036 20042 15048
rect 20441 15045 20453 15048
rect 20487 15045 20499 15079
rect 20441 15039 20499 15045
rect 19260 14980 21220 15008
rect 15841 14943 15899 14949
rect 15841 14909 15853 14943
rect 15887 14940 15899 14943
rect 16301 14943 16359 14949
rect 16301 14940 16313 14943
rect 15887 14912 16313 14940
rect 15887 14909 15899 14912
rect 15841 14903 15899 14909
rect 16301 14909 16313 14912
rect 16347 14909 16359 14943
rect 16301 14903 16359 14909
rect 16669 14943 16727 14949
rect 16669 14909 16681 14943
rect 16715 14909 16727 14943
rect 16669 14903 16727 14909
rect 16853 14943 16911 14949
rect 16853 14909 16865 14943
rect 16899 14909 16911 14943
rect 16853 14903 16911 14909
rect 13964 14844 14688 14872
rect 15120 14872 15148 14900
rect 16684 14872 16712 14903
rect 17126 14900 17132 14952
rect 17184 14900 17190 14952
rect 18138 14900 18144 14952
rect 18196 14940 18202 14952
rect 19061 14943 19119 14949
rect 19061 14940 19073 14943
rect 18196 14912 19073 14940
rect 18196 14900 18202 14912
rect 19061 14909 19073 14912
rect 19107 14940 19119 14943
rect 19242 14940 19248 14952
rect 19107 14912 19248 14940
rect 19107 14909 19119 14912
rect 19061 14903 19119 14909
rect 19242 14900 19248 14912
rect 19300 14900 19306 14952
rect 19518 14900 19524 14952
rect 19576 14900 19582 14952
rect 20806 14940 20812 14952
rect 19628 14912 20812 14940
rect 15120 14844 16712 14872
rect 13964 14832 13970 14844
rect 19334 14832 19340 14884
rect 19392 14872 19398 14884
rect 19628 14881 19656 14912
rect 20806 14900 20812 14912
rect 20864 14940 20870 14952
rect 20993 14943 21051 14949
rect 20993 14940 21005 14943
rect 20864 14912 21005 14940
rect 20864 14900 20870 14912
rect 20993 14909 21005 14912
rect 21039 14909 21051 14943
rect 20993 14903 21051 14909
rect 19613 14875 19671 14881
rect 19613 14872 19625 14875
rect 19392 14844 19625 14872
rect 19392 14832 19398 14844
rect 19613 14841 19625 14844
rect 19659 14841 19671 14875
rect 19613 14835 19671 14841
rect 19794 14832 19800 14884
rect 19852 14872 19858 14884
rect 20165 14875 20223 14881
rect 20165 14872 20177 14875
rect 19852 14844 20177 14872
rect 19852 14832 19858 14844
rect 20165 14841 20177 14844
rect 20211 14841 20223 14875
rect 20165 14835 20223 14841
rect 14090 14804 14096 14816
rect 13464 14776 14096 14804
rect 14090 14764 14096 14776
rect 14148 14764 14154 14816
rect 14182 14764 14188 14816
rect 14240 14764 14246 14816
rect 14550 14764 14556 14816
rect 14608 14804 14614 14816
rect 15102 14804 15108 14816
rect 14608 14776 15108 14804
rect 14608 14764 14614 14776
rect 15102 14764 15108 14776
rect 15160 14764 15166 14816
rect 16206 14764 16212 14816
rect 16264 14764 16270 14816
rect 16298 14764 16304 14816
rect 16356 14804 16362 14816
rect 16577 14807 16635 14813
rect 16577 14804 16589 14807
rect 16356 14776 16589 14804
rect 16356 14764 16362 14776
rect 16577 14773 16589 14776
rect 16623 14773 16635 14807
rect 16577 14767 16635 14773
rect 17402 14764 17408 14816
rect 17460 14804 17466 14816
rect 17497 14807 17555 14813
rect 17497 14804 17509 14807
rect 17460 14776 17509 14804
rect 17460 14764 17466 14776
rect 17497 14773 17509 14776
rect 17543 14773 17555 14807
rect 17497 14767 17555 14773
rect 18690 14764 18696 14816
rect 18748 14764 18754 14816
rect 19518 14764 19524 14816
rect 19576 14804 19582 14816
rect 19978 14804 19984 14816
rect 19576 14776 19984 14804
rect 19576 14764 19582 14776
rect 19978 14764 19984 14776
rect 20036 14764 20042 14816
rect 20073 14807 20131 14813
rect 20073 14773 20085 14807
rect 20119 14804 20131 14807
rect 20346 14804 20352 14816
rect 20119 14776 20352 14804
rect 20119 14773 20131 14776
rect 20073 14767 20131 14773
rect 20346 14764 20352 14776
rect 20404 14764 20410 14816
rect 20438 14764 20444 14816
rect 20496 14804 20502 14816
rect 21192 14813 21220 14980
rect 22554 14968 22560 15020
rect 22612 14968 22618 15020
rect 22278 14900 22284 14952
rect 22336 14940 22342 14952
rect 22462 14940 22468 14952
rect 22336 14912 22468 14940
rect 22336 14900 22342 14912
rect 22462 14900 22468 14912
rect 22520 14900 22526 14952
rect 20625 14807 20683 14813
rect 20625 14804 20637 14807
rect 20496 14776 20637 14804
rect 20496 14764 20502 14776
rect 20625 14773 20637 14776
rect 20671 14773 20683 14807
rect 20625 14767 20683 14773
rect 21177 14807 21235 14813
rect 21177 14773 21189 14807
rect 21223 14804 21235 14807
rect 21358 14804 21364 14816
rect 21223 14776 21364 14804
rect 21223 14773 21235 14776
rect 21177 14767 21235 14773
rect 21358 14764 21364 14776
rect 21416 14764 21422 14816
rect 21818 14764 21824 14816
rect 21876 14804 21882 14816
rect 22097 14807 22155 14813
rect 22097 14804 22109 14807
rect 21876 14776 22109 14804
rect 21876 14764 21882 14776
rect 22097 14773 22109 14776
rect 22143 14773 22155 14807
rect 22097 14767 22155 14773
rect 552 14714 23368 14736
rect 552 14662 4366 14714
rect 4418 14662 4430 14714
rect 4482 14662 4494 14714
rect 4546 14662 4558 14714
rect 4610 14662 4622 14714
rect 4674 14662 4686 14714
rect 4738 14662 10366 14714
rect 10418 14662 10430 14714
rect 10482 14662 10494 14714
rect 10546 14662 10558 14714
rect 10610 14662 10622 14714
rect 10674 14662 10686 14714
rect 10738 14662 16366 14714
rect 16418 14662 16430 14714
rect 16482 14662 16494 14714
rect 16546 14662 16558 14714
rect 16610 14662 16622 14714
rect 16674 14662 16686 14714
rect 16738 14662 22366 14714
rect 22418 14662 22430 14714
rect 22482 14662 22494 14714
rect 22546 14662 22558 14714
rect 22610 14662 22622 14714
rect 22674 14662 22686 14714
rect 22738 14662 23368 14714
rect 552 14640 23368 14662
rect 1397 14603 1455 14609
rect 1397 14569 1409 14603
rect 1443 14600 1455 14603
rect 1854 14600 1860 14612
rect 1443 14572 1860 14600
rect 1443 14569 1455 14572
rect 1397 14563 1455 14569
rect 1854 14560 1860 14572
rect 1912 14560 1918 14612
rect 3418 14560 3424 14612
rect 3476 14560 3482 14612
rect 3973 14603 4031 14609
rect 3973 14569 3985 14603
rect 4019 14600 4031 14603
rect 4062 14600 4068 14612
rect 4019 14572 4068 14600
rect 4019 14569 4031 14572
rect 3973 14563 4031 14569
rect 4062 14560 4068 14572
rect 4120 14560 4126 14612
rect 4246 14560 4252 14612
rect 4304 14560 4310 14612
rect 4890 14560 4896 14612
rect 4948 14600 4954 14612
rect 6178 14600 6184 14612
rect 4948 14572 6184 14600
rect 4948 14560 4954 14572
rect 6178 14560 6184 14572
rect 6236 14560 6242 14612
rect 6546 14560 6552 14612
rect 6604 14600 6610 14612
rect 7561 14603 7619 14609
rect 7561 14600 7573 14603
rect 6604 14572 7573 14600
rect 6604 14560 6610 14572
rect 7561 14569 7573 14572
rect 7607 14569 7619 14603
rect 7561 14563 7619 14569
rect 8386 14560 8392 14612
rect 8444 14600 8450 14612
rect 8481 14603 8539 14609
rect 8481 14600 8493 14603
rect 8444 14572 8493 14600
rect 8444 14560 8450 14572
rect 8481 14569 8493 14572
rect 8527 14569 8539 14603
rect 8481 14563 8539 14569
rect 9033 14603 9091 14609
rect 9033 14569 9045 14603
rect 9079 14569 9091 14603
rect 9033 14563 9091 14569
rect 1305 14535 1363 14541
rect 1305 14501 1317 14535
rect 1351 14532 1363 14535
rect 1762 14532 1768 14544
rect 1351 14504 1768 14532
rect 1351 14501 1363 14504
rect 1305 14495 1363 14501
rect 1762 14492 1768 14504
rect 1820 14492 1826 14544
rect 2590 14532 2596 14544
rect 1964 14504 2596 14532
rect 1026 14424 1032 14476
rect 1084 14424 1090 14476
rect 1118 14424 1124 14476
rect 1176 14424 1182 14476
rect 1578 14424 1584 14476
rect 1636 14464 1642 14476
rect 1964 14464 1992 14504
rect 1636 14436 1992 14464
rect 1636 14424 1642 14436
rect 2038 14424 2044 14476
rect 2096 14424 2102 14476
rect 2332 14473 2360 14504
rect 2590 14492 2596 14504
rect 2648 14492 2654 14544
rect 3694 14492 3700 14544
rect 3752 14532 3758 14544
rect 4798 14532 4804 14544
rect 3752 14504 4804 14532
rect 3752 14492 3758 14504
rect 4798 14492 4804 14504
rect 4856 14532 4862 14544
rect 4985 14535 5043 14541
rect 4985 14532 4997 14535
rect 4856 14504 4997 14532
rect 4856 14492 4862 14504
rect 4985 14501 4997 14504
rect 5031 14501 5043 14535
rect 4985 14495 5043 14501
rect 5353 14535 5411 14541
rect 5353 14501 5365 14535
rect 5399 14532 5411 14535
rect 5442 14532 5448 14544
rect 5399 14504 5448 14532
rect 5399 14501 5411 14504
rect 5353 14495 5411 14501
rect 5442 14492 5448 14504
rect 5500 14492 5506 14544
rect 6730 14492 6736 14544
rect 6788 14532 6794 14544
rect 6788 14504 7236 14532
rect 6788 14492 6794 14504
rect 2317 14467 2375 14473
rect 2317 14433 2329 14467
rect 2363 14433 2375 14467
rect 2317 14427 2375 14433
rect 2958 14424 2964 14476
rect 3016 14424 3022 14476
rect 3142 14424 3148 14476
rect 3200 14464 3206 14476
rect 3605 14467 3663 14473
rect 3605 14464 3617 14467
rect 3200 14436 3617 14464
rect 3200 14424 3206 14436
rect 3605 14433 3617 14436
rect 3651 14433 3663 14467
rect 3605 14427 3663 14433
rect 3789 14467 3847 14473
rect 3789 14433 3801 14467
rect 3835 14464 3847 14467
rect 3878 14464 3884 14476
rect 3835 14436 3884 14464
rect 3835 14433 3847 14436
rect 3789 14427 3847 14433
rect 3878 14424 3884 14436
rect 3936 14424 3942 14476
rect 4522 14424 4528 14476
rect 4580 14424 4586 14476
rect 4614 14424 4620 14476
rect 4672 14424 4678 14476
rect 5166 14424 5172 14476
rect 5224 14464 5230 14476
rect 6086 14464 6092 14476
rect 5224 14436 6092 14464
rect 5224 14424 5230 14436
rect 6086 14424 6092 14436
rect 6144 14424 6150 14476
rect 7009 14467 7067 14473
rect 7009 14433 7021 14467
rect 7055 14464 7067 14467
rect 7098 14464 7104 14476
rect 7055 14436 7104 14464
rect 7055 14433 7067 14436
rect 7009 14427 7067 14433
rect 7098 14424 7104 14436
rect 7156 14424 7162 14476
rect 7208 14464 7236 14504
rect 7926 14492 7932 14544
rect 7984 14492 7990 14544
rect 9048 14532 9076 14563
rect 9214 14560 9220 14612
rect 9272 14600 9278 14612
rect 10042 14600 10048 14612
rect 9272 14572 10048 14600
rect 9272 14560 9278 14572
rect 10042 14560 10048 14572
rect 10100 14560 10106 14612
rect 11054 14560 11060 14612
rect 11112 14600 11118 14612
rect 11333 14603 11391 14609
rect 11333 14600 11345 14603
rect 11112 14572 11345 14600
rect 11112 14560 11118 14572
rect 11333 14569 11345 14572
rect 11379 14600 11391 14603
rect 12250 14600 12256 14612
rect 11379 14572 12256 14600
rect 11379 14569 11391 14572
rect 11333 14563 11391 14569
rect 12250 14560 12256 14572
rect 12308 14560 12314 14612
rect 12802 14600 12808 14612
rect 12636 14572 12808 14600
rect 9306 14532 9312 14544
rect 8588 14504 9312 14532
rect 7466 14464 7472 14476
rect 7208 14436 7472 14464
rect 7451 14434 7472 14436
rect 7466 14424 7472 14434
rect 7524 14424 7530 14476
rect 7745 14467 7803 14473
rect 7745 14433 7757 14467
rect 7791 14464 7803 14467
rect 8202 14464 8208 14476
rect 7791 14436 8208 14464
rect 7791 14433 7803 14436
rect 7745 14427 7803 14433
rect 8202 14424 8208 14436
rect 8260 14424 8266 14476
rect 8389 14467 8447 14473
rect 8389 14433 8401 14467
rect 8435 14464 8447 14467
rect 8478 14464 8484 14476
rect 8435 14436 8484 14464
rect 8435 14433 8447 14436
rect 8389 14427 8447 14433
rect 8478 14424 8484 14436
rect 8536 14424 8542 14476
rect 8588 14473 8616 14504
rect 9306 14492 9312 14504
rect 9364 14532 9370 14544
rect 10594 14532 10600 14544
rect 9364 14504 9812 14532
rect 9364 14492 9370 14504
rect 8573 14467 8631 14473
rect 8573 14433 8585 14467
rect 8619 14433 8631 14467
rect 8573 14427 8631 14433
rect 8665 14467 8723 14473
rect 8665 14433 8677 14467
rect 8711 14464 8723 14467
rect 8754 14464 8760 14476
rect 8711 14436 8760 14464
rect 8711 14433 8723 14436
rect 8665 14427 8723 14433
rect 8754 14424 8760 14436
rect 8812 14424 8818 14476
rect 8846 14424 8852 14476
rect 8904 14424 8910 14476
rect 9214 14424 9220 14476
rect 9272 14424 9278 14476
rect 9398 14424 9404 14476
rect 9456 14424 9462 14476
rect 9582 14424 9588 14476
rect 9640 14424 9646 14476
rect 9674 14424 9680 14476
rect 9732 14424 9738 14476
rect 9784 14473 9812 14504
rect 10152 14504 10600 14532
rect 9769 14467 9827 14473
rect 9769 14433 9781 14467
rect 9815 14433 9827 14467
rect 9769 14427 9827 14433
rect 10042 14424 10048 14476
rect 10100 14464 10106 14476
rect 10152 14473 10180 14504
rect 10594 14492 10600 14504
rect 10652 14492 10658 14544
rect 12161 14535 12219 14541
rect 12161 14501 12173 14535
rect 12207 14532 12219 14535
rect 12636 14532 12664 14572
rect 12802 14560 12808 14572
rect 12860 14560 12866 14612
rect 13170 14560 13176 14612
rect 13228 14600 13234 14612
rect 13630 14600 13636 14612
rect 13228 14572 13636 14600
rect 13228 14560 13234 14572
rect 13630 14560 13636 14572
rect 13688 14560 13694 14612
rect 17310 14560 17316 14612
rect 17368 14600 17374 14612
rect 17405 14603 17463 14609
rect 17405 14600 17417 14603
rect 17368 14572 17417 14600
rect 17368 14560 17374 14572
rect 17405 14569 17417 14572
rect 17451 14569 17463 14603
rect 17405 14563 17463 14569
rect 17678 14560 17684 14612
rect 17736 14560 17742 14612
rect 19242 14560 19248 14612
rect 19300 14600 19306 14612
rect 21266 14600 21272 14612
rect 19300 14572 21272 14600
rect 19300 14560 19306 14572
rect 21266 14560 21272 14572
rect 21324 14560 21330 14612
rect 12207 14504 12664 14532
rect 12207 14501 12219 14504
rect 12161 14495 12219 14501
rect 12710 14492 12716 14544
rect 12768 14532 12774 14544
rect 13725 14535 13783 14541
rect 13725 14532 13737 14535
rect 12768 14504 13737 14532
rect 12768 14492 12774 14504
rect 13725 14501 13737 14504
rect 13771 14501 13783 14535
rect 13725 14495 13783 14501
rect 14734 14492 14740 14544
rect 14792 14532 14798 14544
rect 18690 14532 18696 14544
rect 14792 14504 18696 14532
rect 14792 14492 14798 14504
rect 18690 14492 18696 14504
rect 18748 14492 18754 14544
rect 21358 14492 21364 14544
rect 21416 14492 21422 14544
rect 10137 14467 10195 14473
rect 10137 14464 10149 14467
rect 10100 14436 10149 14464
rect 10100 14424 10106 14436
rect 10137 14433 10149 14436
rect 10183 14433 10195 14467
rect 10137 14427 10195 14433
rect 10321 14467 10379 14473
rect 10321 14433 10333 14467
rect 10367 14464 10379 14467
rect 10962 14464 10968 14476
rect 10367 14436 10968 14464
rect 10367 14433 10379 14436
rect 10321 14427 10379 14433
rect 10962 14424 10968 14436
rect 11020 14424 11026 14476
rect 11517 14467 11575 14473
rect 11517 14433 11529 14467
rect 11563 14464 11575 14467
rect 11698 14464 11704 14476
rect 11563 14436 11704 14464
rect 11563 14433 11575 14436
rect 11517 14427 11575 14433
rect 11698 14424 11704 14436
rect 11756 14424 11762 14476
rect 11790 14424 11796 14476
rect 11848 14424 11854 14476
rect 12342 14424 12348 14476
rect 12400 14464 12406 14476
rect 12618 14464 12624 14476
rect 12400 14436 12624 14464
rect 12400 14424 12406 14436
rect 12618 14424 12624 14436
rect 12676 14424 12682 14476
rect 12802 14424 12808 14476
rect 12860 14424 12866 14476
rect 13262 14464 13268 14476
rect 13004 14436 13268 14464
rect 2406 14356 2412 14408
rect 2464 14356 2470 14408
rect 2866 14356 2872 14408
rect 2924 14356 2930 14408
rect 5813 14399 5871 14405
rect 5813 14396 5825 14399
rect 5290 14368 5825 14396
rect 5813 14365 5825 14368
rect 5859 14365 5871 14399
rect 5813 14359 5871 14365
rect 7193 14399 7251 14405
rect 7193 14365 7205 14399
rect 7239 14396 7251 14399
rect 9950 14396 9956 14408
rect 7239 14368 9956 14396
rect 7239 14365 7251 14368
rect 7193 14359 7251 14365
rect 2685 14331 2743 14337
rect 2685 14297 2697 14331
rect 2731 14328 2743 14331
rect 3510 14328 3516 14340
rect 2731 14300 3516 14328
rect 2731 14297 2743 14300
rect 2685 14291 2743 14297
rect 3510 14288 3516 14300
rect 3568 14288 3574 14340
rect 5828 14328 5856 14359
rect 9950 14356 9956 14368
rect 10008 14356 10014 14408
rect 10410 14356 10416 14408
rect 10468 14396 10474 14408
rect 11606 14396 11612 14408
rect 10468 14368 11612 14396
rect 10468 14356 10474 14368
rect 11606 14356 11612 14368
rect 11664 14356 11670 14408
rect 12066 14356 12072 14408
rect 12124 14356 12130 14408
rect 12434 14356 12440 14408
rect 12492 14396 12498 14408
rect 13004 14396 13032 14436
rect 13262 14424 13268 14436
rect 13320 14424 13326 14476
rect 13998 14424 14004 14476
rect 14056 14424 14062 14476
rect 14182 14424 14188 14476
rect 14240 14464 14246 14476
rect 14645 14467 14703 14473
rect 14645 14464 14657 14467
rect 14240 14436 14657 14464
rect 14240 14424 14246 14436
rect 14645 14433 14657 14436
rect 14691 14433 14703 14467
rect 14645 14427 14703 14433
rect 15010 14424 15016 14476
rect 15068 14464 15074 14476
rect 15289 14467 15347 14473
rect 15289 14464 15301 14467
rect 15068 14436 15301 14464
rect 15068 14424 15074 14436
rect 15289 14433 15301 14436
rect 15335 14433 15347 14467
rect 15289 14427 15347 14433
rect 17589 14467 17647 14473
rect 17589 14433 17601 14467
rect 17635 14433 17647 14467
rect 17589 14427 17647 14433
rect 12492 14368 13032 14396
rect 13081 14399 13139 14405
rect 12492 14356 12498 14368
rect 13081 14365 13093 14399
rect 13127 14396 13139 14399
rect 13170 14396 13176 14408
rect 13127 14368 13176 14396
rect 13127 14365 13139 14368
rect 13081 14359 13139 14365
rect 13170 14356 13176 14368
rect 13228 14356 13234 14408
rect 13909 14399 13967 14405
rect 13909 14365 13921 14399
rect 13955 14365 13967 14399
rect 13909 14359 13967 14365
rect 10134 14328 10140 14340
rect 5828 14300 10140 14328
rect 10134 14288 10140 14300
rect 10192 14288 10198 14340
rect 10318 14288 10324 14340
rect 10376 14328 10382 14340
rect 13924 14328 13952 14359
rect 14366 14356 14372 14408
rect 14424 14356 14430 14408
rect 14737 14399 14795 14405
rect 14737 14365 14749 14399
rect 14783 14365 14795 14399
rect 14737 14359 14795 14365
rect 14752 14328 14780 14359
rect 14918 14356 14924 14408
rect 14976 14396 14982 14408
rect 15105 14399 15163 14405
rect 15105 14396 15117 14399
rect 14976 14368 15117 14396
rect 14976 14356 14982 14368
rect 15105 14365 15117 14368
rect 15151 14365 15163 14399
rect 15105 14359 15163 14365
rect 16758 14328 16764 14340
rect 10376 14300 13860 14328
rect 13924 14300 16764 14328
rect 10376 14288 10382 14300
rect 1854 14220 1860 14272
rect 1912 14220 1918 14272
rect 3142 14220 3148 14272
rect 3200 14260 3206 14272
rect 3237 14263 3295 14269
rect 3237 14260 3249 14263
rect 3200 14232 3249 14260
rect 3200 14220 3206 14232
rect 3237 14229 3249 14232
rect 3283 14229 3295 14263
rect 3237 14223 3295 14229
rect 5534 14220 5540 14272
rect 5592 14220 5598 14272
rect 6825 14263 6883 14269
rect 6825 14229 6837 14263
rect 6871 14260 6883 14263
rect 7006 14260 7012 14272
rect 6871 14232 7012 14260
rect 6871 14229 6883 14232
rect 6825 14223 6883 14229
rect 7006 14220 7012 14232
rect 7064 14220 7070 14272
rect 8386 14220 8392 14272
rect 8444 14260 8450 14272
rect 9766 14260 9772 14272
rect 8444 14232 9772 14260
rect 8444 14220 8450 14232
rect 9766 14220 9772 14232
rect 9824 14220 9830 14272
rect 9950 14220 9956 14272
rect 10008 14260 10014 14272
rect 10045 14263 10103 14269
rect 10045 14260 10057 14263
rect 10008 14232 10057 14260
rect 10008 14220 10014 14232
rect 10045 14229 10057 14232
rect 10091 14229 10103 14263
rect 10045 14223 10103 14229
rect 10229 14263 10287 14269
rect 10229 14229 10241 14263
rect 10275 14260 10287 14263
rect 10502 14260 10508 14272
rect 10275 14232 10508 14260
rect 10275 14229 10287 14232
rect 10229 14223 10287 14229
rect 10502 14220 10508 14232
rect 10560 14260 10566 14272
rect 10778 14260 10784 14272
rect 10560 14232 10784 14260
rect 10560 14220 10566 14232
rect 10778 14220 10784 14232
rect 10836 14220 10842 14272
rect 11054 14220 11060 14272
rect 11112 14260 11118 14272
rect 11330 14260 11336 14272
rect 11112 14232 11336 14260
rect 11112 14220 11118 14232
rect 11330 14220 11336 14232
rect 11388 14260 11394 14272
rect 11609 14263 11667 14269
rect 11609 14260 11621 14263
rect 11388 14232 11621 14260
rect 11388 14220 11394 14232
rect 11609 14229 11621 14232
rect 11655 14229 11667 14263
rect 11609 14223 11667 14229
rect 12618 14220 12624 14272
rect 12676 14220 12682 14272
rect 13832 14260 13860 14300
rect 16758 14288 16764 14300
rect 16816 14288 16822 14340
rect 17126 14288 17132 14340
rect 17184 14328 17190 14340
rect 17604 14328 17632 14427
rect 17678 14424 17684 14476
rect 17736 14424 17742 14476
rect 17865 14467 17923 14473
rect 17865 14433 17877 14467
rect 17911 14464 17923 14467
rect 18414 14464 18420 14476
rect 17911 14436 18420 14464
rect 17911 14433 17923 14436
rect 17865 14427 17923 14433
rect 18414 14424 18420 14436
rect 18472 14464 18478 14476
rect 18966 14464 18972 14476
rect 18472 14436 18972 14464
rect 18472 14424 18478 14436
rect 18966 14424 18972 14436
rect 19024 14424 19030 14476
rect 19978 14464 19984 14476
rect 19076 14436 19984 14464
rect 18690 14356 18696 14408
rect 18748 14396 18754 14408
rect 19076 14405 19104 14436
rect 19978 14424 19984 14436
rect 20036 14424 20042 14476
rect 20165 14467 20223 14473
rect 20165 14433 20177 14467
rect 20211 14433 20223 14467
rect 20165 14427 20223 14433
rect 19061 14399 19119 14405
rect 19061 14396 19073 14399
rect 18748 14368 19073 14396
rect 18748 14356 18754 14368
rect 19061 14365 19073 14368
rect 19107 14365 19119 14399
rect 19061 14359 19119 14365
rect 19334 14356 19340 14408
rect 19392 14356 19398 14408
rect 19886 14356 19892 14408
rect 19944 14396 19950 14408
rect 20180 14396 20208 14427
rect 20346 14424 20352 14476
rect 20404 14424 20410 14476
rect 20438 14424 20444 14476
rect 20496 14424 20502 14476
rect 21174 14424 21180 14476
rect 21232 14464 21238 14476
rect 21545 14467 21603 14473
rect 21545 14464 21557 14467
rect 21232 14436 21557 14464
rect 21232 14424 21238 14436
rect 21545 14433 21557 14436
rect 21591 14464 21603 14467
rect 21910 14464 21916 14476
rect 21591 14436 21916 14464
rect 21591 14433 21603 14436
rect 21545 14427 21603 14433
rect 21910 14424 21916 14436
rect 21968 14424 21974 14476
rect 22002 14424 22008 14476
rect 22060 14424 22066 14476
rect 22097 14467 22155 14473
rect 22097 14433 22109 14467
rect 22143 14433 22155 14467
rect 22097 14427 22155 14433
rect 19944 14368 20208 14396
rect 21729 14399 21787 14405
rect 19944 14356 19950 14368
rect 21729 14365 21741 14399
rect 21775 14396 21787 14399
rect 22112 14396 22140 14427
rect 22278 14424 22284 14476
rect 22336 14424 22342 14476
rect 21775 14368 22140 14396
rect 21775 14365 21787 14368
rect 21729 14359 21787 14365
rect 19242 14328 19248 14340
rect 17184 14300 19248 14328
rect 17184 14288 17190 14300
rect 19242 14288 19248 14300
rect 19300 14288 19306 14340
rect 14550 14260 14556 14272
rect 13832 14232 14556 14260
rect 14550 14220 14556 14232
rect 14608 14220 14614 14272
rect 14826 14220 14832 14272
rect 14884 14260 14890 14272
rect 15013 14263 15071 14269
rect 15013 14260 15025 14263
rect 14884 14232 15025 14260
rect 14884 14220 14890 14232
rect 15013 14229 15025 14232
rect 15059 14229 15071 14263
rect 15013 14223 15071 14229
rect 15102 14220 15108 14272
rect 15160 14260 15166 14272
rect 15473 14263 15531 14269
rect 15473 14260 15485 14263
rect 15160 14232 15485 14260
rect 15160 14220 15166 14232
rect 15473 14229 15485 14232
rect 15519 14229 15531 14263
rect 15473 14223 15531 14229
rect 15838 14220 15844 14272
rect 15896 14260 15902 14272
rect 19518 14260 19524 14272
rect 15896 14232 19524 14260
rect 15896 14220 15902 14232
rect 19518 14220 19524 14232
rect 19576 14220 19582 14272
rect 19981 14263 20039 14269
rect 19981 14229 19993 14263
rect 20027 14260 20039 14263
rect 20438 14260 20444 14272
rect 20027 14232 20444 14260
rect 20027 14229 20039 14232
rect 19981 14223 20039 14229
rect 20438 14220 20444 14232
rect 20496 14220 20502 14272
rect 21634 14220 21640 14272
rect 21692 14260 21698 14272
rect 21821 14263 21879 14269
rect 21821 14260 21833 14263
rect 21692 14232 21833 14260
rect 21692 14220 21698 14232
rect 21821 14229 21833 14232
rect 21867 14229 21879 14263
rect 21821 14223 21879 14229
rect 22189 14263 22247 14269
rect 22189 14229 22201 14263
rect 22235 14260 22247 14263
rect 22462 14260 22468 14272
rect 22235 14232 22468 14260
rect 22235 14229 22247 14232
rect 22189 14223 22247 14229
rect 22462 14220 22468 14232
rect 22520 14220 22526 14272
rect 552 14170 23368 14192
rect 552 14118 1366 14170
rect 1418 14118 1430 14170
rect 1482 14118 1494 14170
rect 1546 14118 1558 14170
rect 1610 14118 1622 14170
rect 1674 14118 1686 14170
rect 1738 14118 7366 14170
rect 7418 14118 7430 14170
rect 7482 14118 7494 14170
rect 7546 14118 7558 14170
rect 7610 14118 7622 14170
rect 7674 14118 7686 14170
rect 7738 14118 13366 14170
rect 13418 14118 13430 14170
rect 13482 14118 13494 14170
rect 13546 14118 13558 14170
rect 13610 14118 13622 14170
rect 13674 14118 13686 14170
rect 13738 14118 19366 14170
rect 19418 14118 19430 14170
rect 19482 14118 19494 14170
rect 19546 14118 19558 14170
rect 19610 14118 19622 14170
rect 19674 14118 19686 14170
rect 19738 14118 23368 14170
rect 552 14096 23368 14118
rect 2958 14016 2964 14068
rect 3016 14016 3022 14068
rect 4062 14016 4068 14068
rect 4120 14016 4126 14068
rect 5997 14059 6055 14065
rect 5997 14025 6009 14059
rect 6043 14056 6055 14059
rect 6822 14056 6828 14068
rect 6043 14028 6828 14056
rect 6043 14025 6055 14028
rect 5997 14019 6055 14025
rect 6822 14016 6828 14028
rect 6880 14016 6886 14068
rect 9766 14016 9772 14068
rect 9824 14056 9830 14068
rect 10410 14056 10416 14068
rect 9824 14028 10416 14056
rect 9824 14016 9830 14028
rect 10410 14016 10416 14028
rect 10468 14016 10474 14068
rect 10781 14059 10839 14065
rect 10781 14025 10793 14059
rect 10827 14056 10839 14059
rect 12342 14056 12348 14068
rect 10827 14028 12348 14056
rect 10827 14025 10839 14028
rect 10781 14019 10839 14025
rect 12342 14016 12348 14028
rect 12400 14016 12406 14068
rect 12529 14059 12587 14065
rect 12529 14025 12541 14059
rect 12575 14056 12587 14059
rect 12802 14056 12808 14068
rect 12575 14028 12808 14056
rect 12575 14025 12587 14028
rect 12529 14019 12587 14025
rect 12802 14016 12808 14028
rect 12860 14056 12866 14068
rect 13354 14056 13360 14068
rect 12860 14028 13360 14056
rect 12860 14016 12866 14028
rect 13354 14016 13360 14028
rect 13412 14016 13418 14068
rect 13909 14059 13967 14065
rect 13909 14025 13921 14059
rect 13955 14056 13967 14059
rect 14366 14056 14372 14068
rect 13955 14028 14372 14056
rect 13955 14025 13967 14028
rect 13909 14019 13967 14025
rect 14366 14016 14372 14028
rect 14424 14016 14430 14068
rect 15470 14016 15476 14068
rect 15528 14056 15534 14068
rect 15528 14028 17264 14056
rect 15528 14016 15534 14028
rect 2682 13948 2688 14000
rect 2740 13988 2746 14000
rect 2869 13991 2927 13997
rect 2869 13988 2881 13991
rect 2740 13960 2881 13988
rect 2740 13948 2746 13960
rect 2869 13957 2881 13960
rect 2915 13988 2927 13991
rect 4080 13988 4108 14016
rect 2915 13960 4108 13988
rect 2915 13957 2927 13960
rect 2869 13951 2927 13957
rect 4522 13948 4528 14000
rect 4580 13988 4586 14000
rect 5074 13988 5080 14000
rect 4580 13960 5080 13988
rect 4580 13948 4586 13960
rect 5074 13948 5080 13960
rect 5132 13948 5138 14000
rect 8110 13948 8116 14000
rect 8168 13948 8174 14000
rect 9861 13991 9919 13997
rect 9861 13957 9873 13991
rect 9907 13988 9919 13991
rect 10686 13988 10692 14000
rect 9907 13960 10692 13988
rect 9907 13957 9919 13960
rect 9861 13951 9919 13957
rect 10686 13948 10692 13960
rect 10744 13948 10750 14000
rect 10965 13991 11023 13997
rect 10965 13957 10977 13991
rect 11011 13988 11023 13991
rect 11238 13988 11244 14000
rect 11011 13960 11244 13988
rect 11011 13957 11023 13960
rect 10965 13951 11023 13957
rect 11238 13948 11244 13960
rect 11296 13948 11302 14000
rect 11790 13948 11796 14000
rect 11848 13988 11854 14000
rect 13081 13991 13139 13997
rect 13081 13988 13093 13991
rect 11848 13960 13093 13988
rect 11848 13948 11854 13960
rect 13081 13957 13093 13960
rect 13127 13957 13139 13991
rect 13081 13951 13139 13957
rect 13725 13991 13783 13997
rect 13725 13957 13737 13991
rect 13771 13988 13783 13991
rect 16761 13991 16819 13997
rect 13771 13960 16712 13988
rect 13771 13957 13783 13960
rect 13725 13951 13783 13957
rect 3050 13880 3056 13932
rect 3108 13880 3114 13932
rect 842 13812 848 13864
rect 900 13852 906 13864
rect 1118 13852 1124 13864
rect 900 13824 1124 13852
rect 900 13812 906 13824
rect 1118 13812 1124 13824
rect 1176 13812 1182 13864
rect 1210 13812 1216 13864
rect 1268 13852 1274 13864
rect 1305 13855 1363 13861
rect 1305 13852 1317 13855
rect 1268 13824 1317 13852
rect 1268 13812 1274 13824
rect 1305 13821 1317 13824
rect 1351 13821 1363 13855
rect 1305 13815 1363 13821
rect 1572 13855 1630 13861
rect 1572 13821 1584 13855
rect 1618 13852 1630 13855
rect 1854 13852 1860 13864
rect 1618 13824 1860 13852
rect 1618 13821 1630 13824
rect 1572 13815 1630 13821
rect 1854 13812 1860 13824
rect 1912 13812 1918 13864
rect 2777 13855 2835 13861
rect 2777 13821 2789 13855
rect 2823 13821 2835 13855
rect 2777 13815 2835 13821
rect 1026 13744 1032 13796
rect 1084 13784 1090 13796
rect 2406 13784 2412 13796
rect 1084 13756 2412 13784
rect 1084 13744 1090 13756
rect 2406 13744 2412 13756
rect 2464 13784 2470 13796
rect 2792 13784 2820 13815
rect 3602 13812 3608 13864
rect 3660 13852 3666 13864
rect 3697 13855 3755 13861
rect 3697 13852 3709 13855
rect 3660 13824 3709 13852
rect 3660 13812 3666 13824
rect 3697 13821 3709 13824
rect 3743 13821 3755 13855
rect 3697 13815 3755 13821
rect 3881 13855 3939 13861
rect 3881 13821 3893 13855
rect 3927 13852 3939 13855
rect 3970 13852 3976 13864
rect 3927 13824 3976 13852
rect 3927 13821 3939 13824
rect 3881 13815 3939 13821
rect 3970 13812 3976 13824
rect 4028 13812 4034 13864
rect 5074 13812 5080 13864
rect 5132 13852 5138 13864
rect 5813 13855 5871 13861
rect 5813 13852 5825 13855
rect 5132 13824 5825 13852
rect 5132 13812 5138 13824
rect 5813 13821 5825 13824
rect 5859 13852 5871 13855
rect 7193 13855 7251 13861
rect 5859 13824 6776 13852
rect 5859 13821 5871 13824
rect 5813 13815 5871 13821
rect 2464 13756 2820 13784
rect 6748 13784 6776 13824
rect 7193 13821 7205 13855
rect 7239 13852 7251 13855
rect 7374 13852 7380 13864
rect 7239 13824 7380 13852
rect 7239 13821 7251 13824
rect 7193 13815 7251 13821
rect 7374 13812 7380 13824
rect 7432 13812 7438 13864
rect 7650 13812 7656 13864
rect 7708 13852 7714 13864
rect 7852 13852 7880 13906
rect 8754 13880 8760 13932
rect 8812 13880 8818 13932
rect 12161 13923 12219 13929
rect 12161 13920 12173 13923
rect 9683 13892 12173 13920
rect 8772 13852 8800 13880
rect 7708 13824 8800 13852
rect 7708 13812 7714 13824
rect 8938 13812 8944 13864
rect 8996 13812 9002 13864
rect 9398 13812 9404 13864
rect 9456 13852 9462 13864
rect 9683 13854 9711 13892
rect 12161 13889 12173 13892
rect 12207 13889 12219 13923
rect 12986 13920 12992 13932
rect 12161 13883 12219 13889
rect 12360 13892 12992 13920
rect 9600 13852 9711 13854
rect 9456 13826 9711 13852
rect 10137 13855 10195 13861
rect 9456 13824 9628 13826
rect 9456 13812 9462 13824
rect 10137 13821 10149 13855
rect 10183 13852 10195 13855
rect 10183 13821 10196 13852
rect 10137 13815 10196 13821
rect 7101 13787 7159 13793
rect 7101 13784 7113 13787
rect 6748 13756 7113 13784
rect 2464 13744 2470 13756
rect 7101 13753 7113 13756
rect 7147 13753 7159 13787
rect 7101 13747 7159 13753
rect 7558 13744 7564 13796
rect 7616 13784 7622 13796
rect 8849 13787 8907 13793
rect 8849 13784 8861 13787
rect 7616 13756 8861 13784
rect 7616 13744 7622 13756
rect 8849 13753 8861 13756
rect 8895 13753 8907 13787
rect 8849 13747 8907 13753
rect 9306 13744 9312 13796
rect 9364 13744 9370 13796
rect 9677 13787 9735 13793
rect 9677 13753 9689 13787
rect 9723 13784 9735 13787
rect 9766 13784 9772 13796
rect 9723 13756 9772 13784
rect 9723 13753 9735 13756
rect 9677 13747 9735 13753
rect 9766 13744 9772 13756
rect 9824 13744 9830 13796
rect 10168 13784 10196 13815
rect 10226 13812 10232 13864
rect 10284 13852 10290 13864
rect 10413 13855 10471 13861
rect 10413 13852 10425 13855
rect 10284 13824 10425 13852
rect 10284 13812 10290 13824
rect 10413 13821 10425 13824
rect 10459 13821 10471 13855
rect 10781 13855 10839 13861
rect 10781 13852 10793 13855
rect 10413 13815 10471 13821
rect 10520 13824 10793 13852
rect 10520 13784 10548 13824
rect 10781 13821 10793 13824
rect 10827 13821 10839 13855
rect 10781 13815 10839 13821
rect 11609 13855 11667 13861
rect 11609 13821 11621 13855
rect 11655 13821 11667 13855
rect 11609 13815 11667 13821
rect 10168 13756 10548 13784
rect 10244 13728 10272 13756
rect 10594 13744 10600 13796
rect 10652 13784 10658 13796
rect 11330 13784 11336 13796
rect 10652 13756 11336 13784
rect 10652 13744 10658 13756
rect 11330 13744 11336 13756
rect 11388 13744 11394 13796
rect 11624 13784 11652 13815
rect 11698 13812 11704 13864
rect 11756 13852 11762 13864
rect 12360 13861 12388 13892
rect 12986 13880 12992 13892
rect 13044 13880 13050 13932
rect 13740 13920 13768 13951
rect 15381 13923 15439 13929
rect 15381 13920 15393 13923
rect 13188 13892 13768 13920
rect 14660 13892 15056 13920
rect 11885 13855 11943 13861
rect 11885 13852 11897 13855
rect 11756 13824 11897 13852
rect 11756 13812 11762 13824
rect 11885 13821 11897 13824
rect 11931 13821 11943 13855
rect 11885 13815 11943 13821
rect 12345 13855 12403 13861
rect 12345 13821 12357 13855
rect 12391 13821 12403 13855
rect 12345 13815 12403 13821
rect 12621 13855 12679 13861
rect 12621 13821 12633 13855
rect 12667 13852 12679 13855
rect 12802 13852 12808 13864
rect 12667 13824 12808 13852
rect 12667 13821 12679 13824
rect 12621 13815 12679 13821
rect 12802 13812 12808 13824
rect 12860 13812 12866 13864
rect 12897 13855 12955 13861
rect 12897 13821 12909 13855
rect 12943 13852 12955 13855
rect 13188 13852 13216 13892
rect 12943 13824 13216 13852
rect 12943 13821 12955 13824
rect 12897 13815 12955 13821
rect 13262 13812 13268 13864
rect 13320 13852 13326 13864
rect 13357 13855 13415 13861
rect 13357 13852 13369 13855
rect 13320 13824 13369 13852
rect 13320 13812 13326 13824
rect 13357 13821 13369 13824
rect 13403 13852 13415 13855
rect 13541 13855 13599 13861
rect 13541 13852 13553 13855
rect 13403 13824 13553 13852
rect 13403 13821 13415 13824
rect 13357 13815 13415 13821
rect 13541 13821 13553 13824
rect 13587 13821 13599 13855
rect 13541 13815 13599 13821
rect 13814 13812 13820 13864
rect 13872 13812 13878 13864
rect 13906 13812 13912 13864
rect 13964 13852 13970 13864
rect 14660 13861 14688 13892
rect 14001 13855 14059 13861
rect 14001 13852 14013 13855
rect 13964 13824 14013 13852
rect 13964 13812 13970 13824
rect 14001 13821 14013 13824
rect 14047 13821 14059 13855
rect 14001 13815 14059 13821
rect 14645 13855 14703 13861
rect 14645 13821 14657 13855
rect 14691 13821 14703 13855
rect 14645 13815 14703 13821
rect 14734 13812 14740 13864
rect 14792 13852 14798 13864
rect 15028 13861 15056 13892
rect 15212 13892 15393 13920
rect 14921 13855 14979 13861
rect 14921 13852 14933 13855
rect 14792 13824 14933 13852
rect 14792 13812 14798 13824
rect 14921 13821 14933 13824
rect 14967 13821 14979 13855
rect 14921 13815 14979 13821
rect 15013 13855 15071 13861
rect 15013 13821 15025 13855
rect 15059 13852 15071 13855
rect 15102 13852 15108 13864
rect 15059 13824 15108 13852
rect 15059 13821 15071 13824
rect 15013 13815 15071 13821
rect 15102 13812 15108 13824
rect 15160 13812 15166 13864
rect 15212 13861 15240 13892
rect 15381 13889 15393 13892
rect 15427 13889 15439 13923
rect 15381 13883 15439 13889
rect 16114 13880 16120 13932
rect 16172 13920 16178 13932
rect 16390 13920 16396 13932
rect 16172 13892 16396 13920
rect 16172 13880 16178 13892
rect 16390 13880 16396 13892
rect 16448 13880 16454 13932
rect 15197 13855 15255 13861
rect 15197 13821 15209 13855
rect 15243 13821 15255 13855
rect 15197 13815 15255 13821
rect 15286 13812 15292 13864
rect 15344 13812 15350 13864
rect 15470 13812 15476 13864
rect 15528 13812 15534 13864
rect 15930 13812 15936 13864
rect 15988 13852 15994 13864
rect 16025 13855 16083 13861
rect 16025 13852 16037 13855
rect 15988 13824 16037 13852
rect 15988 13812 15994 13824
rect 16025 13821 16037 13824
rect 16071 13852 16083 13855
rect 16071 13824 16160 13852
rect 16071 13821 16083 13824
rect 16025 13815 16083 13821
rect 12066 13784 12072 13796
rect 11624 13756 12072 13784
rect 12066 13744 12072 13756
rect 12124 13784 12130 13796
rect 12713 13787 12771 13793
rect 12713 13784 12725 13787
rect 12124 13756 12725 13784
rect 12124 13744 12130 13756
rect 12713 13753 12725 13756
rect 12759 13753 12771 13787
rect 14461 13787 14519 13793
rect 14461 13784 14473 13787
rect 12713 13747 12771 13753
rect 13004 13756 14473 13784
rect 1213 13719 1271 13725
rect 1213 13685 1225 13719
rect 1259 13716 1271 13719
rect 1302 13716 1308 13728
rect 1259 13688 1308 13716
rect 1259 13685 1271 13688
rect 1213 13679 1271 13685
rect 1302 13676 1308 13688
rect 1360 13676 1366 13728
rect 2590 13676 2596 13728
rect 2648 13716 2654 13728
rect 2685 13719 2743 13725
rect 2685 13716 2697 13719
rect 2648 13688 2697 13716
rect 2648 13676 2654 13688
rect 2685 13685 2697 13688
rect 2731 13685 2743 13719
rect 2685 13679 2743 13685
rect 3878 13676 3884 13728
rect 3936 13716 3942 13728
rect 4065 13719 4123 13725
rect 4065 13716 4077 13719
rect 3936 13688 4077 13716
rect 3936 13676 3942 13688
rect 4065 13685 4077 13688
rect 4111 13685 4123 13719
rect 4065 13679 4123 13685
rect 6825 13719 6883 13725
rect 6825 13685 6837 13719
rect 6871 13716 6883 13719
rect 7466 13716 7472 13728
rect 6871 13688 7472 13716
rect 6871 13685 6883 13688
rect 6825 13679 6883 13685
rect 7466 13676 7472 13688
rect 7524 13676 7530 13728
rect 7929 13719 7987 13725
rect 7929 13685 7941 13719
rect 7975 13716 7987 13719
rect 8294 13716 8300 13728
rect 7975 13688 8300 13716
rect 7975 13685 7987 13688
rect 7929 13679 7987 13685
rect 8294 13676 8300 13688
rect 8352 13676 8358 13728
rect 8573 13719 8631 13725
rect 8573 13685 8585 13719
rect 8619 13716 8631 13719
rect 8662 13716 8668 13728
rect 8619 13688 8668 13716
rect 8619 13685 8631 13688
rect 8573 13679 8631 13685
rect 8662 13676 8668 13688
rect 8720 13716 8726 13728
rect 9214 13716 9220 13728
rect 8720 13688 9220 13716
rect 8720 13676 8726 13688
rect 9214 13676 9220 13688
rect 9272 13716 9278 13728
rect 10042 13716 10048 13728
rect 9272 13688 10048 13716
rect 9272 13676 9278 13688
rect 10042 13676 10048 13688
rect 10100 13676 10106 13728
rect 10226 13676 10232 13728
rect 10284 13676 10290 13728
rect 10318 13676 10324 13728
rect 10376 13676 10382 13728
rect 10502 13676 10508 13728
rect 10560 13716 10566 13728
rect 11698 13716 11704 13728
rect 10560 13688 11704 13716
rect 10560 13676 10566 13688
rect 11698 13676 11704 13688
rect 11756 13676 11762 13728
rect 12250 13676 12256 13728
rect 12308 13716 12314 13728
rect 13004 13716 13032 13756
rect 14461 13753 14473 13756
rect 14507 13753 14519 13787
rect 16132 13784 16160 13824
rect 16206 13812 16212 13864
rect 16264 13852 16270 13864
rect 16485 13855 16543 13861
rect 16485 13852 16497 13855
rect 16264 13824 16497 13852
rect 16264 13812 16270 13824
rect 16485 13821 16497 13824
rect 16531 13821 16543 13855
rect 16485 13815 16543 13821
rect 16301 13787 16359 13793
rect 16301 13784 16313 13787
rect 16132 13756 16313 13784
rect 14461 13747 14519 13753
rect 16301 13753 16313 13756
rect 16347 13753 16359 13787
rect 16684 13784 16712 13960
rect 16761 13957 16773 13991
rect 16807 13988 16819 13991
rect 16942 13988 16948 14000
rect 16807 13960 16948 13988
rect 16807 13957 16819 13960
rect 16761 13951 16819 13957
rect 16942 13948 16948 13960
rect 17000 13948 17006 14000
rect 17126 13920 17132 13932
rect 16960 13892 17132 13920
rect 16761 13855 16819 13861
rect 16761 13821 16773 13855
rect 16807 13852 16819 13855
rect 16850 13852 16856 13864
rect 16807 13824 16856 13852
rect 16807 13821 16819 13824
rect 16761 13815 16819 13821
rect 16850 13812 16856 13824
rect 16908 13812 16914 13864
rect 16960 13861 16988 13892
rect 17126 13880 17132 13892
rect 17184 13880 17190 13932
rect 17236 13920 17264 14028
rect 19334 14016 19340 14068
rect 19392 14056 19398 14068
rect 21634 14056 21640 14068
rect 19392 14028 21640 14056
rect 19392 14016 19398 14028
rect 21634 14016 21640 14028
rect 21692 14016 21698 14068
rect 19610 13988 19616 14000
rect 17880 13960 19616 13988
rect 17313 13923 17371 13929
rect 17313 13920 17325 13923
rect 17236 13892 17325 13920
rect 17313 13889 17325 13892
rect 17359 13920 17371 13923
rect 17770 13920 17776 13932
rect 17359 13892 17776 13920
rect 17359 13889 17371 13892
rect 17313 13883 17371 13889
rect 17770 13880 17776 13892
rect 17828 13880 17834 13932
rect 16945 13855 17003 13861
rect 16945 13821 16957 13855
rect 16991 13821 17003 13855
rect 16945 13815 17003 13821
rect 17037 13855 17095 13861
rect 17037 13821 17049 13855
rect 17083 13852 17095 13855
rect 17880 13852 17908 13960
rect 19610 13948 19616 13960
rect 19668 13948 19674 14000
rect 20346 13988 20352 14000
rect 20088 13960 20352 13988
rect 19153 13923 19211 13929
rect 19153 13889 19165 13923
rect 19199 13920 19211 13923
rect 19429 13923 19487 13929
rect 19429 13920 19441 13923
rect 19199 13892 19441 13920
rect 19199 13889 19211 13892
rect 19153 13883 19211 13889
rect 19429 13889 19441 13892
rect 19475 13889 19487 13923
rect 19702 13920 19708 13932
rect 19429 13883 19487 13889
rect 19628 13892 19708 13920
rect 17083 13824 17908 13852
rect 17083 13821 17095 13824
rect 17037 13815 17095 13821
rect 17052 13784 17080 13815
rect 18230 13812 18236 13864
rect 18288 13852 18294 13864
rect 18288 13824 18736 13852
rect 18288 13812 18294 13824
rect 16684 13756 17080 13784
rect 16301 13747 16359 13753
rect 18414 13744 18420 13796
rect 18472 13744 18478 13796
rect 18708 13784 18736 13824
rect 18782 13812 18788 13864
rect 18840 13852 18846 13864
rect 19061 13855 19119 13861
rect 19061 13852 19073 13855
rect 18840 13824 19073 13852
rect 18840 13812 18846 13824
rect 19061 13821 19073 13824
rect 19107 13821 19119 13855
rect 19061 13815 19119 13821
rect 19334 13812 19340 13864
rect 19392 13812 19398 13864
rect 19628 13861 19656 13892
rect 19702 13880 19708 13892
rect 19760 13920 19766 13932
rect 19978 13920 19984 13932
rect 19760 13892 19984 13920
rect 19760 13880 19766 13892
rect 19978 13880 19984 13892
rect 20036 13880 20042 13932
rect 19521 13855 19579 13861
rect 19521 13852 19533 13855
rect 19444 13824 19533 13852
rect 19444 13784 19472 13824
rect 19521 13821 19533 13824
rect 19567 13821 19579 13855
rect 19521 13815 19579 13821
rect 19613 13855 19671 13861
rect 19613 13821 19625 13855
rect 19659 13821 19671 13855
rect 19613 13815 19671 13821
rect 19797 13855 19855 13861
rect 19797 13821 19809 13855
rect 19843 13821 19855 13855
rect 19797 13815 19855 13821
rect 19889 13855 19947 13861
rect 19889 13821 19901 13855
rect 19935 13852 19947 13855
rect 20088 13852 20116 13960
rect 20346 13948 20352 13960
rect 20404 13948 20410 14000
rect 20717 13991 20775 13997
rect 20717 13988 20729 13991
rect 20456 13960 20729 13988
rect 20254 13880 20260 13932
rect 20312 13920 20318 13932
rect 20456 13920 20484 13960
rect 20717 13957 20729 13960
rect 20763 13957 20775 13991
rect 20717 13951 20775 13957
rect 20806 13948 20812 14000
rect 20864 13988 20870 14000
rect 22097 13991 22155 13997
rect 22097 13988 22109 13991
rect 20864 13960 22109 13988
rect 20864 13948 20870 13960
rect 22097 13957 22109 13960
rect 22143 13957 22155 13991
rect 22097 13951 22155 13957
rect 21545 13923 21603 13929
rect 21545 13920 21557 13923
rect 20312 13892 20484 13920
rect 21192 13892 21557 13920
rect 20312 13880 20318 13892
rect 20349 13855 20407 13861
rect 20349 13852 20361 13855
rect 19935 13824 20116 13852
rect 20180 13824 20361 13852
rect 19935 13821 19947 13824
rect 19889 13815 19947 13821
rect 18708 13756 19472 13784
rect 19812 13784 19840 13815
rect 20180 13784 20208 13824
rect 20349 13821 20361 13824
rect 20395 13852 20407 13855
rect 20530 13852 20536 13864
rect 20395 13824 20536 13852
rect 20395 13821 20407 13824
rect 20349 13815 20407 13821
rect 20530 13812 20536 13824
rect 20588 13852 20594 13864
rect 21085 13855 21143 13861
rect 21085 13852 21097 13855
rect 20588 13824 21097 13852
rect 20588 13812 20594 13824
rect 21085 13821 21097 13824
rect 21131 13821 21143 13855
rect 21085 13815 21143 13821
rect 21192 13784 21220 13892
rect 21545 13889 21557 13892
rect 21591 13889 21603 13923
rect 21545 13883 21603 13889
rect 22005 13923 22063 13929
rect 22005 13889 22017 13923
rect 22051 13920 22063 13923
rect 22373 13923 22431 13929
rect 22373 13920 22385 13923
rect 22051 13892 22385 13920
rect 22051 13889 22063 13892
rect 22005 13883 22063 13889
rect 22373 13889 22385 13892
rect 22419 13889 22431 13923
rect 22373 13883 22431 13889
rect 21634 13812 21640 13864
rect 21692 13812 21698 13864
rect 22462 13812 22468 13864
rect 22520 13812 22526 13864
rect 19812 13756 20208 13784
rect 20548 13756 21220 13784
rect 20548 13728 20576 13756
rect 12308 13688 13032 13716
rect 13173 13719 13231 13725
rect 12308 13676 12314 13688
rect 13173 13685 13185 13719
rect 13219 13716 13231 13719
rect 14550 13716 14556 13728
rect 13219 13688 14556 13716
rect 13219 13685 13231 13688
rect 13173 13679 13231 13685
rect 14550 13676 14556 13688
rect 14608 13676 14614 13728
rect 14829 13719 14887 13725
rect 14829 13685 14841 13719
rect 14875 13716 14887 13719
rect 15102 13716 15108 13728
rect 14875 13688 15108 13716
rect 14875 13685 14887 13688
rect 14829 13679 14887 13685
rect 15102 13676 15108 13688
rect 15160 13676 15166 13728
rect 16206 13676 16212 13728
rect 16264 13676 16270 13728
rect 16390 13676 16396 13728
rect 16448 13716 16454 13728
rect 16669 13719 16727 13725
rect 16669 13716 16681 13719
rect 16448 13688 16681 13716
rect 16448 13676 16454 13688
rect 16669 13685 16681 13688
rect 16715 13685 16727 13719
rect 16669 13679 16727 13685
rect 16758 13676 16764 13728
rect 16816 13716 16822 13728
rect 17543 13719 17601 13725
rect 17543 13716 17555 13719
rect 16816 13688 17555 13716
rect 16816 13676 16822 13688
rect 17543 13685 17555 13688
rect 17589 13716 17601 13719
rect 17678 13716 17684 13728
rect 17589 13688 17684 13716
rect 17589 13685 17601 13688
rect 17543 13679 17601 13685
rect 17678 13676 17684 13688
rect 17736 13676 17742 13728
rect 18690 13676 18696 13728
rect 18748 13676 18754 13728
rect 19794 13676 19800 13728
rect 19852 13716 19858 13728
rect 19889 13719 19947 13725
rect 19889 13716 19901 13719
rect 19852 13688 19901 13716
rect 19852 13676 19858 13688
rect 19889 13685 19901 13688
rect 19935 13685 19947 13719
rect 19889 13679 19947 13685
rect 19978 13676 19984 13728
rect 20036 13676 20042 13728
rect 20530 13676 20536 13728
rect 20588 13676 20594 13728
rect 20625 13719 20683 13725
rect 20625 13685 20637 13719
rect 20671 13716 20683 13719
rect 21174 13716 21180 13728
rect 20671 13688 21180 13716
rect 20671 13685 20683 13688
rect 20625 13679 20683 13685
rect 21174 13676 21180 13688
rect 21232 13676 21238 13728
rect 552 13626 23368 13648
rect 552 13574 4366 13626
rect 4418 13574 4430 13626
rect 4482 13574 4494 13626
rect 4546 13574 4558 13626
rect 4610 13574 4622 13626
rect 4674 13574 4686 13626
rect 4738 13574 10366 13626
rect 10418 13574 10430 13626
rect 10482 13574 10494 13626
rect 10546 13574 10558 13626
rect 10610 13574 10622 13626
rect 10674 13574 10686 13626
rect 10738 13574 16366 13626
rect 16418 13574 16430 13626
rect 16482 13574 16494 13626
rect 16546 13574 16558 13626
rect 16610 13574 16622 13626
rect 16674 13574 16686 13626
rect 16738 13574 22366 13626
rect 22418 13574 22430 13626
rect 22482 13574 22494 13626
rect 22546 13574 22558 13626
rect 22610 13574 22622 13626
rect 22674 13574 22686 13626
rect 22738 13574 23368 13626
rect 552 13552 23368 13574
rect 1302 13472 1308 13524
rect 1360 13512 1366 13524
rect 1857 13515 1915 13521
rect 1857 13512 1869 13515
rect 1360 13484 1869 13512
rect 1360 13472 1366 13484
rect 1857 13481 1869 13484
rect 1903 13481 1915 13515
rect 1857 13475 1915 13481
rect 2038 13472 2044 13524
rect 2096 13472 2102 13524
rect 2590 13472 2596 13524
rect 2648 13512 2654 13524
rect 2648 13484 3188 13512
rect 2648 13472 2654 13484
rect 1118 13404 1124 13456
rect 1176 13444 1182 13456
rect 1213 13447 1271 13453
rect 1213 13444 1225 13447
rect 1176 13416 1225 13444
rect 1176 13404 1182 13416
rect 1213 13413 1225 13416
rect 1259 13413 1271 13447
rect 1213 13407 1271 13413
rect 2869 13447 2927 13453
rect 2869 13413 2881 13447
rect 2915 13444 2927 13447
rect 3050 13444 3056 13456
rect 2915 13416 3056 13444
rect 2915 13413 2927 13416
rect 2869 13407 2927 13413
rect 3050 13404 3056 13416
rect 3108 13404 3114 13456
rect 842 13336 848 13388
rect 900 13336 906 13388
rect 1489 13379 1547 13385
rect 1489 13345 1501 13379
rect 1535 13376 1547 13379
rect 1762 13376 1768 13388
rect 1535 13348 1768 13376
rect 1535 13345 1547 13348
rect 1489 13339 1547 13345
rect 1762 13336 1768 13348
rect 1820 13336 1826 13388
rect 2406 13336 2412 13388
rect 2464 13376 2470 13388
rect 3160 13385 3188 13484
rect 6178 13472 6184 13524
rect 6236 13512 6242 13524
rect 6273 13515 6331 13521
rect 6273 13512 6285 13515
rect 6236 13484 6285 13512
rect 6236 13472 6242 13484
rect 6273 13481 6285 13484
rect 6319 13512 6331 13515
rect 7558 13512 7564 13524
rect 6319 13484 7564 13512
rect 6319 13481 6331 13484
rect 6273 13475 6331 13481
rect 7558 13472 7564 13484
rect 7616 13472 7622 13524
rect 7834 13472 7840 13524
rect 7892 13512 7898 13524
rect 8018 13512 8024 13524
rect 7892 13484 8024 13512
rect 7892 13472 7898 13484
rect 8018 13472 8024 13484
rect 8076 13472 8082 13524
rect 8662 13472 8668 13524
rect 8720 13472 8726 13524
rect 9674 13472 9680 13524
rect 9732 13512 9738 13524
rect 9861 13515 9919 13521
rect 9861 13512 9873 13515
rect 9732 13484 9873 13512
rect 9732 13472 9738 13484
rect 9861 13481 9873 13484
rect 9907 13481 9919 13515
rect 9861 13475 9919 13481
rect 10226 13472 10232 13524
rect 10284 13512 10290 13524
rect 10597 13515 10655 13521
rect 10597 13512 10609 13515
rect 10284 13484 10609 13512
rect 10284 13472 10290 13484
rect 10597 13481 10609 13484
rect 10643 13481 10655 13515
rect 10597 13475 10655 13481
rect 10965 13515 11023 13521
rect 10965 13481 10977 13515
rect 11011 13481 11023 13515
rect 10965 13475 11023 13481
rect 4614 13404 4620 13456
rect 4672 13444 4678 13456
rect 5350 13444 5356 13456
rect 4672 13416 5356 13444
rect 4672 13404 4678 13416
rect 5350 13404 5356 13416
rect 5408 13404 5414 13456
rect 5534 13404 5540 13456
rect 5592 13444 5598 13456
rect 6549 13447 6607 13453
rect 6549 13444 6561 13447
rect 5592 13416 6561 13444
rect 5592 13404 5598 13416
rect 6549 13413 6561 13416
rect 6595 13413 6607 13447
rect 6549 13407 6607 13413
rect 6914 13404 6920 13456
rect 6972 13444 6978 13456
rect 7009 13447 7067 13453
rect 7009 13444 7021 13447
rect 6972 13416 7021 13444
rect 6972 13404 6978 13416
rect 7009 13413 7021 13416
rect 7055 13413 7067 13447
rect 7009 13407 7067 13413
rect 7098 13404 7104 13456
rect 7156 13444 7162 13456
rect 7377 13447 7435 13453
rect 7377 13444 7389 13447
rect 7156 13416 7389 13444
rect 7156 13404 7162 13416
rect 7377 13413 7389 13416
rect 7423 13444 7435 13447
rect 7466 13444 7472 13456
rect 7423 13416 7472 13444
rect 7423 13413 7435 13416
rect 7377 13407 7435 13413
rect 7466 13404 7472 13416
rect 7524 13444 7530 13456
rect 9306 13444 9312 13456
rect 7524 13416 9312 13444
rect 7524 13404 7530 13416
rect 9306 13404 9312 13416
rect 9364 13404 9370 13456
rect 10134 13444 10140 13456
rect 9600 13416 10140 13444
rect 2593 13379 2651 13385
rect 2593 13376 2605 13379
rect 2464 13348 2605 13376
rect 2464 13336 2470 13348
rect 2593 13345 2605 13348
rect 2639 13345 2651 13379
rect 2593 13339 2651 13345
rect 3145 13379 3203 13385
rect 3145 13345 3157 13379
rect 3191 13345 3203 13379
rect 3145 13339 3203 13345
rect 2225 13311 2283 13317
rect 2225 13277 2237 13311
rect 2271 13308 2283 13311
rect 2498 13308 2504 13320
rect 2271 13280 2504 13308
rect 2271 13277 2283 13280
rect 2225 13271 2283 13277
rect 2498 13268 2504 13280
rect 2556 13268 2562 13320
rect 2608 13240 2636 13339
rect 3602 13336 3608 13388
rect 3660 13336 3666 13388
rect 4246 13336 4252 13388
rect 4304 13336 4310 13388
rect 4982 13336 4988 13388
rect 5040 13376 5046 13388
rect 5813 13379 5871 13385
rect 5813 13376 5825 13379
rect 5040 13348 5825 13376
rect 5040 13336 5046 13348
rect 5813 13345 5825 13348
rect 5859 13345 5871 13379
rect 5813 13339 5871 13345
rect 6641 13379 6699 13385
rect 6641 13345 6653 13379
rect 6687 13376 6699 13379
rect 6687 13348 8156 13376
rect 6687 13345 6699 13348
rect 6641 13339 6699 13345
rect 2682 13268 2688 13320
rect 2740 13268 2746 13320
rect 3697 13311 3755 13317
rect 3697 13277 3709 13311
rect 3743 13308 3755 13311
rect 3973 13311 4031 13317
rect 3743 13280 3924 13308
rect 3743 13277 3755 13280
rect 3697 13271 3755 13277
rect 2961 13243 3019 13249
rect 2961 13240 2973 13243
rect 1228 13212 1900 13240
rect 2608 13212 2973 13240
rect 1228 13181 1256 13212
rect 1213 13175 1271 13181
rect 1213 13141 1225 13175
rect 1259 13141 1271 13175
rect 1213 13135 1271 13141
rect 1397 13175 1455 13181
rect 1397 13141 1409 13175
rect 1443 13172 1455 13175
rect 1762 13172 1768 13184
rect 1443 13144 1768 13172
rect 1443 13141 1455 13144
rect 1397 13135 1455 13141
rect 1762 13132 1768 13144
rect 1820 13132 1826 13184
rect 1872 13181 1900 13212
rect 2961 13209 2973 13212
rect 3007 13209 3019 13243
rect 2961 13203 3019 13209
rect 1857 13175 1915 13181
rect 1857 13141 1869 13175
rect 1903 13172 1915 13175
rect 2130 13172 2136 13184
rect 1903 13144 2136 13172
rect 1903 13141 1915 13144
rect 1857 13135 1915 13141
rect 2130 13132 2136 13144
rect 2188 13132 2194 13184
rect 3896 13172 3924 13280
rect 3973 13277 3985 13311
rect 4019 13308 4031 13311
rect 4154 13308 4160 13320
rect 4019 13280 4160 13308
rect 4019 13277 4031 13280
rect 3973 13271 4031 13277
rect 4154 13268 4160 13280
rect 4212 13268 4218 13320
rect 7650 13308 7656 13320
rect 7314 13280 7656 13308
rect 7650 13268 7656 13280
rect 7708 13268 7714 13320
rect 8128 13308 8156 13348
rect 8294 13336 8300 13388
rect 8352 13376 8358 13388
rect 8481 13379 8539 13385
rect 8481 13376 8493 13379
rect 8352 13348 8493 13376
rect 8352 13336 8358 13348
rect 8481 13345 8493 13348
rect 8527 13345 8539 13379
rect 8481 13339 8539 13345
rect 9214 13336 9220 13388
rect 9272 13336 9278 13388
rect 9401 13379 9459 13385
rect 9401 13345 9413 13379
rect 9447 13345 9459 13379
rect 9401 13339 9459 13345
rect 9030 13308 9036 13320
rect 8128 13280 9036 13308
rect 9030 13268 9036 13280
rect 9088 13268 9094 13320
rect 9416 13308 9444 13339
rect 9490 13336 9496 13388
rect 9548 13336 9554 13388
rect 9600 13385 9628 13416
rect 10134 13404 10140 13416
rect 10192 13404 10198 13456
rect 9585 13379 9643 13385
rect 9585 13345 9597 13379
rect 9631 13345 9643 13379
rect 9585 13339 9643 13345
rect 9674 13336 9680 13388
rect 9732 13376 9738 13388
rect 10244 13385 10272 13472
rect 10980 13444 11008 13475
rect 11330 13472 11336 13524
rect 11388 13512 11394 13524
rect 11388 13484 16344 13512
rect 11388 13472 11394 13484
rect 10704 13416 11008 13444
rect 10229 13379 10287 13385
rect 9732 13348 10196 13376
rect 9732 13336 9738 13348
rect 10168 13308 10196 13348
rect 10229 13345 10241 13379
rect 10275 13345 10287 13379
rect 10229 13339 10287 13345
rect 10502 13336 10508 13388
rect 10560 13336 10566 13388
rect 10704 13308 10732 13416
rect 11698 13404 11704 13456
rect 11756 13404 11762 13456
rect 11790 13404 11796 13456
rect 11848 13404 11854 13456
rect 11977 13447 12035 13453
rect 11977 13413 11989 13447
rect 12023 13444 12035 13447
rect 12342 13444 12348 13456
rect 12023 13416 12348 13444
rect 12023 13413 12035 13416
rect 11977 13407 12035 13413
rect 12342 13404 12348 13416
rect 12400 13404 12406 13456
rect 12544 13416 13952 13444
rect 10781 13379 10839 13385
rect 10781 13345 10793 13379
rect 10827 13376 10839 13379
rect 11054 13376 11060 13388
rect 10827 13348 11060 13376
rect 10827 13345 10839 13348
rect 10781 13339 10839 13345
rect 11054 13336 11060 13348
rect 11112 13336 11118 13388
rect 11238 13336 11244 13388
rect 11296 13336 11302 13388
rect 11333 13379 11391 13385
rect 11333 13345 11345 13379
rect 11379 13376 11391 13379
rect 11609 13379 11667 13385
rect 11609 13376 11621 13379
rect 11379 13348 11621 13376
rect 11379 13345 11391 13348
rect 11333 13339 11391 13345
rect 11609 13345 11621 13348
rect 11655 13345 11667 13379
rect 11609 13339 11667 13345
rect 9416 13280 9996 13308
rect 10168 13280 10732 13308
rect 4617 13243 4675 13249
rect 4617 13209 4629 13243
rect 4663 13240 4675 13243
rect 5350 13240 5356 13252
rect 4663 13212 5356 13240
rect 4663 13209 4675 13212
rect 4617 13203 4675 13209
rect 5350 13200 5356 13212
rect 5408 13200 5414 13252
rect 5997 13243 6055 13249
rect 5997 13209 6009 13243
rect 6043 13240 6055 13243
rect 6178 13240 6184 13252
rect 6043 13212 6184 13240
rect 6043 13209 6055 13212
rect 5997 13203 6055 13209
rect 6178 13200 6184 13212
rect 6236 13200 6242 13252
rect 7561 13243 7619 13249
rect 7561 13209 7573 13243
rect 7607 13240 7619 13243
rect 9766 13240 9772 13252
rect 7607 13212 9772 13240
rect 7607 13209 7619 13212
rect 7561 13203 7619 13209
rect 9766 13200 9772 13212
rect 9824 13200 9830 13252
rect 9968 13249 9996 13280
rect 10962 13268 10968 13320
rect 11020 13308 11026 13320
rect 11149 13311 11207 13317
rect 11149 13308 11161 13311
rect 11020 13280 11161 13308
rect 11020 13268 11026 13280
rect 11149 13277 11161 13280
rect 11195 13277 11207 13311
rect 11149 13271 11207 13277
rect 11425 13311 11483 13317
rect 11425 13277 11437 13311
rect 11471 13308 11483 13311
rect 11716 13308 11744 13404
rect 12250 13336 12256 13388
rect 12308 13376 12314 13388
rect 12544 13385 12572 13416
rect 12437 13379 12495 13385
rect 12437 13376 12449 13379
rect 12308 13348 12449 13376
rect 12308 13336 12314 13348
rect 12437 13345 12449 13348
rect 12483 13345 12495 13379
rect 12437 13339 12495 13345
rect 12529 13379 12587 13385
rect 12529 13345 12541 13379
rect 12575 13345 12587 13379
rect 12529 13339 12587 13345
rect 12544 13308 12572 13339
rect 12710 13336 12716 13388
rect 12768 13376 12774 13388
rect 13924 13385 13952 13416
rect 14090 13404 14096 13456
rect 14148 13444 14154 13456
rect 15286 13444 15292 13456
rect 14148 13416 15292 13444
rect 14148 13404 14154 13416
rect 15286 13404 15292 13416
rect 15344 13404 15350 13456
rect 13081 13379 13139 13385
rect 13081 13376 13093 13379
rect 12768 13348 13093 13376
rect 12768 13336 12774 13348
rect 13081 13345 13093 13348
rect 13127 13345 13139 13379
rect 13081 13339 13139 13345
rect 13909 13379 13967 13385
rect 13909 13345 13921 13379
rect 13955 13345 13967 13379
rect 13909 13339 13967 13345
rect 15102 13336 15108 13388
rect 15160 13336 15166 13388
rect 16316 13385 16344 13484
rect 16574 13472 16580 13524
rect 16632 13512 16638 13524
rect 16669 13515 16727 13521
rect 16669 13512 16681 13515
rect 16632 13484 16681 13512
rect 16632 13472 16638 13484
rect 16669 13481 16681 13484
rect 16715 13481 16727 13515
rect 17034 13512 17040 13524
rect 16669 13475 16727 13481
rect 16868 13484 17040 13512
rect 16301 13379 16359 13385
rect 16301 13345 16313 13379
rect 16347 13345 16359 13379
rect 16301 13339 16359 13345
rect 16761 13379 16819 13385
rect 16761 13345 16773 13379
rect 16807 13376 16819 13379
rect 16868 13376 16896 13484
rect 17034 13472 17040 13484
rect 17092 13472 17098 13524
rect 19429 13515 19487 13521
rect 19429 13481 19441 13515
rect 19475 13512 19487 13515
rect 19702 13512 19708 13524
rect 19475 13484 19708 13512
rect 19475 13481 19487 13484
rect 19429 13475 19487 13481
rect 19702 13472 19708 13484
rect 19760 13472 19766 13524
rect 16960 13416 17540 13444
rect 16960 13385 16988 13416
rect 17512 13388 17540 13416
rect 18598 13404 18604 13456
rect 18656 13444 18662 13456
rect 19886 13444 19892 13456
rect 18656 13416 19892 13444
rect 18656 13404 18662 13416
rect 19886 13404 19892 13416
rect 19944 13404 19950 13456
rect 16807 13348 16896 13376
rect 16945 13379 17003 13385
rect 16807 13345 16819 13348
rect 16761 13339 16819 13345
rect 16945 13345 16957 13379
rect 16991 13345 17003 13379
rect 16945 13339 17003 13345
rect 17034 13336 17040 13388
rect 17092 13376 17098 13388
rect 17221 13379 17279 13385
rect 17221 13376 17233 13379
rect 17092 13348 17233 13376
rect 17092 13336 17098 13348
rect 17221 13345 17233 13348
rect 17267 13345 17279 13379
rect 17221 13339 17279 13345
rect 17494 13336 17500 13388
rect 17552 13336 17558 13388
rect 17678 13336 17684 13388
rect 17736 13336 17742 13388
rect 17770 13336 17776 13388
rect 17828 13376 17834 13388
rect 17957 13379 18015 13385
rect 17957 13376 17969 13379
rect 17828 13348 17969 13376
rect 17828 13336 17834 13348
rect 17957 13345 17969 13348
rect 18003 13345 18015 13379
rect 17957 13339 18015 13345
rect 19610 13336 19616 13388
rect 19668 13376 19674 13388
rect 20530 13376 20536 13388
rect 19668 13348 20536 13376
rect 19668 13336 19674 13348
rect 20530 13336 20536 13348
rect 20588 13336 20594 13388
rect 11471 13280 11744 13308
rect 12268 13280 12572 13308
rect 11471 13277 11483 13280
rect 11425 13271 11483 13277
rect 12268 13252 12296 13280
rect 12802 13268 12808 13320
rect 12860 13268 12866 13320
rect 13354 13268 13360 13320
rect 13412 13308 13418 13320
rect 13817 13311 13875 13317
rect 13817 13308 13829 13311
rect 13412 13280 13829 13308
rect 13412 13268 13418 13280
rect 13817 13277 13829 13280
rect 13863 13277 13875 13311
rect 13817 13271 13875 13277
rect 14734 13268 14740 13320
rect 14792 13308 14798 13320
rect 15013 13311 15071 13317
rect 15013 13308 15025 13311
rect 14792 13280 15025 13308
rect 14792 13268 14798 13280
rect 15013 13277 15025 13280
rect 15059 13277 15071 13311
rect 15013 13271 15071 13277
rect 15194 13268 15200 13320
rect 15252 13308 15258 13320
rect 16209 13311 16267 13317
rect 16209 13308 16221 13311
rect 15252 13280 16221 13308
rect 15252 13268 15258 13280
rect 16209 13277 16221 13280
rect 16255 13308 16267 13311
rect 16666 13308 16672 13320
rect 16255 13280 16672 13308
rect 16255 13277 16267 13280
rect 16209 13271 16267 13277
rect 16666 13268 16672 13280
rect 16724 13268 16730 13320
rect 16853 13311 16911 13317
rect 16853 13277 16865 13311
rect 16899 13308 16911 13311
rect 17865 13311 17923 13317
rect 17865 13308 17877 13311
rect 16899 13280 17877 13308
rect 16899 13277 16911 13280
rect 16853 13271 16911 13277
rect 17865 13277 17877 13280
rect 17911 13277 17923 13311
rect 18598 13308 18604 13320
rect 17865 13271 17923 13277
rect 18340 13280 18604 13308
rect 9953 13243 10011 13249
rect 9953 13209 9965 13243
rect 9999 13209 10011 13243
rect 9953 13203 10011 13209
rect 12250 13200 12256 13252
rect 12308 13200 12314 13252
rect 13722 13240 13728 13252
rect 12636 13212 13728 13240
rect 3970 13172 3976 13184
rect 3896 13144 3976 13172
rect 3970 13132 3976 13144
rect 4028 13172 4034 13184
rect 5442 13172 5448 13184
rect 4028 13144 5448 13172
rect 4028 13132 4034 13144
rect 5442 13132 5448 13144
rect 5500 13132 5506 13184
rect 10134 13132 10140 13184
rect 10192 13132 10198 13184
rect 11606 13132 11612 13184
rect 11664 13172 11670 13184
rect 12636 13172 12664 13212
rect 13722 13200 13728 13212
rect 13780 13200 13786 13252
rect 15102 13200 15108 13252
rect 15160 13240 15166 13252
rect 18340 13240 18368 13280
rect 18598 13268 18604 13280
rect 18656 13268 18662 13320
rect 15160 13212 18368 13240
rect 15160 13200 15166 13212
rect 18414 13200 18420 13252
rect 18472 13240 18478 13252
rect 20806 13240 20812 13252
rect 18472 13212 20812 13240
rect 18472 13200 18478 13212
rect 20806 13200 20812 13212
rect 20864 13200 20870 13252
rect 11664 13144 12664 13172
rect 12713 13175 12771 13181
rect 11664 13132 11670 13144
rect 12713 13141 12725 13175
rect 12759 13172 12771 13175
rect 12986 13172 12992 13184
rect 12759 13144 12992 13172
rect 12759 13141 12771 13144
rect 12713 13135 12771 13141
rect 12986 13132 12992 13144
rect 13044 13132 13050 13184
rect 14182 13132 14188 13184
rect 14240 13132 14246 13184
rect 14829 13175 14887 13181
rect 14829 13141 14841 13175
rect 14875 13172 14887 13175
rect 14918 13172 14924 13184
rect 14875 13144 14924 13172
rect 14875 13141 14887 13144
rect 14829 13135 14887 13141
rect 14918 13132 14924 13144
rect 14976 13132 14982 13184
rect 15194 13132 15200 13184
rect 15252 13172 15258 13184
rect 17037 13175 17095 13181
rect 17037 13172 17049 13175
rect 15252 13144 17049 13172
rect 15252 13132 15258 13144
rect 17037 13141 17049 13144
rect 17083 13141 17095 13175
rect 17037 13135 17095 13141
rect 17126 13132 17132 13184
rect 17184 13172 17190 13184
rect 17586 13172 17592 13184
rect 17184 13144 17592 13172
rect 17184 13132 17190 13144
rect 17586 13132 17592 13144
rect 17644 13132 17650 13184
rect 18233 13175 18291 13181
rect 18233 13141 18245 13175
rect 18279 13172 18291 13175
rect 18874 13172 18880 13184
rect 18279 13144 18880 13172
rect 18279 13141 18291 13144
rect 18233 13135 18291 13141
rect 18874 13132 18880 13144
rect 18932 13132 18938 13184
rect 20070 13132 20076 13184
rect 20128 13172 20134 13184
rect 20254 13172 20260 13184
rect 20128 13144 20260 13172
rect 20128 13132 20134 13144
rect 20254 13132 20260 13144
rect 20312 13132 20318 13184
rect 20714 13132 20720 13184
rect 20772 13172 20778 13184
rect 21082 13172 21088 13184
rect 20772 13144 21088 13172
rect 20772 13132 20778 13144
rect 21082 13132 21088 13144
rect 21140 13132 21146 13184
rect 552 13082 23368 13104
rect 552 13030 1366 13082
rect 1418 13030 1430 13082
rect 1482 13030 1494 13082
rect 1546 13030 1558 13082
rect 1610 13030 1622 13082
rect 1674 13030 1686 13082
rect 1738 13030 7366 13082
rect 7418 13030 7430 13082
rect 7482 13030 7494 13082
rect 7546 13030 7558 13082
rect 7610 13030 7622 13082
rect 7674 13030 7686 13082
rect 7738 13030 13366 13082
rect 13418 13030 13430 13082
rect 13482 13030 13494 13082
rect 13546 13030 13558 13082
rect 13610 13030 13622 13082
rect 13674 13030 13686 13082
rect 13738 13030 19366 13082
rect 19418 13030 19430 13082
rect 19482 13030 19494 13082
rect 19546 13030 19558 13082
rect 19610 13030 19622 13082
rect 19674 13030 19686 13082
rect 19738 13030 23368 13082
rect 552 13008 23368 13030
rect 842 12928 848 12980
rect 900 12968 906 12980
rect 937 12971 995 12977
rect 937 12968 949 12971
rect 900 12940 949 12968
rect 900 12928 906 12940
rect 937 12937 949 12940
rect 983 12937 995 12971
rect 937 12931 995 12937
rect 1121 12971 1179 12977
rect 1121 12937 1133 12971
rect 1167 12937 1179 12971
rect 5074 12968 5080 12980
rect 1121 12931 1179 12937
rect 2746 12940 5080 12968
rect 750 12860 756 12912
rect 808 12900 814 12912
rect 1136 12900 1164 12931
rect 808 12872 1164 12900
rect 808 12860 814 12872
rect 1670 12860 1676 12912
rect 1728 12900 1734 12912
rect 2314 12900 2320 12912
rect 1728 12872 2320 12900
rect 1728 12860 1734 12872
rect 2314 12860 2320 12872
rect 2372 12860 2378 12912
rect 658 12792 664 12844
rect 716 12832 722 12844
rect 2746 12832 2774 12940
rect 5074 12928 5080 12940
rect 5132 12928 5138 12980
rect 6733 12971 6791 12977
rect 6733 12937 6745 12971
rect 6779 12968 6791 12971
rect 7190 12968 7196 12980
rect 6779 12940 7196 12968
rect 6779 12937 6791 12940
rect 6733 12931 6791 12937
rect 7190 12928 7196 12940
rect 7248 12928 7254 12980
rect 8754 12968 8760 12980
rect 7392 12940 8760 12968
rect 6270 12860 6276 12912
rect 6328 12900 6334 12912
rect 7392 12900 7420 12940
rect 8754 12928 8760 12940
rect 8812 12928 8818 12980
rect 9214 12928 9220 12980
rect 9272 12968 9278 12980
rect 9493 12971 9551 12977
rect 9493 12968 9505 12971
rect 9272 12940 9505 12968
rect 9272 12928 9278 12940
rect 9493 12937 9505 12940
rect 9539 12937 9551 12971
rect 9493 12931 9551 12937
rect 10962 12928 10968 12980
rect 11020 12928 11026 12980
rect 11885 12971 11943 12977
rect 11885 12968 11897 12971
rect 11072 12940 11897 12968
rect 6328 12872 7420 12900
rect 7469 12903 7527 12909
rect 6328 12860 6334 12872
rect 7469 12869 7481 12903
rect 7515 12900 7527 12903
rect 7834 12900 7840 12912
rect 7515 12872 7840 12900
rect 7515 12869 7527 12872
rect 7469 12863 7527 12869
rect 7834 12860 7840 12872
rect 7892 12860 7898 12912
rect 9953 12903 10011 12909
rect 9953 12869 9965 12903
rect 9999 12900 10011 12903
rect 10042 12900 10048 12912
rect 9999 12872 10048 12900
rect 9999 12869 10011 12872
rect 9953 12863 10011 12869
rect 10042 12860 10048 12872
rect 10100 12860 10106 12912
rect 10502 12860 10508 12912
rect 10560 12900 10566 12912
rect 11072 12900 11100 12940
rect 11885 12937 11897 12940
rect 11931 12937 11943 12971
rect 11885 12931 11943 12937
rect 11609 12903 11667 12909
rect 11609 12900 11621 12903
rect 10560 12872 11100 12900
rect 11164 12872 11621 12900
rect 10560 12860 10566 12872
rect 6822 12832 6828 12844
rect 716 12804 2774 12832
rect 6118 12804 6828 12832
rect 716 12792 722 12804
rect 6822 12792 6828 12804
rect 6880 12792 6886 12844
rect 6914 12792 6920 12844
rect 6972 12832 6978 12844
rect 7009 12835 7067 12841
rect 7009 12832 7021 12835
rect 6972 12804 7021 12832
rect 6972 12792 6978 12804
rect 7009 12801 7021 12804
rect 7055 12832 7067 12835
rect 11164 12832 11192 12872
rect 11609 12869 11621 12872
rect 11655 12869 11667 12903
rect 11900 12900 11928 12931
rect 11974 12928 11980 12980
rect 12032 12968 12038 12980
rect 14645 12971 14703 12977
rect 14645 12968 14657 12971
rect 12032 12940 14657 12968
rect 12032 12928 12038 12940
rect 14645 12937 14657 12940
rect 14691 12937 14703 12971
rect 19429 12971 19487 12977
rect 19429 12968 19441 12971
rect 14645 12931 14703 12937
rect 15396 12940 19441 12968
rect 11900 12872 12572 12900
rect 11609 12863 11667 12869
rect 11330 12832 11336 12844
rect 7055 12804 7512 12832
rect 7055 12801 7067 12804
rect 7009 12795 7067 12801
rect 7484 12776 7512 12804
rect 10060 12804 11192 12832
rect 1026 12724 1032 12776
rect 1084 12739 1090 12776
rect 1084 12733 1133 12739
rect 1084 12724 1087 12733
rect 1044 12702 1087 12724
rect 1075 12699 1087 12702
rect 1121 12699 1133 12733
rect 2038 12724 2044 12776
rect 2096 12764 2102 12776
rect 2593 12767 2651 12773
rect 2593 12764 2605 12767
rect 2096 12736 2605 12764
rect 2096 12724 2102 12736
rect 2593 12733 2605 12736
rect 2639 12733 2651 12767
rect 2593 12727 2651 12733
rect 2958 12724 2964 12776
rect 3016 12764 3022 12776
rect 3421 12767 3479 12773
rect 3421 12764 3433 12767
rect 3016 12736 3433 12764
rect 3016 12724 3022 12736
rect 3421 12733 3433 12736
rect 3467 12733 3479 12767
rect 3421 12727 3479 12733
rect 3605 12767 3663 12773
rect 3605 12733 3617 12767
rect 3651 12764 3663 12767
rect 3651 12736 3832 12764
rect 3651 12733 3663 12736
rect 3605 12727 3663 12733
rect 1075 12693 1133 12699
rect 1305 12699 1363 12705
rect 1305 12665 1317 12699
rect 1351 12696 1363 12699
rect 1486 12696 1492 12708
rect 1351 12668 1492 12696
rect 1351 12665 1363 12668
rect 1305 12659 1363 12665
rect 1486 12656 1492 12668
rect 1544 12656 1550 12708
rect 2133 12699 2191 12705
rect 2133 12665 2145 12699
rect 2179 12696 2191 12699
rect 2222 12696 2228 12708
rect 2179 12668 2228 12696
rect 2179 12665 2191 12668
rect 2133 12659 2191 12665
rect 2222 12656 2228 12668
rect 2280 12656 2286 12708
rect 2314 12656 2320 12708
rect 2372 12656 2378 12708
rect 3326 12656 3332 12708
rect 3384 12696 3390 12708
rect 3697 12699 3755 12705
rect 3697 12696 3709 12699
rect 3384 12668 3709 12696
rect 3384 12656 3390 12668
rect 3697 12665 3709 12668
rect 3743 12665 3755 12699
rect 3804 12696 3832 12736
rect 3878 12724 3884 12776
rect 3936 12724 3942 12776
rect 4154 12724 4160 12776
rect 4212 12724 4218 12776
rect 4614 12724 4620 12776
rect 4672 12724 4678 12776
rect 4982 12724 4988 12776
rect 5040 12764 5046 12776
rect 6549 12767 6607 12773
rect 6549 12764 6561 12767
rect 5040 12736 6561 12764
rect 5040 12724 5046 12736
rect 6549 12733 6561 12736
rect 6595 12733 6607 12767
rect 6549 12727 6607 12733
rect 7101 12767 7159 12773
rect 7101 12733 7113 12767
rect 7147 12764 7159 12767
rect 7190 12764 7196 12776
rect 7147 12736 7196 12764
rect 7147 12733 7159 12736
rect 7101 12727 7159 12733
rect 7190 12724 7196 12736
rect 7248 12724 7254 12776
rect 7466 12724 7472 12776
rect 7524 12724 7530 12776
rect 7561 12767 7619 12773
rect 7561 12733 7573 12767
rect 7607 12733 7619 12767
rect 7561 12727 7619 12733
rect 8573 12767 8631 12773
rect 8573 12733 8585 12767
rect 8619 12764 8631 12767
rect 8662 12764 8668 12776
rect 8619 12736 8668 12764
rect 8619 12733 8631 12736
rect 8573 12727 8631 12733
rect 3970 12696 3976 12708
rect 3804 12668 3976 12696
rect 3697 12659 3755 12665
rect 3970 12656 3976 12668
rect 4028 12656 4034 12708
rect 4065 12699 4123 12705
rect 4065 12665 4077 12699
rect 4111 12696 4123 12699
rect 4246 12696 4252 12708
rect 4111 12668 4252 12696
rect 4111 12665 4123 12668
rect 4065 12659 4123 12665
rect 4246 12656 4252 12668
rect 4304 12656 4310 12708
rect 1946 12588 1952 12640
rect 2004 12588 2010 12640
rect 2406 12588 2412 12640
rect 2464 12588 2470 12640
rect 3513 12631 3571 12637
rect 3513 12597 3525 12631
rect 3559 12628 3571 12631
rect 3602 12628 3608 12640
rect 3559 12600 3608 12628
rect 3559 12597 3571 12600
rect 3513 12591 3571 12597
rect 3602 12588 3608 12600
rect 3660 12588 3666 12640
rect 4154 12588 4160 12640
rect 4212 12628 4218 12640
rect 4632 12628 4660 12724
rect 4890 12656 4896 12708
rect 4948 12696 4954 12708
rect 5353 12699 5411 12705
rect 5353 12696 5365 12699
rect 4948 12668 5365 12696
rect 4948 12656 4954 12668
rect 5353 12665 5365 12668
rect 5399 12665 5411 12699
rect 5353 12659 5411 12665
rect 5445 12699 5503 12705
rect 5445 12665 5457 12699
rect 5491 12665 5503 12699
rect 5445 12659 5503 12665
rect 4212 12600 4660 12628
rect 4801 12631 4859 12637
rect 4212 12588 4218 12600
rect 4801 12597 4813 12631
rect 4847 12628 4859 12631
rect 4982 12628 4988 12640
rect 4847 12600 4988 12628
rect 4847 12597 4859 12600
rect 4801 12591 4859 12597
rect 4982 12588 4988 12600
rect 5040 12588 5046 12640
rect 5074 12588 5080 12640
rect 5132 12588 5138 12640
rect 5166 12588 5172 12640
rect 5224 12628 5230 12640
rect 5460 12628 5488 12659
rect 5534 12656 5540 12708
rect 5592 12696 5598 12708
rect 5813 12699 5871 12705
rect 5813 12696 5825 12699
rect 5592 12668 5825 12696
rect 5592 12656 5598 12668
rect 5813 12665 5825 12668
rect 5859 12665 5871 12699
rect 5813 12659 5871 12665
rect 6178 12656 6184 12708
rect 6236 12656 6242 12708
rect 7208 12696 7236 12724
rect 7576 12696 7604 12727
rect 8662 12724 8668 12736
rect 8720 12724 8726 12776
rect 8757 12767 8815 12773
rect 8757 12733 8769 12767
rect 8803 12733 8815 12767
rect 8757 12727 8815 12733
rect 8386 12696 8392 12708
rect 7208 12668 7604 12696
rect 7668 12668 8392 12696
rect 5224 12600 5488 12628
rect 6365 12631 6423 12637
rect 5224 12588 5230 12600
rect 6365 12597 6377 12631
rect 6411 12628 6423 12631
rect 6454 12628 6460 12640
rect 6411 12600 6460 12628
rect 6411 12597 6423 12600
rect 6365 12591 6423 12597
rect 6454 12588 6460 12600
rect 6512 12588 6518 12640
rect 6730 12588 6736 12640
rect 6788 12628 6794 12640
rect 7668 12628 7696 12668
rect 8386 12656 8392 12668
rect 8444 12656 8450 12708
rect 8772 12696 8800 12727
rect 9674 12724 9680 12776
rect 9732 12724 9738 12776
rect 10060 12773 10088 12804
rect 9769 12767 9827 12773
rect 9769 12733 9781 12767
rect 9815 12764 9827 12767
rect 10045 12767 10103 12773
rect 9815 12736 9996 12764
rect 9815 12733 9827 12736
rect 9769 12727 9827 12733
rect 9968 12696 9996 12736
rect 10045 12733 10057 12767
rect 10091 12733 10103 12767
rect 10045 12727 10103 12733
rect 10137 12767 10195 12773
rect 10137 12733 10149 12767
rect 10183 12764 10195 12767
rect 10226 12764 10232 12776
rect 10183 12736 10232 12764
rect 10183 12733 10195 12736
rect 10137 12727 10195 12733
rect 10226 12724 10232 12736
rect 10284 12724 10290 12776
rect 10321 12767 10379 12773
rect 10321 12733 10333 12767
rect 10367 12764 10379 12767
rect 10502 12764 10508 12776
rect 10367 12736 10508 12764
rect 10367 12733 10379 12736
rect 10321 12727 10379 12733
rect 10502 12724 10508 12736
rect 10560 12724 10566 12776
rect 11164 12773 11192 12804
rect 11256 12804 11336 12832
rect 11256 12773 11284 12804
rect 11330 12792 11336 12804
rect 11388 12792 11394 12844
rect 11425 12835 11483 12841
rect 11425 12801 11437 12835
rect 11471 12832 11483 12835
rect 12544 12832 12572 12872
rect 12618 12860 12624 12912
rect 12676 12900 12682 12912
rect 13081 12903 13139 12909
rect 13081 12900 13093 12903
rect 12676 12872 13093 12900
rect 12676 12860 12682 12872
rect 13081 12869 13093 12872
rect 13127 12869 13139 12903
rect 14458 12900 14464 12912
rect 13081 12863 13139 12869
rect 13188 12872 14464 12900
rect 13188 12832 13216 12872
rect 14458 12860 14464 12872
rect 14516 12860 14522 12912
rect 14553 12903 14611 12909
rect 14553 12869 14565 12903
rect 14599 12869 14611 12903
rect 14553 12863 14611 12869
rect 11471 12804 12480 12832
rect 12544 12804 13216 12832
rect 14093 12835 14151 12841
rect 11471 12801 11483 12804
rect 11425 12795 11483 12801
rect 11149 12767 11207 12773
rect 11149 12733 11161 12767
rect 11195 12733 11207 12767
rect 11149 12727 11207 12733
rect 11241 12767 11299 12773
rect 11241 12733 11253 12767
rect 11287 12733 11299 12767
rect 11517 12767 11575 12773
rect 11517 12764 11529 12767
rect 11241 12727 11299 12733
rect 11440 12736 11529 12764
rect 8772 12668 9812 12696
rect 9968 12668 10364 12696
rect 9784 12640 9812 12668
rect 6788 12600 7696 12628
rect 7745 12631 7803 12637
rect 6788 12588 6794 12600
rect 7745 12597 7757 12631
rect 7791 12628 7803 12631
rect 8294 12628 8300 12640
rect 7791 12600 8300 12628
rect 7791 12597 7803 12600
rect 7745 12591 7803 12597
rect 8294 12588 8300 12600
rect 8352 12588 8358 12640
rect 8665 12631 8723 12637
rect 8665 12597 8677 12631
rect 8711 12628 8723 12631
rect 8846 12628 8852 12640
rect 8711 12600 8852 12628
rect 8711 12597 8723 12600
rect 8665 12591 8723 12597
rect 8846 12588 8852 12600
rect 8904 12588 8910 12640
rect 9766 12588 9772 12640
rect 9824 12588 9830 12640
rect 10336 12637 10364 12668
rect 11440 12640 11468 12736
rect 11517 12733 11529 12736
rect 11563 12733 11575 12767
rect 11517 12727 11575 12733
rect 12066 12724 12072 12776
rect 12124 12724 12130 12776
rect 12342 12724 12348 12776
rect 12400 12724 12406 12776
rect 12452 12764 12480 12804
rect 14093 12801 14105 12835
rect 14139 12801 14151 12835
rect 14568 12832 14596 12863
rect 15102 12860 15108 12912
rect 15160 12900 15166 12912
rect 15197 12903 15255 12909
rect 15197 12900 15209 12903
rect 15160 12872 15209 12900
rect 15160 12860 15166 12872
rect 15197 12869 15209 12872
rect 15243 12869 15255 12903
rect 15197 12863 15255 12869
rect 15010 12832 15016 12844
rect 14568 12804 15016 12832
rect 14093 12795 14151 12801
rect 12452 12736 12756 12764
rect 10321 12631 10379 12637
rect 10321 12597 10333 12631
rect 10367 12628 10379 12631
rect 11422 12628 11428 12640
rect 10367 12600 11428 12628
rect 10367 12597 10379 12600
rect 10321 12591 10379 12597
rect 11422 12588 11428 12600
rect 11480 12588 11486 12640
rect 12161 12631 12219 12637
rect 12161 12597 12173 12631
rect 12207 12628 12219 12631
rect 12434 12628 12440 12640
rect 12207 12600 12440 12628
rect 12207 12597 12219 12600
rect 12161 12591 12219 12597
rect 12434 12588 12440 12600
rect 12492 12588 12498 12640
rect 12728 12628 12756 12736
rect 12802 12724 12808 12776
rect 12860 12764 12866 12776
rect 12897 12767 12955 12773
rect 12897 12764 12909 12767
rect 12860 12736 12909 12764
rect 12860 12724 12866 12736
rect 12897 12733 12909 12736
rect 12943 12733 12955 12767
rect 12897 12727 12955 12733
rect 14108 12696 14136 12795
rect 15010 12792 15016 12804
rect 15068 12832 15074 12844
rect 15068 12804 15148 12832
rect 15068 12792 15074 12804
rect 14182 12724 14188 12776
rect 14240 12764 14246 12776
rect 15120 12773 15148 12804
rect 15396 12776 15424 12940
rect 19429 12937 19441 12940
rect 19475 12937 19487 12971
rect 19429 12931 19487 12937
rect 19886 12928 19892 12980
rect 19944 12968 19950 12980
rect 19944 12940 20576 12968
rect 19944 12928 19950 12940
rect 16853 12903 16911 12909
rect 16853 12869 16865 12903
rect 16899 12900 16911 12903
rect 17218 12900 17224 12912
rect 16899 12872 17224 12900
rect 16899 12869 16911 12872
rect 16853 12863 16911 12869
rect 17218 12860 17224 12872
rect 17276 12900 17282 12912
rect 17405 12903 17463 12909
rect 17405 12900 17417 12903
rect 17276 12872 17417 12900
rect 17276 12860 17282 12872
rect 17405 12869 17417 12872
rect 17451 12869 17463 12903
rect 17405 12863 17463 12869
rect 18506 12860 18512 12912
rect 18564 12900 18570 12912
rect 20073 12903 20131 12909
rect 20073 12900 20085 12903
rect 18564 12872 20085 12900
rect 18564 12860 18570 12872
rect 20073 12869 20085 12872
rect 20119 12869 20131 12903
rect 20073 12863 20131 12869
rect 17589 12835 17647 12841
rect 16960 12804 17356 12832
rect 16960 12776 16988 12804
rect 14829 12767 14887 12773
rect 14829 12764 14841 12767
rect 14240 12736 14841 12764
rect 14240 12724 14246 12736
rect 14829 12733 14841 12736
rect 14875 12733 14887 12767
rect 14829 12727 14887 12733
rect 15105 12767 15163 12773
rect 15105 12733 15117 12767
rect 15151 12733 15163 12767
rect 15105 12727 15163 12733
rect 15378 12724 15384 12776
rect 15436 12724 15442 12776
rect 15470 12724 15476 12776
rect 15528 12764 15534 12776
rect 16761 12767 16819 12773
rect 16761 12764 16773 12767
rect 15528 12736 16773 12764
rect 15528 12724 15534 12736
rect 16761 12733 16773 12736
rect 16807 12764 16819 12767
rect 16850 12764 16856 12776
rect 16807 12736 16856 12764
rect 16807 12733 16819 12736
rect 16761 12727 16819 12733
rect 16850 12724 16856 12736
rect 16908 12724 16914 12776
rect 16942 12724 16948 12776
rect 17000 12724 17006 12776
rect 17328 12773 17356 12804
rect 17589 12801 17601 12835
rect 17635 12801 17647 12835
rect 17589 12795 17647 12801
rect 17037 12767 17095 12773
rect 17037 12733 17049 12767
rect 17083 12733 17095 12767
rect 17037 12727 17095 12733
rect 17313 12767 17371 12773
rect 17313 12733 17325 12767
rect 17359 12733 17371 12767
rect 17313 12727 17371 12733
rect 15013 12699 15071 12705
rect 15013 12696 15025 12699
rect 14108 12668 15025 12696
rect 15013 12665 15025 12668
rect 15059 12696 15071 12699
rect 15194 12696 15200 12708
rect 15059 12668 15200 12696
rect 15059 12665 15071 12668
rect 15013 12659 15071 12665
rect 15194 12656 15200 12668
rect 15252 12656 15258 12708
rect 15286 12656 15292 12708
rect 15344 12656 15350 12708
rect 17052 12696 17080 12727
rect 17604 12696 17632 12795
rect 18782 12792 18788 12844
rect 18840 12792 18846 12844
rect 19245 12835 19303 12841
rect 19245 12801 19257 12835
rect 19291 12832 19303 12835
rect 19426 12832 19432 12844
rect 19291 12804 19432 12832
rect 19291 12801 19303 12804
rect 19245 12795 19303 12801
rect 19426 12792 19432 12804
rect 19484 12792 19490 12844
rect 20438 12792 20444 12844
rect 20496 12832 20502 12844
rect 20548 12841 20576 12940
rect 20533 12835 20591 12841
rect 20533 12832 20545 12835
rect 20496 12804 20545 12832
rect 20496 12792 20502 12804
rect 20533 12801 20545 12804
rect 20579 12801 20591 12835
rect 20533 12795 20591 12801
rect 20717 12835 20775 12841
rect 20717 12801 20729 12835
rect 20763 12832 20775 12835
rect 20990 12832 20996 12844
rect 20763 12804 20996 12832
rect 20763 12801 20775 12804
rect 20717 12795 20775 12801
rect 20990 12792 20996 12804
rect 21048 12792 21054 12844
rect 18874 12724 18880 12776
rect 18932 12764 18938 12776
rect 19518 12773 19524 12776
rect 19337 12767 19395 12773
rect 19337 12764 19349 12767
rect 18932 12736 19349 12764
rect 18932 12724 18938 12736
rect 19337 12733 19349 12736
rect 19383 12733 19395 12767
rect 19514 12764 19524 12773
rect 19479 12736 19524 12764
rect 19337 12727 19395 12733
rect 19514 12727 19524 12736
rect 19518 12724 19524 12727
rect 19576 12724 19582 12776
rect 19886 12724 19892 12776
rect 19944 12724 19950 12776
rect 20070 12724 20076 12776
rect 20128 12724 20134 12776
rect 20806 12724 20812 12776
rect 20864 12724 20870 12776
rect 21361 12767 21419 12773
rect 21361 12733 21373 12767
rect 21407 12764 21419 12767
rect 21407 12736 21772 12764
rect 21407 12733 21419 12736
rect 21361 12727 21419 12733
rect 21744 12708 21772 12736
rect 17052 12668 21404 12696
rect 14366 12628 14372 12640
rect 12728 12600 14372 12628
rect 14366 12588 14372 12600
rect 14424 12588 14430 12640
rect 14458 12588 14464 12640
rect 14516 12628 14522 12640
rect 16022 12628 16028 12640
rect 14516 12600 16028 12628
rect 14516 12588 14522 12600
rect 16022 12588 16028 12600
rect 16080 12588 16086 12640
rect 17126 12588 17132 12640
rect 17184 12628 17190 12640
rect 17221 12631 17279 12637
rect 17221 12628 17233 12631
rect 17184 12600 17233 12628
rect 17184 12588 17190 12600
rect 17221 12597 17233 12600
rect 17267 12597 17279 12631
rect 17221 12591 17279 12597
rect 17586 12588 17592 12640
rect 17644 12588 17650 12640
rect 18782 12588 18788 12640
rect 18840 12628 18846 12640
rect 19288 12628 19294 12640
rect 18840 12600 19294 12628
rect 18840 12588 18846 12600
rect 19288 12588 19294 12600
rect 19346 12588 19352 12640
rect 21177 12631 21235 12637
rect 21177 12597 21189 12631
rect 21223 12628 21235 12631
rect 21266 12628 21272 12640
rect 21223 12600 21272 12628
rect 21223 12597 21235 12600
rect 21177 12591 21235 12597
rect 21266 12588 21272 12600
rect 21324 12588 21330 12640
rect 21376 12628 21404 12668
rect 21450 12656 21456 12708
rect 21508 12696 21514 12708
rect 21606 12699 21664 12705
rect 21606 12696 21618 12699
rect 21508 12668 21618 12696
rect 21508 12656 21514 12668
rect 21606 12665 21618 12668
rect 21652 12665 21664 12699
rect 21606 12659 21664 12665
rect 21726 12656 21732 12708
rect 21784 12656 21790 12708
rect 21818 12628 21824 12640
rect 21376 12600 21824 12628
rect 21818 12588 21824 12600
rect 21876 12588 21882 12640
rect 22094 12588 22100 12640
rect 22152 12628 22158 12640
rect 22741 12631 22799 12637
rect 22741 12628 22753 12631
rect 22152 12600 22753 12628
rect 22152 12588 22158 12600
rect 22741 12597 22753 12600
rect 22787 12597 22799 12631
rect 22741 12591 22799 12597
rect 552 12538 23368 12560
rect 552 12486 4366 12538
rect 4418 12486 4430 12538
rect 4482 12486 4494 12538
rect 4546 12486 4558 12538
rect 4610 12486 4622 12538
rect 4674 12486 4686 12538
rect 4738 12486 10366 12538
rect 10418 12486 10430 12538
rect 10482 12486 10494 12538
rect 10546 12486 10558 12538
rect 10610 12486 10622 12538
rect 10674 12486 10686 12538
rect 10738 12486 16366 12538
rect 16418 12486 16430 12538
rect 16482 12486 16494 12538
rect 16546 12486 16558 12538
rect 16610 12486 16622 12538
rect 16674 12486 16686 12538
rect 16738 12486 22366 12538
rect 22418 12486 22430 12538
rect 22482 12486 22494 12538
rect 22546 12486 22558 12538
rect 22610 12486 22622 12538
rect 22674 12486 22686 12538
rect 22738 12486 23368 12538
rect 552 12464 23368 12486
rect 937 12427 995 12433
rect 937 12393 949 12427
rect 983 12424 995 12427
rect 1026 12424 1032 12436
rect 983 12396 1032 12424
rect 983 12393 995 12396
rect 937 12387 995 12393
rect 1026 12384 1032 12396
rect 1084 12384 1090 12436
rect 1765 12427 1823 12433
rect 1765 12393 1777 12427
rect 1811 12424 1823 12427
rect 1946 12424 1952 12436
rect 1811 12396 1952 12424
rect 1811 12393 1823 12396
rect 1765 12387 1823 12393
rect 1946 12384 1952 12396
rect 2004 12384 2010 12436
rect 2222 12384 2228 12436
rect 2280 12384 2286 12436
rect 3694 12384 3700 12436
rect 3752 12384 3758 12436
rect 4890 12424 4896 12436
rect 4264 12396 4896 12424
rect 1670 12356 1676 12368
rect 1136 12328 1676 12356
rect 1136 12297 1164 12328
rect 1670 12316 1676 12328
rect 1728 12316 1734 12368
rect 1121 12291 1179 12297
rect 1121 12257 1133 12291
rect 1167 12257 1179 12291
rect 1121 12251 1179 12257
rect 1210 12248 1216 12300
rect 1268 12288 1274 12300
rect 2041 12291 2099 12297
rect 2041 12288 2053 12291
rect 1268 12260 2053 12288
rect 1268 12248 1274 12260
rect 2041 12257 2053 12260
rect 2087 12257 2099 12291
rect 2240 12288 2268 12384
rect 2308 12359 2366 12365
rect 2308 12325 2320 12359
rect 2354 12356 2366 12359
rect 2406 12356 2412 12368
rect 2354 12328 2412 12356
rect 2354 12325 2366 12328
rect 2308 12319 2366 12325
rect 2406 12316 2412 12328
rect 2464 12316 2470 12368
rect 3712 12356 3740 12384
rect 4062 12356 4068 12368
rect 3712 12328 4068 12356
rect 4062 12316 4068 12328
rect 4120 12316 4126 12368
rect 2041 12251 2099 12257
rect 2148 12260 2268 12288
rect 1305 12223 1363 12229
rect 1305 12189 1317 12223
rect 1351 12220 1363 12223
rect 2148 12220 2176 12260
rect 3418 12248 3424 12300
rect 3476 12288 3482 12300
rect 3513 12291 3571 12297
rect 3513 12288 3525 12291
rect 3476 12260 3525 12288
rect 3476 12248 3482 12260
rect 3513 12257 3525 12260
rect 3559 12257 3571 12291
rect 3513 12251 3571 12257
rect 3602 12248 3608 12300
rect 3660 12288 3666 12300
rect 3697 12291 3755 12297
rect 3697 12288 3709 12291
rect 3660 12260 3709 12288
rect 3660 12248 3666 12260
rect 3697 12257 3709 12260
rect 3743 12257 3755 12291
rect 3697 12251 3755 12257
rect 3789 12291 3847 12297
rect 3789 12257 3801 12291
rect 3835 12257 3847 12291
rect 3789 12251 3847 12257
rect 1351 12192 2176 12220
rect 3804 12220 3832 12251
rect 3878 12248 3884 12300
rect 3936 12288 3942 12300
rect 4154 12288 4160 12300
rect 3936 12260 4160 12288
rect 3936 12248 3942 12260
rect 4154 12248 4160 12260
rect 4212 12248 4218 12300
rect 4264 12297 4292 12396
rect 4890 12384 4896 12396
rect 4948 12424 4954 12436
rect 6270 12424 6276 12436
rect 4948 12396 6276 12424
rect 4948 12384 4954 12396
rect 6270 12384 6276 12396
rect 6328 12384 6334 12436
rect 7466 12384 7472 12436
rect 7524 12424 7530 12436
rect 9674 12424 9680 12436
rect 7524 12396 9680 12424
rect 7524 12384 7530 12396
rect 9674 12384 9680 12396
rect 9732 12384 9738 12436
rect 11422 12384 11428 12436
rect 11480 12424 11486 12436
rect 15194 12424 15200 12436
rect 11480 12396 15200 12424
rect 11480 12384 11486 12396
rect 15194 12384 15200 12396
rect 15252 12384 15258 12436
rect 15289 12427 15347 12433
rect 15289 12393 15301 12427
rect 15335 12424 15347 12427
rect 15378 12424 15384 12436
rect 15335 12396 15384 12424
rect 15335 12393 15347 12396
rect 15289 12387 15347 12393
rect 15378 12384 15384 12396
rect 15436 12384 15442 12436
rect 15746 12384 15752 12436
rect 15804 12424 15810 12436
rect 16298 12424 16304 12436
rect 15804 12396 16304 12424
rect 15804 12384 15810 12396
rect 16298 12384 16304 12396
rect 16356 12384 16362 12436
rect 17037 12427 17095 12433
rect 16408 12396 16988 12424
rect 4433 12359 4491 12365
rect 4433 12325 4445 12359
rect 4479 12356 4491 12359
rect 4709 12359 4767 12365
rect 4479 12328 4660 12356
rect 4479 12325 4491 12328
rect 4433 12319 4491 12325
rect 4249 12291 4307 12297
rect 4249 12257 4261 12291
rect 4295 12257 4307 12291
rect 4249 12251 4307 12257
rect 4338 12248 4344 12300
rect 4396 12248 4402 12300
rect 4632 12297 4660 12328
rect 4709 12325 4721 12359
rect 4755 12356 4767 12359
rect 7745 12359 7803 12365
rect 7745 12356 7757 12359
rect 4755 12328 6040 12356
rect 4755 12325 4767 12328
rect 4709 12319 4767 12325
rect 4525 12291 4583 12297
rect 4525 12257 4537 12291
rect 4571 12257 4583 12291
rect 4525 12251 4583 12257
rect 4617 12291 4675 12297
rect 4617 12257 4629 12291
rect 4663 12257 4675 12291
rect 4617 12251 4675 12257
rect 4801 12291 4859 12297
rect 4801 12257 4813 12291
rect 4847 12288 4859 12291
rect 5074 12288 5080 12300
rect 4847 12260 5080 12288
rect 4847 12257 4859 12260
rect 4801 12251 4859 12257
rect 3804 12192 4292 12220
rect 1351 12189 1363 12192
rect 1305 12183 1363 12189
rect 4264 12164 4292 12192
rect 842 12112 848 12164
rect 900 12152 906 12164
rect 1026 12152 1032 12164
rect 900 12124 1032 12152
rect 900 12112 906 12124
rect 1026 12112 1032 12124
rect 1084 12152 1090 12164
rect 1397 12155 1455 12161
rect 1397 12152 1409 12155
rect 1084 12124 1409 12152
rect 1084 12112 1090 12124
rect 1397 12121 1409 12124
rect 1443 12121 1455 12155
rect 1397 12115 1455 12121
rect 1949 12155 2007 12161
rect 1949 12121 1961 12155
rect 1995 12152 2007 12155
rect 2038 12152 2044 12164
rect 1995 12124 2044 12152
rect 1995 12121 2007 12124
rect 1949 12115 2007 12121
rect 2038 12112 2044 12124
rect 2096 12112 2102 12164
rect 3421 12155 3479 12161
rect 3421 12121 3433 12155
rect 3467 12152 3479 12155
rect 4154 12152 4160 12164
rect 3467 12124 4160 12152
rect 3467 12121 3479 12124
rect 3421 12115 3479 12121
rect 1765 12087 1823 12093
rect 1765 12053 1777 12087
rect 1811 12084 1823 12087
rect 2222 12084 2228 12096
rect 1811 12056 2228 12084
rect 1811 12053 1823 12056
rect 1765 12047 1823 12053
rect 2222 12044 2228 12056
rect 2280 12044 2286 12096
rect 2774 12044 2780 12096
rect 2832 12084 2838 12096
rect 3436 12084 3464 12115
rect 4154 12112 4160 12124
rect 4212 12112 4218 12164
rect 4246 12112 4252 12164
rect 4304 12112 4310 12164
rect 4540 12152 4568 12251
rect 4632 12220 4660 12251
rect 5074 12248 5080 12260
rect 5132 12288 5138 12300
rect 6012 12297 6040 12328
rect 7024 12328 7757 12356
rect 7024 12300 7052 12328
rect 7745 12325 7757 12328
rect 7791 12325 7803 12359
rect 8478 12356 8484 12368
rect 7745 12319 7803 12325
rect 8312 12328 8484 12356
rect 5445 12291 5503 12297
rect 5445 12288 5457 12291
rect 5132 12260 5457 12288
rect 5132 12248 5138 12260
rect 5445 12257 5457 12260
rect 5491 12257 5503 12291
rect 5445 12251 5503 12257
rect 5997 12291 6055 12297
rect 5997 12257 6009 12291
rect 6043 12257 6055 12291
rect 5997 12251 6055 12257
rect 6549 12291 6607 12297
rect 6549 12257 6561 12291
rect 6595 12257 6607 12291
rect 6549 12251 6607 12257
rect 4893 12223 4951 12229
rect 4893 12220 4905 12223
rect 4632 12192 4905 12220
rect 4893 12189 4905 12192
rect 4939 12189 4951 12223
rect 5537 12223 5595 12229
rect 4893 12183 4951 12189
rect 5092 12192 5488 12220
rect 5092 12152 5120 12192
rect 4540 12124 5120 12152
rect 5169 12155 5227 12161
rect 5169 12121 5181 12155
rect 5215 12152 5227 12155
rect 5258 12152 5264 12164
rect 5215 12124 5264 12152
rect 5215 12121 5227 12124
rect 5169 12115 5227 12121
rect 5258 12112 5264 12124
rect 5316 12112 5322 12164
rect 5460 12152 5488 12192
rect 5537 12189 5549 12223
rect 5583 12220 5595 12223
rect 5902 12220 5908 12232
rect 5583 12192 5908 12220
rect 5583 12189 5595 12192
rect 5537 12183 5595 12189
rect 5902 12180 5908 12192
rect 5960 12180 5966 12232
rect 6564 12220 6592 12251
rect 6730 12248 6736 12300
rect 6788 12248 6794 12300
rect 7006 12248 7012 12300
rect 7064 12248 7070 12300
rect 7285 12291 7343 12297
rect 7285 12257 7297 12291
rect 7331 12257 7343 12291
rect 7285 12251 7343 12257
rect 6012 12192 6592 12220
rect 6641 12223 6699 12229
rect 5810 12152 5816 12164
rect 5460 12124 5816 12152
rect 5810 12112 5816 12124
rect 5868 12112 5874 12164
rect 2832 12056 3464 12084
rect 3697 12087 3755 12093
rect 2832 12044 2838 12056
rect 3697 12053 3709 12087
rect 3743 12084 3755 12087
rect 3786 12084 3792 12096
rect 3743 12056 3792 12084
rect 3743 12053 3755 12056
rect 3697 12047 3755 12053
rect 3786 12044 3792 12056
rect 3844 12044 3850 12096
rect 3970 12044 3976 12096
rect 4028 12044 4034 12096
rect 4062 12044 4068 12096
rect 4120 12044 4126 12096
rect 4264 12084 4292 12112
rect 6012 12084 6040 12192
rect 6641 12189 6653 12223
rect 6687 12220 6699 12223
rect 7300 12220 7328 12251
rect 7466 12248 7472 12300
rect 7524 12248 7530 12300
rect 8312 12297 8340 12328
rect 8478 12316 8484 12328
rect 8536 12356 8542 12368
rect 8536 12328 9168 12356
rect 8536 12316 8542 12328
rect 7561 12291 7619 12297
rect 7561 12257 7573 12291
rect 7607 12257 7619 12291
rect 7561 12251 7619 12257
rect 8297 12291 8355 12297
rect 8297 12257 8309 12291
rect 8343 12257 8355 12291
rect 8297 12251 8355 12257
rect 7576 12220 7604 12251
rect 8386 12248 8392 12300
rect 8444 12248 8450 12300
rect 8570 12248 8576 12300
rect 8628 12288 8634 12300
rect 8665 12291 8723 12297
rect 8665 12288 8677 12291
rect 8628 12260 8677 12288
rect 8628 12248 8634 12260
rect 8665 12257 8677 12260
rect 8711 12257 8723 12291
rect 8665 12251 8723 12257
rect 8757 12291 8815 12297
rect 8757 12257 8769 12291
rect 8803 12257 8815 12291
rect 8757 12251 8815 12257
rect 6687 12192 7604 12220
rect 6687 12189 6699 12192
rect 6641 12183 6699 12189
rect 6365 12155 6423 12161
rect 6365 12121 6377 12155
rect 6411 12152 6423 12155
rect 7006 12152 7012 12164
rect 6411 12124 7012 12152
rect 6411 12121 6423 12124
rect 6365 12115 6423 12121
rect 7006 12112 7012 12124
rect 7064 12112 7070 12164
rect 8772 12096 8800 12251
rect 8846 12248 8852 12300
rect 8904 12248 8910 12300
rect 9140 12297 9168 12328
rect 11054 12316 11060 12368
rect 11112 12356 11118 12368
rect 12066 12356 12072 12368
rect 11112 12328 12072 12356
rect 11112 12316 11118 12328
rect 9125 12291 9183 12297
rect 9125 12257 9137 12291
rect 9171 12288 9183 12291
rect 11606 12288 11612 12300
rect 9171 12260 11612 12288
rect 9171 12257 9183 12260
rect 9125 12251 9183 12257
rect 11606 12248 11612 12260
rect 11664 12248 11670 12300
rect 11716 12297 11744 12328
rect 12066 12316 12072 12328
rect 12124 12316 12130 12368
rect 12710 12356 12716 12368
rect 12406 12328 12716 12356
rect 11701 12291 11759 12297
rect 11701 12257 11713 12291
rect 11747 12257 11759 12291
rect 11701 12251 11759 12257
rect 11790 12248 11796 12300
rect 11848 12248 11854 12300
rect 12406 12288 12434 12328
rect 11900 12260 12434 12288
rect 9214 12180 9220 12232
rect 9272 12220 9278 12232
rect 11900 12220 11928 12260
rect 9272 12192 11928 12220
rect 9272 12180 9278 12192
rect 12250 12180 12256 12232
rect 12308 12180 12314 12232
rect 12544 12229 12572 12328
rect 12710 12316 12716 12328
rect 12768 12316 12774 12368
rect 14090 12356 14096 12368
rect 12820 12328 14096 12356
rect 12621 12291 12679 12297
rect 12621 12257 12633 12291
rect 12667 12288 12679 12291
rect 12820 12288 12848 12328
rect 14090 12316 14096 12328
rect 14148 12316 14154 12368
rect 14826 12316 14832 12368
rect 14884 12356 14890 12368
rect 15473 12359 15531 12365
rect 15473 12356 15485 12359
rect 14884 12328 15485 12356
rect 14884 12316 14890 12328
rect 15473 12325 15485 12328
rect 15519 12325 15531 12359
rect 15930 12356 15936 12368
rect 15473 12319 15531 12325
rect 15580 12328 15936 12356
rect 12667 12260 12848 12288
rect 13357 12291 13415 12297
rect 12667 12257 12679 12260
rect 12621 12251 12679 12257
rect 13357 12257 13369 12291
rect 13403 12288 13415 12291
rect 14458 12288 14464 12300
rect 13403 12260 14464 12288
rect 13403 12257 13415 12260
rect 13357 12251 13415 12257
rect 14108 12232 14136 12260
rect 14458 12248 14464 12260
rect 14516 12248 14522 12300
rect 15010 12248 15016 12300
rect 15068 12288 15074 12300
rect 15105 12291 15163 12297
rect 15105 12288 15117 12291
rect 15068 12260 15117 12288
rect 15068 12248 15074 12260
rect 15105 12257 15117 12260
rect 15151 12257 15163 12291
rect 15105 12251 15163 12257
rect 15286 12248 15292 12300
rect 15344 12288 15350 12300
rect 15381 12291 15439 12297
rect 15381 12288 15393 12291
rect 15344 12260 15393 12288
rect 15344 12248 15350 12260
rect 15381 12257 15393 12260
rect 15427 12288 15439 12291
rect 15580 12288 15608 12328
rect 15930 12316 15936 12328
rect 15988 12316 15994 12368
rect 16408 12356 16436 12396
rect 16316 12328 16436 12356
rect 16316 12300 16344 12328
rect 16482 12316 16488 12368
rect 16540 12316 16546 12368
rect 16592 12328 16804 12356
rect 15427 12260 15608 12288
rect 15657 12291 15715 12297
rect 15427 12257 15439 12260
rect 15381 12251 15439 12257
rect 15657 12257 15669 12291
rect 15703 12257 15715 12291
rect 15657 12251 15715 12257
rect 12529 12223 12587 12229
rect 12529 12189 12541 12223
rect 12575 12189 12587 12223
rect 12529 12183 12587 12189
rect 12989 12223 13047 12229
rect 12989 12189 13001 12223
rect 13035 12220 13047 12223
rect 13262 12220 13268 12232
rect 13035 12192 13268 12220
rect 13035 12189 13047 12192
rect 12989 12183 13047 12189
rect 13262 12180 13268 12192
rect 13320 12180 13326 12232
rect 14090 12180 14096 12232
rect 14148 12180 14154 12232
rect 14274 12180 14280 12232
rect 14332 12220 14338 12232
rect 15672 12220 15700 12251
rect 16298 12248 16304 12300
rect 16356 12248 16362 12300
rect 16390 12248 16396 12300
rect 16448 12248 16454 12300
rect 14332 12192 15700 12220
rect 14332 12180 14338 12192
rect 9030 12112 9036 12164
rect 9088 12152 9094 12164
rect 10778 12152 10784 12164
rect 9088 12124 10784 12152
rect 9088 12112 9094 12124
rect 10778 12112 10784 12124
rect 10836 12112 10842 12164
rect 10870 12112 10876 12164
rect 10928 12152 10934 12164
rect 12066 12152 12072 12164
rect 10928 12124 12072 12152
rect 10928 12112 10934 12124
rect 12066 12112 12072 12124
rect 12124 12112 12130 12164
rect 12618 12112 12624 12164
rect 12676 12152 12682 12164
rect 12676 12124 14780 12152
rect 12676 12112 12682 12124
rect 14752 12096 14780 12124
rect 4264 12056 6040 12084
rect 6638 12044 6644 12096
rect 6696 12084 6702 12096
rect 6825 12087 6883 12093
rect 6825 12084 6837 12087
rect 6696 12056 6837 12084
rect 6696 12044 6702 12056
rect 6825 12053 6837 12056
rect 6871 12053 6883 12087
rect 6825 12047 6883 12053
rect 7098 12044 7104 12096
rect 7156 12084 7162 12096
rect 7929 12087 7987 12093
rect 7929 12084 7941 12087
rect 7156 12056 7941 12084
rect 7156 12044 7162 12056
rect 7929 12053 7941 12056
rect 7975 12053 7987 12087
rect 7929 12047 7987 12053
rect 8570 12044 8576 12096
rect 8628 12044 8634 12096
rect 8754 12044 8760 12096
rect 8812 12044 8818 12096
rect 8846 12044 8852 12096
rect 8904 12084 8910 12096
rect 8941 12087 8999 12093
rect 8941 12084 8953 12087
rect 8904 12056 8953 12084
rect 8904 12044 8910 12056
rect 8941 12053 8953 12056
rect 8987 12053 8999 12087
rect 8941 12047 8999 12053
rect 9766 12044 9772 12096
rect 9824 12084 9830 12096
rect 11422 12084 11428 12096
rect 9824 12056 11428 12084
rect 9824 12044 9830 12056
rect 11422 12044 11428 12056
rect 11480 12044 11486 12096
rect 13633 12087 13691 12093
rect 13633 12053 13645 12087
rect 13679 12084 13691 12087
rect 13814 12084 13820 12096
rect 13679 12056 13820 12084
rect 13679 12053 13691 12056
rect 13633 12047 13691 12053
rect 13814 12044 13820 12056
rect 13872 12044 13878 12096
rect 14734 12044 14740 12096
rect 14792 12084 14798 12096
rect 14921 12087 14979 12093
rect 14921 12084 14933 12087
rect 14792 12056 14933 12084
rect 14792 12044 14798 12056
rect 14921 12053 14933 12056
rect 14967 12053 14979 12087
rect 14921 12047 14979 12053
rect 15010 12044 15016 12096
rect 15068 12084 15074 12096
rect 15120 12084 15148 12192
rect 15654 12112 15660 12164
rect 15712 12152 15718 12164
rect 16592 12152 16620 12328
rect 16776 12297 16804 12328
rect 16669 12291 16727 12297
rect 16669 12257 16681 12291
rect 16715 12257 16727 12291
rect 16669 12251 16727 12257
rect 16761 12291 16819 12297
rect 16761 12257 16773 12291
rect 16807 12257 16819 12291
rect 16761 12251 16819 12257
rect 16684 12220 16712 12251
rect 16850 12248 16856 12300
rect 16908 12248 16914 12300
rect 16684 12192 16896 12220
rect 16868 12161 16896 12192
rect 15712 12124 16620 12152
rect 16853 12155 16911 12161
rect 15712 12112 15718 12124
rect 16853 12121 16865 12155
rect 16899 12121 16911 12155
rect 16960 12152 16988 12396
rect 17037 12393 17049 12427
rect 17083 12424 17095 12427
rect 17586 12424 17592 12436
rect 17083 12396 17592 12424
rect 17083 12393 17095 12396
rect 17037 12387 17095 12393
rect 17586 12384 17592 12396
rect 17644 12384 17650 12436
rect 17770 12384 17776 12436
rect 17828 12424 17834 12436
rect 18233 12427 18291 12433
rect 18233 12424 18245 12427
rect 17828 12396 18245 12424
rect 17828 12384 17834 12396
rect 18233 12393 18245 12396
rect 18279 12393 18291 12427
rect 18233 12387 18291 12393
rect 18417 12427 18475 12433
rect 18417 12393 18429 12427
rect 18463 12424 18475 12427
rect 18690 12424 18696 12436
rect 18463 12396 18696 12424
rect 18463 12393 18475 12396
rect 18417 12387 18475 12393
rect 18432 12356 18460 12387
rect 18690 12384 18696 12396
rect 18748 12384 18754 12436
rect 19886 12384 19892 12436
rect 19944 12384 19950 12436
rect 20346 12384 20352 12436
rect 20404 12384 20410 12436
rect 21450 12384 21456 12436
rect 21508 12384 21514 12436
rect 19904 12356 19932 12384
rect 17788 12328 18460 12356
rect 19352 12328 19932 12356
rect 17126 12248 17132 12300
rect 17184 12248 17190 12300
rect 17788 12297 17816 12328
rect 17773 12291 17831 12297
rect 17773 12257 17785 12291
rect 17819 12257 17831 12291
rect 17773 12251 17831 12257
rect 17957 12291 18015 12297
rect 17957 12257 17969 12291
rect 18003 12257 18015 12291
rect 17957 12251 18015 12257
rect 17972 12220 18000 12251
rect 18046 12248 18052 12300
rect 18104 12248 18110 12300
rect 18322 12248 18328 12300
rect 18380 12248 18386 12300
rect 18601 12291 18659 12297
rect 18601 12257 18613 12291
rect 18647 12288 18659 12291
rect 18690 12288 18696 12300
rect 18647 12260 18696 12288
rect 18647 12257 18659 12260
rect 18601 12251 18659 12257
rect 18690 12248 18696 12260
rect 18748 12248 18754 12300
rect 19352 12297 19380 12328
rect 19245 12291 19303 12297
rect 19245 12257 19257 12291
rect 19291 12257 19303 12291
rect 19245 12251 19303 12257
rect 19337 12291 19395 12297
rect 19337 12257 19349 12291
rect 19383 12257 19395 12291
rect 19337 12251 19395 12257
rect 18340 12220 18368 12248
rect 17972 12192 18368 12220
rect 19260 12220 19288 12251
rect 19426 12248 19432 12300
rect 19484 12248 19490 12300
rect 19518 12248 19524 12300
rect 19576 12248 19582 12300
rect 19978 12248 19984 12300
rect 20036 12288 20042 12300
rect 20073 12291 20131 12297
rect 20073 12288 20085 12291
rect 20036 12260 20085 12288
rect 20036 12248 20042 12260
rect 20073 12257 20085 12260
rect 20119 12257 20131 12291
rect 20073 12251 20131 12257
rect 20162 12220 20168 12232
rect 19260 12192 20168 12220
rect 20162 12180 20168 12192
rect 20220 12180 20226 12232
rect 20254 12180 20260 12232
rect 20312 12220 20318 12232
rect 20364 12220 20392 12384
rect 21634 12316 21640 12368
rect 21692 12356 21698 12368
rect 21692 12328 23060 12356
rect 21692 12316 21698 12328
rect 20717 12291 20775 12297
rect 20717 12257 20729 12291
rect 20763 12288 20775 12291
rect 20806 12288 20812 12300
rect 20763 12260 20812 12288
rect 20763 12257 20775 12260
rect 20717 12251 20775 12257
rect 20806 12248 20812 12260
rect 20864 12248 20870 12300
rect 21266 12248 21272 12300
rect 21324 12248 21330 12300
rect 21726 12248 21732 12300
rect 21784 12288 21790 12300
rect 23032 12297 23060 12328
rect 22750 12291 22808 12297
rect 22750 12288 22762 12291
rect 21784 12260 22762 12288
rect 21784 12248 21790 12260
rect 22750 12257 22762 12260
rect 22796 12257 22808 12291
rect 22750 12251 22808 12257
rect 23017 12291 23075 12297
rect 23017 12257 23029 12291
rect 23063 12257 23075 12291
rect 23017 12251 23075 12257
rect 20312 12192 20392 12220
rect 20312 12180 20318 12192
rect 20438 12180 20444 12232
rect 20496 12220 20502 12232
rect 20533 12223 20591 12229
rect 20533 12220 20545 12223
rect 20496 12192 20545 12220
rect 20496 12180 20502 12192
rect 20533 12189 20545 12192
rect 20579 12189 20591 12223
rect 20533 12183 20591 12189
rect 19518 12152 19524 12164
rect 16960 12124 19524 12152
rect 16853 12115 16911 12121
rect 19518 12112 19524 12124
rect 19576 12112 19582 12164
rect 20548 12152 20576 12183
rect 20622 12180 20628 12232
rect 20680 12180 20686 12232
rect 21818 12152 21824 12164
rect 20548 12124 21824 12152
rect 21818 12112 21824 12124
rect 21876 12112 21882 12164
rect 15068 12056 15148 12084
rect 15068 12044 15074 12056
rect 15470 12044 15476 12096
rect 15528 12084 15534 12096
rect 15841 12087 15899 12093
rect 15841 12084 15853 12087
rect 15528 12056 15853 12084
rect 15528 12044 15534 12056
rect 15841 12053 15853 12056
rect 15887 12053 15899 12087
rect 15841 12047 15899 12053
rect 16022 12044 16028 12096
rect 16080 12084 16086 12096
rect 16117 12087 16175 12093
rect 16117 12084 16129 12087
rect 16080 12056 16129 12084
rect 16080 12044 16086 12056
rect 16117 12053 16129 12056
rect 16163 12053 16175 12087
rect 16117 12047 16175 12053
rect 16390 12044 16396 12096
rect 16448 12084 16454 12096
rect 17310 12084 17316 12096
rect 16448 12056 17316 12084
rect 16448 12044 16454 12056
rect 17310 12044 17316 12056
rect 17368 12084 17374 12096
rect 17770 12084 17776 12096
rect 17368 12056 17776 12084
rect 17368 12044 17374 12056
rect 17770 12044 17776 12056
rect 17828 12044 17834 12096
rect 17957 12087 18015 12093
rect 17957 12053 17969 12087
rect 18003 12084 18015 12087
rect 18138 12084 18144 12096
rect 18003 12056 18144 12084
rect 18003 12053 18015 12056
rect 17957 12047 18015 12053
rect 18138 12044 18144 12056
rect 18196 12044 18202 12096
rect 18782 12044 18788 12096
rect 18840 12044 18846 12096
rect 18874 12044 18880 12096
rect 18932 12084 18938 12096
rect 19061 12087 19119 12093
rect 19061 12084 19073 12087
rect 18932 12056 19073 12084
rect 18932 12044 18938 12056
rect 19061 12053 19073 12056
rect 19107 12053 19119 12087
rect 19061 12047 19119 12053
rect 21085 12087 21143 12093
rect 21085 12053 21097 12087
rect 21131 12084 21143 12087
rect 21450 12084 21456 12096
rect 21131 12056 21456 12084
rect 21131 12053 21143 12056
rect 21085 12047 21143 12053
rect 21450 12044 21456 12056
rect 21508 12044 21514 12096
rect 21542 12044 21548 12096
rect 21600 12084 21606 12096
rect 21637 12087 21695 12093
rect 21637 12084 21649 12087
rect 21600 12056 21649 12084
rect 21600 12044 21606 12056
rect 21637 12053 21649 12056
rect 21683 12053 21695 12087
rect 21637 12047 21695 12053
rect 552 11994 23368 12016
rect 552 11942 1366 11994
rect 1418 11942 1430 11994
rect 1482 11942 1494 11994
rect 1546 11942 1558 11994
rect 1610 11942 1622 11994
rect 1674 11942 1686 11994
rect 1738 11942 7366 11994
rect 7418 11942 7430 11994
rect 7482 11942 7494 11994
rect 7546 11942 7558 11994
rect 7610 11942 7622 11994
rect 7674 11942 7686 11994
rect 7738 11942 13366 11994
rect 13418 11942 13430 11994
rect 13482 11942 13494 11994
rect 13546 11942 13558 11994
rect 13610 11942 13622 11994
rect 13674 11942 13686 11994
rect 13738 11942 19366 11994
rect 19418 11942 19430 11994
rect 19482 11942 19494 11994
rect 19546 11942 19558 11994
rect 19610 11942 19622 11994
rect 19674 11942 19686 11994
rect 19738 11942 23368 11994
rect 552 11920 23368 11942
rect 1121 11883 1179 11889
rect 1121 11849 1133 11883
rect 1167 11880 1179 11883
rect 2409 11883 2467 11889
rect 2409 11880 2421 11883
rect 1167 11852 2421 11880
rect 1167 11849 1179 11852
rect 1121 11843 1179 11849
rect 2409 11849 2421 11852
rect 2455 11849 2467 11883
rect 2409 11843 2467 11849
rect 3712 11852 4292 11880
rect 934 11772 940 11824
rect 992 11812 998 11824
rect 1302 11812 1308 11824
rect 992 11784 1308 11812
rect 992 11772 998 11784
rect 1302 11772 1308 11784
rect 1360 11772 1366 11824
rect 1118 11704 1124 11756
rect 1176 11744 1182 11756
rect 1397 11747 1455 11753
rect 1397 11744 1409 11747
rect 1176 11716 1409 11744
rect 1176 11704 1182 11716
rect 1397 11713 1409 11716
rect 1443 11713 1455 11747
rect 1397 11707 1455 11713
rect 1578 11704 1584 11756
rect 1636 11704 1642 11756
rect 1670 11704 1676 11756
rect 1728 11704 1734 11756
rect 1765 11747 1823 11753
rect 1765 11713 1777 11747
rect 1811 11713 1823 11747
rect 1946 11744 1952 11756
rect 1765 11707 1823 11713
rect 1872 11716 1952 11744
rect 750 11636 756 11688
rect 808 11676 814 11688
rect 1780 11676 1808 11707
rect 1872 11685 1900 11716
rect 1946 11704 1952 11716
rect 2004 11704 2010 11756
rect 2884 11716 3556 11744
rect 808 11648 1808 11676
rect 1857 11679 1915 11685
rect 808 11636 814 11648
rect 842 11568 848 11620
rect 900 11608 906 11620
rect 1118 11617 1124 11620
rect 1105 11611 1124 11617
rect 900 11580 1072 11608
rect 900 11568 906 11580
rect 934 11500 940 11552
rect 992 11500 998 11552
rect 1044 11540 1072 11580
rect 1105 11577 1117 11611
rect 1105 11571 1124 11577
rect 1118 11568 1124 11571
rect 1176 11568 1182 11620
rect 1302 11568 1308 11620
rect 1360 11568 1366 11620
rect 1688 11608 1716 11648
rect 1857 11645 1869 11679
rect 1903 11645 1915 11679
rect 2225 11679 2283 11685
rect 2225 11676 2237 11679
rect 1857 11639 1915 11645
rect 1964 11648 2237 11676
rect 1762 11608 1768 11620
rect 1688 11580 1768 11608
rect 1762 11568 1768 11580
rect 1820 11608 1826 11620
rect 1964 11608 1992 11648
rect 2225 11645 2237 11648
rect 2271 11645 2283 11679
rect 2225 11639 2283 11645
rect 2774 11636 2780 11688
rect 2832 11636 2838 11688
rect 2884 11685 2912 11716
rect 2869 11679 2927 11685
rect 2869 11645 2881 11679
rect 2915 11645 2927 11679
rect 2869 11639 2927 11645
rect 3053 11679 3111 11685
rect 3053 11645 3065 11679
rect 3099 11676 3111 11679
rect 3418 11676 3424 11688
rect 3099 11648 3424 11676
rect 3099 11645 3111 11648
rect 3053 11639 3111 11645
rect 3418 11636 3424 11648
rect 3476 11636 3482 11688
rect 1820 11580 1992 11608
rect 2041 11611 2099 11617
rect 1820 11568 1826 11580
rect 2041 11577 2053 11611
rect 2087 11577 2099 11611
rect 3237 11611 3295 11617
rect 3237 11608 3249 11611
rect 2041 11571 2099 11577
rect 2746 11580 3249 11608
rect 1946 11540 1952 11552
rect 1044 11512 1952 11540
rect 1946 11500 1952 11512
rect 2004 11540 2010 11552
rect 2056 11540 2084 11571
rect 2746 11552 2774 11580
rect 3237 11577 3249 11580
rect 3283 11577 3295 11611
rect 3237 11571 3295 11577
rect 2004 11512 2084 11540
rect 2004 11500 2010 11512
rect 2682 11500 2688 11552
rect 2740 11512 2774 11552
rect 3528 11540 3556 11716
rect 3712 11685 3740 11852
rect 4264 11756 4292 11852
rect 5074 11840 5080 11892
rect 5132 11840 5138 11892
rect 5350 11840 5356 11892
rect 5408 11880 5414 11892
rect 9766 11880 9772 11892
rect 5408 11852 9772 11880
rect 5408 11840 5414 11852
rect 9766 11840 9772 11852
rect 9824 11840 9830 11892
rect 9858 11840 9864 11892
rect 9916 11880 9922 11892
rect 10045 11883 10103 11889
rect 10045 11880 10057 11883
rect 9916 11852 10057 11880
rect 9916 11840 9922 11852
rect 10045 11849 10057 11852
rect 10091 11849 10103 11883
rect 12158 11880 12164 11892
rect 10045 11843 10103 11849
rect 10152 11852 12164 11880
rect 8754 11772 8760 11824
rect 8812 11812 8818 11824
rect 10152 11812 10180 11852
rect 12158 11840 12164 11852
rect 12216 11840 12222 11892
rect 14274 11840 14280 11892
rect 14332 11880 14338 11892
rect 16298 11880 16304 11892
rect 14332 11852 16304 11880
rect 14332 11840 14338 11852
rect 16298 11840 16304 11852
rect 16356 11840 16362 11892
rect 16850 11840 16856 11892
rect 16908 11840 16914 11892
rect 16942 11840 16948 11892
rect 17000 11840 17006 11892
rect 17586 11840 17592 11892
rect 17644 11840 17650 11892
rect 18782 11840 18788 11892
rect 18840 11840 18846 11892
rect 19521 11883 19579 11889
rect 19521 11849 19533 11883
rect 19567 11880 19579 11883
rect 19886 11880 19892 11892
rect 19567 11852 19892 11880
rect 19567 11849 19579 11852
rect 19521 11843 19579 11849
rect 19886 11840 19892 11852
rect 19944 11840 19950 11892
rect 19978 11840 19984 11892
rect 20036 11840 20042 11892
rect 20070 11840 20076 11892
rect 20128 11840 20134 11892
rect 21637 11883 21695 11889
rect 21637 11849 21649 11883
rect 21683 11880 21695 11883
rect 21726 11880 21732 11892
rect 21683 11852 21732 11880
rect 21683 11849 21695 11852
rect 21637 11843 21695 11849
rect 21726 11840 21732 11852
rect 21784 11840 21790 11892
rect 12434 11812 12440 11824
rect 8812 11784 8984 11812
rect 8812 11772 8818 11784
rect 3786 11704 3792 11756
rect 3844 11744 3850 11756
rect 3844 11716 4016 11744
rect 3844 11704 3850 11716
rect 3697 11679 3755 11685
rect 3697 11645 3709 11679
rect 3743 11645 3755 11679
rect 3697 11639 3755 11645
rect 3881 11679 3939 11685
rect 3881 11645 3893 11679
rect 3927 11645 3939 11679
rect 3988 11676 4016 11716
rect 4246 11704 4252 11756
rect 4304 11704 4310 11756
rect 4338 11704 4344 11756
rect 4396 11744 4402 11756
rect 4982 11744 4988 11756
rect 4396 11716 4988 11744
rect 4396 11704 4402 11716
rect 4982 11704 4988 11716
rect 5040 11744 5046 11756
rect 8846 11744 8852 11756
rect 5040 11716 5488 11744
rect 5040 11704 5046 11716
rect 4157 11679 4215 11685
rect 4157 11676 4169 11679
rect 3988 11648 4169 11676
rect 3881 11639 3939 11645
rect 4157 11645 4169 11648
rect 4203 11645 4215 11679
rect 4157 11639 4215 11645
rect 4801 11679 4859 11685
rect 4801 11645 4813 11679
rect 4847 11676 4859 11679
rect 4890 11676 4896 11688
rect 4847 11648 4896 11676
rect 4847 11645 4859 11648
rect 4801 11639 4859 11645
rect 3602 11568 3608 11620
rect 3660 11608 3666 11620
rect 3896 11608 3924 11639
rect 4890 11636 4896 11648
rect 4948 11636 4954 11688
rect 5460 11685 5488 11716
rect 7576 11716 8852 11744
rect 5445 11679 5503 11685
rect 5445 11645 5457 11679
rect 5491 11645 5503 11679
rect 5445 11639 5503 11645
rect 6086 11636 6092 11688
rect 6144 11676 6150 11688
rect 7282 11676 7288 11688
rect 6144 11648 7288 11676
rect 6144 11636 6150 11648
rect 7282 11636 7288 11648
rect 7340 11636 7346 11688
rect 3660 11580 3924 11608
rect 5261 11611 5319 11617
rect 3660 11568 3666 11580
rect 5261 11577 5273 11611
rect 5307 11608 5319 11611
rect 5350 11608 5356 11620
rect 5307 11580 5356 11608
rect 5307 11577 5319 11580
rect 5261 11571 5319 11577
rect 5350 11568 5356 11580
rect 5408 11608 5414 11620
rect 7576 11608 7604 11716
rect 8846 11704 8852 11716
rect 8904 11704 8910 11756
rect 8956 11753 8984 11784
rect 9048 11784 10180 11812
rect 11900 11784 12440 11812
rect 8941 11747 8999 11753
rect 8941 11713 8953 11747
rect 8987 11713 8999 11747
rect 8941 11707 8999 11713
rect 8478 11636 8484 11688
rect 8536 11676 8542 11688
rect 8573 11679 8631 11685
rect 8573 11676 8585 11679
rect 8536 11648 8585 11676
rect 8536 11636 8542 11648
rect 8573 11645 8585 11648
rect 8619 11645 8631 11679
rect 8573 11639 8631 11645
rect 8754 11636 8760 11688
rect 8812 11676 8818 11688
rect 9048 11685 9076 11784
rect 9401 11747 9459 11753
rect 9401 11713 9413 11747
rect 9447 11713 9459 11747
rect 9953 11747 10011 11753
rect 9953 11744 9965 11747
rect 9401 11707 9459 11713
rect 9692 11716 9965 11744
rect 9033 11679 9091 11685
rect 9033 11676 9045 11679
rect 8812 11648 9045 11676
rect 8812 11636 8818 11648
rect 9033 11645 9045 11648
rect 9079 11645 9091 11679
rect 9416 11676 9444 11707
rect 9692 11685 9720 11716
rect 9953 11713 9965 11716
rect 9999 11713 10011 11747
rect 9953 11707 10011 11713
rect 11422 11704 11428 11756
rect 11480 11704 11486 11756
rect 11514 11704 11520 11756
rect 11572 11704 11578 11756
rect 11900 11753 11928 11784
rect 12434 11772 12440 11784
rect 12492 11812 12498 11824
rect 12894 11812 12900 11824
rect 12492 11784 12900 11812
rect 12492 11772 12498 11784
rect 12894 11772 12900 11784
rect 12952 11772 12958 11824
rect 13722 11772 13728 11824
rect 13780 11812 13786 11824
rect 13780 11784 15884 11812
rect 13780 11772 13786 11784
rect 11885 11747 11943 11753
rect 11885 11713 11897 11747
rect 11931 11713 11943 11747
rect 11885 11707 11943 11713
rect 12161 11747 12219 11753
rect 12161 11713 12173 11747
rect 12207 11744 12219 11747
rect 12207 11716 12480 11744
rect 12207 11713 12219 11716
rect 12161 11707 12219 11713
rect 9677 11679 9735 11685
rect 9677 11676 9689 11679
rect 9416 11648 9689 11676
rect 9033 11639 9091 11645
rect 9677 11645 9689 11648
rect 9723 11645 9735 11679
rect 9677 11639 9735 11645
rect 9858 11636 9864 11688
rect 9916 11636 9922 11688
rect 10229 11679 10287 11685
rect 10229 11645 10241 11679
rect 10275 11645 10287 11679
rect 10229 11639 10287 11645
rect 10413 11679 10471 11685
rect 10413 11645 10425 11679
rect 10459 11676 10471 11679
rect 10505 11679 10563 11685
rect 10505 11676 10517 11679
rect 10459 11648 10517 11676
rect 10459 11645 10471 11648
rect 10413 11639 10471 11645
rect 10505 11645 10517 11648
rect 10551 11645 10563 11679
rect 10505 11639 10563 11645
rect 10781 11679 10839 11685
rect 10781 11645 10793 11679
rect 10827 11676 10839 11679
rect 11146 11676 11152 11688
rect 10827 11648 11152 11676
rect 10827 11645 10839 11648
rect 10781 11639 10839 11645
rect 5408 11580 7604 11608
rect 5408 11568 5414 11580
rect 7650 11568 7656 11620
rect 7708 11608 7714 11620
rect 10244 11608 10272 11639
rect 11146 11636 11152 11648
rect 11204 11636 11210 11688
rect 11241 11679 11299 11685
rect 11241 11645 11253 11679
rect 11287 11676 11299 11679
rect 11330 11676 11336 11688
rect 11287 11648 11336 11676
rect 11287 11645 11299 11648
rect 11241 11639 11299 11645
rect 11330 11636 11336 11648
rect 11388 11636 11394 11688
rect 11790 11636 11796 11688
rect 11848 11636 11854 11688
rect 12342 11608 12348 11620
rect 7708 11580 12348 11608
rect 7708 11568 7714 11580
rect 12342 11568 12348 11580
rect 12400 11568 12406 11620
rect 12452 11608 12480 11716
rect 13078 11704 13084 11756
rect 13136 11744 13142 11756
rect 13136 11716 13768 11744
rect 13136 11704 13142 11716
rect 12986 11636 12992 11688
rect 13044 11636 13050 11688
rect 13262 11636 13268 11688
rect 13320 11636 13326 11688
rect 13740 11685 13768 11716
rect 13832 11716 14320 11744
rect 13832 11688 13860 11716
rect 13725 11679 13783 11685
rect 13725 11645 13737 11679
rect 13771 11645 13783 11679
rect 13725 11639 13783 11645
rect 13078 11608 13084 11620
rect 12452 11580 13084 11608
rect 13078 11568 13084 11580
rect 13136 11568 13142 11620
rect 13740 11608 13768 11639
rect 13814 11636 13820 11688
rect 13872 11636 13878 11688
rect 14001 11679 14059 11685
rect 14001 11645 14013 11679
rect 14047 11676 14059 11679
rect 14182 11676 14188 11688
rect 14047 11648 14188 11676
rect 14047 11645 14059 11648
rect 14001 11639 14059 11645
rect 14182 11636 14188 11648
rect 14240 11636 14246 11688
rect 14292 11685 14320 11716
rect 14366 11704 14372 11756
rect 14424 11744 14430 11756
rect 14424 11716 14596 11744
rect 14424 11704 14430 11716
rect 14277 11679 14335 11685
rect 14277 11645 14289 11679
rect 14323 11645 14335 11679
rect 14277 11639 14335 11645
rect 14461 11679 14519 11685
rect 14461 11645 14473 11679
rect 14507 11645 14519 11679
rect 14461 11639 14519 11645
rect 14476 11608 14504 11639
rect 13740 11580 14504 11608
rect 14568 11608 14596 11716
rect 15010 11704 15016 11756
rect 15068 11744 15074 11756
rect 15068 11716 15148 11744
rect 15068 11704 15074 11716
rect 14826 11636 14832 11688
rect 14884 11676 14890 11688
rect 15120 11685 15148 11716
rect 15194 11704 15200 11756
rect 15252 11744 15258 11756
rect 15381 11747 15439 11753
rect 15381 11744 15393 11747
rect 15252 11716 15393 11744
rect 15252 11704 15258 11716
rect 15381 11713 15393 11716
rect 15427 11713 15439 11747
rect 15381 11707 15439 11713
rect 15470 11704 15476 11756
rect 15528 11704 15534 11756
rect 15562 11704 15568 11756
rect 15620 11704 15626 11756
rect 15856 11744 15884 11784
rect 15930 11772 15936 11824
rect 15988 11812 15994 11824
rect 17957 11815 18015 11821
rect 15988 11784 17908 11812
rect 15988 11772 15994 11784
rect 15856 11716 17448 11744
rect 14921 11679 14979 11685
rect 14921 11676 14933 11679
rect 14884 11648 14933 11676
rect 14884 11636 14890 11648
rect 14921 11645 14933 11648
rect 14967 11645 14979 11679
rect 14921 11639 14979 11645
rect 15105 11679 15163 11685
rect 15105 11645 15117 11679
rect 15151 11645 15163 11679
rect 15105 11639 15163 11645
rect 15289 11679 15347 11685
rect 15289 11645 15301 11679
rect 15335 11676 15347 11679
rect 15746 11676 15752 11688
rect 15335 11648 15752 11676
rect 15335 11645 15347 11648
rect 15289 11639 15347 11645
rect 15746 11636 15752 11648
rect 15804 11636 15810 11688
rect 16574 11636 16580 11688
rect 16632 11636 16638 11688
rect 16666 11636 16672 11688
rect 16724 11636 16730 11688
rect 16868 11685 16896 11716
rect 16853 11679 16911 11685
rect 16853 11645 16865 11679
rect 16899 11645 16911 11679
rect 16853 11639 16911 11645
rect 17126 11636 17132 11688
rect 17184 11636 17190 11688
rect 17420 11685 17448 11716
rect 17494 11704 17500 11756
rect 17552 11704 17558 11756
rect 17681 11747 17739 11753
rect 17681 11713 17693 11747
rect 17727 11744 17739 11747
rect 17770 11744 17776 11756
rect 17727 11716 17776 11744
rect 17727 11713 17739 11716
rect 17681 11707 17739 11713
rect 17770 11704 17776 11716
rect 17828 11704 17834 11756
rect 17880 11744 17908 11784
rect 17957 11781 17969 11815
rect 18003 11812 18015 11815
rect 19153 11815 19211 11821
rect 19153 11812 19165 11815
rect 18003 11784 19165 11812
rect 18003 11781 18015 11784
rect 17957 11775 18015 11781
rect 19153 11781 19165 11784
rect 19199 11781 19211 11815
rect 19996 11812 20024 11840
rect 20165 11815 20223 11821
rect 20165 11812 20177 11815
rect 19996 11784 20177 11812
rect 19153 11775 19211 11781
rect 20165 11781 20177 11784
rect 20211 11781 20223 11815
rect 21082 11812 21088 11824
rect 20165 11775 20223 11781
rect 20272 11784 21088 11812
rect 17880 11716 17984 11744
rect 17405 11679 17463 11685
rect 17405 11645 17417 11679
rect 17451 11645 17463 11679
rect 17512 11676 17540 11704
rect 17865 11679 17923 11685
rect 17865 11676 17877 11679
rect 17512 11648 17877 11676
rect 17405 11639 17463 11645
rect 17865 11645 17877 11648
rect 17911 11645 17923 11679
rect 17956 11676 17984 11716
rect 18138 11704 18144 11756
rect 18196 11744 18202 11756
rect 18693 11747 18751 11753
rect 18693 11744 18705 11747
rect 18196 11716 18705 11744
rect 18196 11704 18202 11716
rect 18693 11713 18705 11716
rect 18739 11713 18751 11747
rect 18874 11744 18880 11756
rect 18693 11707 18751 11713
rect 18800 11716 18880 11744
rect 18233 11679 18291 11685
rect 17956 11648 18184 11676
rect 17865 11639 17923 11645
rect 15013 11611 15071 11617
rect 14568 11580 14872 11608
rect 14844 11552 14872 11580
rect 15013 11577 15025 11611
rect 15059 11608 15071 11611
rect 15470 11608 15476 11620
rect 15059 11580 15476 11608
rect 15059 11577 15071 11580
rect 15013 11571 15071 11577
rect 15470 11568 15476 11580
rect 15528 11568 15534 11620
rect 16684 11608 16712 11636
rect 16942 11608 16948 11620
rect 16684 11580 16948 11608
rect 16942 11568 16948 11580
rect 17000 11568 17006 11620
rect 17420 11608 17448 11639
rect 17773 11611 17831 11617
rect 17420 11580 17724 11608
rect 3970 11540 3976 11552
rect 3528 11512 3976 11540
rect 2740 11500 2746 11512
rect 3970 11500 3976 11512
rect 4028 11500 4034 11552
rect 4246 11500 4252 11552
rect 4304 11540 4310 11552
rect 4525 11543 4583 11549
rect 4525 11540 4537 11543
rect 4304 11512 4537 11540
rect 4304 11500 4310 11512
rect 4525 11509 4537 11512
rect 4571 11509 4583 11543
rect 4525 11503 4583 11509
rect 4617 11543 4675 11549
rect 4617 11509 4629 11543
rect 4663 11540 4675 11543
rect 4982 11540 4988 11552
rect 4663 11512 4988 11540
rect 4663 11509 4675 11512
rect 4617 11503 4675 11509
rect 4982 11500 4988 11512
rect 5040 11500 5046 11552
rect 5074 11500 5080 11552
rect 5132 11540 5138 11552
rect 5534 11540 5540 11552
rect 5132 11512 5540 11540
rect 5132 11500 5138 11512
rect 5534 11500 5540 11512
rect 5592 11500 5598 11552
rect 5810 11500 5816 11552
rect 5868 11540 5874 11552
rect 8389 11543 8447 11549
rect 8389 11540 8401 11543
rect 5868 11512 8401 11540
rect 5868 11500 5874 11512
rect 8389 11509 8401 11512
rect 8435 11540 8447 11543
rect 9582 11540 9588 11552
rect 8435 11512 9588 11540
rect 8435 11509 8447 11512
rect 8389 11503 8447 11509
rect 9582 11500 9588 11512
rect 9640 11500 9646 11552
rect 9769 11543 9827 11549
rect 9769 11509 9781 11543
rect 9815 11540 9827 11543
rect 10597 11543 10655 11549
rect 10597 11540 10609 11543
rect 9815 11512 10609 11540
rect 9815 11509 9827 11512
rect 9769 11503 9827 11509
rect 10597 11509 10609 11512
rect 10643 11509 10655 11543
rect 10597 11503 10655 11509
rect 10962 11500 10968 11552
rect 11020 11500 11026 11552
rect 11054 11500 11060 11552
rect 11112 11500 11118 11552
rect 12802 11500 12808 11552
rect 12860 11500 12866 11552
rect 13173 11543 13231 11549
rect 13173 11509 13185 11543
rect 13219 11540 13231 11543
rect 14090 11540 14096 11552
rect 13219 11512 14096 11540
rect 13219 11509 13231 11512
rect 13173 11503 13231 11509
rect 14090 11500 14096 11512
rect 14148 11500 14154 11552
rect 14182 11500 14188 11552
rect 14240 11500 14246 11552
rect 14369 11543 14427 11549
rect 14369 11509 14381 11543
rect 14415 11540 14427 11543
rect 14458 11540 14464 11552
rect 14415 11512 14464 11540
rect 14415 11509 14427 11512
rect 14369 11503 14427 11509
rect 14458 11500 14464 11512
rect 14516 11500 14522 11552
rect 14826 11500 14832 11552
rect 14884 11500 14890 11552
rect 15562 11500 15568 11552
rect 15620 11540 15626 11552
rect 15749 11543 15807 11549
rect 15749 11540 15761 11543
rect 15620 11512 15761 11540
rect 15620 11500 15626 11512
rect 15749 11509 15761 11512
rect 15795 11509 15807 11543
rect 15749 11503 15807 11509
rect 17221 11543 17279 11549
rect 17221 11509 17233 11543
rect 17267 11540 17279 11543
rect 17402 11540 17408 11552
rect 17267 11512 17408 11540
rect 17267 11509 17279 11512
rect 17221 11503 17279 11509
rect 17402 11500 17408 11512
rect 17460 11500 17466 11552
rect 17696 11540 17724 11580
rect 17773 11577 17785 11611
rect 17819 11608 17831 11611
rect 18046 11608 18052 11620
rect 17819 11580 18052 11608
rect 17819 11577 17831 11580
rect 17773 11571 17831 11577
rect 18046 11568 18052 11580
rect 18104 11568 18110 11620
rect 18156 11617 18184 11648
rect 18233 11645 18245 11679
rect 18279 11676 18291 11679
rect 18800 11676 18828 11716
rect 18874 11704 18880 11716
rect 18932 11704 18938 11756
rect 19334 11704 19340 11756
rect 19392 11704 19398 11756
rect 19426 11704 19432 11756
rect 19484 11744 19490 11756
rect 19886 11744 19892 11756
rect 19484 11716 19892 11744
rect 19484 11704 19490 11716
rect 19886 11704 19892 11716
rect 19944 11744 19950 11756
rect 19981 11747 20039 11753
rect 19981 11744 19993 11747
rect 19944 11716 19993 11744
rect 19944 11704 19950 11716
rect 19981 11713 19993 11716
rect 20027 11713 20039 11747
rect 20272 11744 20300 11784
rect 21082 11772 21088 11784
rect 21140 11772 21146 11824
rect 20622 11744 20628 11756
rect 19981 11707 20039 11713
rect 20088 11716 20300 11744
rect 20548 11716 20628 11744
rect 18279 11648 18828 11676
rect 18969 11679 19027 11685
rect 18279 11645 18291 11648
rect 18233 11639 18291 11645
rect 18969 11645 18981 11679
rect 19015 11645 19027 11679
rect 18969 11639 19027 11645
rect 18141 11611 18199 11617
rect 18141 11577 18153 11611
rect 18187 11608 18199 11611
rect 18690 11608 18696 11620
rect 18187 11580 18696 11608
rect 18187 11577 18199 11580
rect 18141 11571 18199 11577
rect 18690 11568 18696 11580
rect 18748 11568 18754 11620
rect 18984 11540 19012 11639
rect 19058 11636 19064 11688
rect 19116 11676 19122 11688
rect 19242 11676 19248 11688
rect 19116 11648 19248 11676
rect 19116 11636 19122 11648
rect 19242 11636 19248 11648
rect 19300 11636 19306 11688
rect 19613 11679 19671 11685
rect 19613 11645 19625 11679
rect 19659 11676 19671 11679
rect 20088 11676 20116 11716
rect 20162 11676 20168 11688
rect 19659 11648 20168 11676
rect 19659 11645 19671 11648
rect 19613 11639 19671 11645
rect 20162 11636 20168 11648
rect 20220 11636 20226 11688
rect 20254 11636 20260 11688
rect 20312 11636 20318 11688
rect 19337 11611 19395 11617
rect 19337 11608 19349 11611
rect 19076 11580 19349 11608
rect 19076 11552 19104 11580
rect 19337 11577 19349 11580
rect 19383 11577 19395 11611
rect 19337 11571 19395 11577
rect 19978 11568 19984 11620
rect 20036 11608 20042 11620
rect 20272 11608 20300 11636
rect 20036 11580 20300 11608
rect 20036 11568 20042 11580
rect 17696 11512 19012 11540
rect 19058 11500 19064 11552
rect 19116 11500 19122 11552
rect 20254 11500 20260 11552
rect 20312 11540 20318 11552
rect 20548 11540 20576 11716
rect 20622 11704 20628 11716
rect 20680 11704 20686 11756
rect 21542 11744 21548 11756
rect 21376 11716 21548 11744
rect 20898 11636 20904 11688
rect 20956 11636 20962 11688
rect 21376 11685 21404 11716
rect 21542 11704 21548 11716
rect 21600 11744 21606 11756
rect 21600 11716 22232 11744
rect 21600 11704 21606 11716
rect 21361 11679 21419 11685
rect 21361 11645 21373 11679
rect 21407 11645 21419 11679
rect 21361 11639 21419 11645
rect 21450 11636 21456 11688
rect 21508 11636 21514 11688
rect 21913 11679 21971 11685
rect 21913 11645 21925 11679
rect 21959 11676 21971 11679
rect 22094 11676 22100 11688
rect 21959 11648 22100 11676
rect 21959 11645 21971 11648
rect 21913 11639 21971 11645
rect 22094 11636 22100 11648
rect 22152 11636 22158 11688
rect 22204 11685 22232 11716
rect 22189 11679 22247 11685
rect 22189 11645 22201 11679
rect 22235 11645 22247 11679
rect 22189 11639 22247 11645
rect 22278 11636 22284 11688
rect 22336 11676 22342 11688
rect 22465 11679 22523 11685
rect 22465 11676 22477 11679
rect 22336 11648 22477 11676
rect 22336 11636 22342 11648
rect 22465 11645 22477 11648
rect 22511 11645 22523 11679
rect 22465 11639 22523 11645
rect 20622 11568 20628 11620
rect 20680 11608 20686 11620
rect 21269 11611 21327 11617
rect 21269 11608 21281 11611
rect 20680 11580 21281 11608
rect 20680 11568 20686 11580
rect 21269 11577 21281 11580
rect 21315 11577 21327 11611
rect 21269 11571 21327 11577
rect 21542 11568 21548 11620
rect 21600 11608 21606 11620
rect 21600 11580 22048 11608
rect 21600 11568 21606 11580
rect 20312 11512 20576 11540
rect 20312 11500 20318 11512
rect 20714 11500 20720 11552
rect 20772 11500 20778 11552
rect 21726 11500 21732 11552
rect 21784 11500 21790 11552
rect 22020 11549 22048 11580
rect 22005 11543 22063 11549
rect 22005 11509 22017 11543
rect 22051 11509 22063 11543
rect 22005 11503 22063 11509
rect 22186 11500 22192 11552
rect 22244 11540 22250 11552
rect 22281 11543 22339 11549
rect 22281 11540 22293 11543
rect 22244 11512 22293 11540
rect 22244 11500 22250 11512
rect 22281 11509 22293 11512
rect 22327 11509 22339 11543
rect 22281 11503 22339 11509
rect 552 11450 23368 11472
rect 552 11398 4366 11450
rect 4418 11398 4430 11450
rect 4482 11398 4494 11450
rect 4546 11398 4558 11450
rect 4610 11398 4622 11450
rect 4674 11398 4686 11450
rect 4738 11398 10366 11450
rect 10418 11398 10430 11450
rect 10482 11398 10494 11450
rect 10546 11398 10558 11450
rect 10610 11398 10622 11450
rect 10674 11398 10686 11450
rect 10738 11398 16366 11450
rect 16418 11398 16430 11450
rect 16482 11398 16494 11450
rect 16546 11398 16558 11450
rect 16610 11398 16622 11450
rect 16674 11398 16686 11450
rect 16738 11398 22366 11450
rect 22418 11398 22430 11450
rect 22482 11398 22494 11450
rect 22546 11398 22558 11450
rect 22610 11398 22622 11450
rect 22674 11398 22686 11450
rect 22738 11398 23368 11450
rect 552 11376 23368 11398
rect 1670 11296 1676 11348
rect 1728 11336 1734 11348
rect 2314 11336 2320 11348
rect 1728 11308 2320 11336
rect 1728 11296 1734 11308
rect 2314 11296 2320 11308
rect 2372 11296 2378 11348
rect 2777 11339 2835 11345
rect 2777 11305 2789 11339
rect 2823 11336 2835 11339
rect 2958 11336 2964 11348
rect 2823 11308 2964 11336
rect 2823 11305 2835 11308
rect 2777 11299 2835 11305
rect 2958 11296 2964 11308
rect 3016 11336 3022 11348
rect 3694 11336 3700 11348
rect 3016 11308 3700 11336
rect 3016 11296 3022 11308
rect 3694 11296 3700 11308
rect 3752 11296 3758 11348
rect 4525 11339 4583 11345
rect 4525 11305 4537 11339
rect 4571 11336 4583 11339
rect 4890 11336 4896 11348
rect 4571 11308 4896 11336
rect 4571 11305 4583 11308
rect 4525 11299 4583 11305
rect 3418 11268 3424 11280
rect 3068 11240 3424 11268
rect 1118 11200 1124 11212
rect 1044 11172 1124 11200
rect 842 11092 848 11144
rect 900 11132 906 11144
rect 1044 11141 1072 11172
rect 1118 11160 1124 11172
rect 1176 11160 1182 11212
rect 1302 11209 1308 11212
rect 1296 11163 1308 11209
rect 1302 11160 1308 11163
rect 1360 11160 1366 11212
rect 2593 11203 2651 11209
rect 2593 11169 2605 11203
rect 2639 11200 2651 11203
rect 2774 11200 2780 11212
rect 2639 11172 2780 11200
rect 2639 11169 2651 11172
rect 2593 11163 2651 11169
rect 2774 11160 2780 11172
rect 2832 11160 2838 11212
rect 3068 11209 3096 11240
rect 3418 11228 3424 11240
rect 3476 11268 3482 11280
rect 3881 11271 3939 11277
rect 3881 11268 3893 11271
rect 3476 11240 3893 11268
rect 3476 11228 3482 11240
rect 3881 11237 3893 11240
rect 3927 11237 3939 11271
rect 3881 11231 3939 11237
rect 3053 11203 3111 11209
rect 3053 11169 3065 11203
rect 3099 11169 3111 11203
rect 3053 11163 3111 11169
rect 3237 11203 3295 11209
rect 3237 11169 3249 11203
rect 3283 11169 3295 11203
rect 3237 11163 3295 11169
rect 1029 11135 1087 11141
rect 1029 11132 1041 11135
rect 900 11104 1041 11132
rect 900 11092 906 11104
rect 1029 11101 1041 11104
rect 1075 11101 1087 11135
rect 1029 11095 1087 11101
rect 2869 11135 2927 11141
rect 2869 11101 2881 11135
rect 2915 11132 2927 11135
rect 3142 11132 3148 11144
rect 2915 11104 3148 11132
rect 2915 11101 2927 11104
rect 2869 11095 2927 11101
rect 3142 11092 3148 11104
rect 3200 11092 3206 11144
rect 2406 10956 2412 11008
rect 2464 10956 2470 11008
rect 3142 10956 3148 11008
rect 3200 10996 3206 11008
rect 3252 10996 3280 11163
rect 3326 11160 3332 11212
rect 3384 11160 3390 11212
rect 3605 11203 3663 11209
rect 3605 11169 3617 11203
rect 3651 11200 3663 11203
rect 3694 11200 3700 11212
rect 3651 11172 3700 11200
rect 3651 11169 3663 11172
rect 3605 11163 3663 11169
rect 3694 11160 3700 11172
rect 3752 11160 3758 11212
rect 3789 11203 3847 11209
rect 3789 11169 3801 11203
rect 3835 11200 3847 11203
rect 4065 11203 4123 11209
rect 4065 11200 4077 11203
rect 3835 11172 4077 11200
rect 3835 11169 3847 11172
rect 3789 11163 3847 11169
rect 4065 11169 4077 11172
rect 4111 11169 4123 11203
rect 4065 11163 4123 11169
rect 4080 11064 4108 11163
rect 4154 11160 4160 11212
rect 4212 11200 4218 11212
rect 4341 11203 4399 11209
rect 4341 11200 4353 11203
rect 4212 11172 4353 11200
rect 4212 11160 4218 11172
rect 4341 11169 4353 11172
rect 4387 11169 4399 11203
rect 4341 11163 4399 11169
rect 4249 11135 4307 11141
rect 4249 11101 4261 11135
rect 4295 11132 4307 11135
rect 4540 11132 4568 11299
rect 4890 11296 4896 11308
rect 4948 11296 4954 11348
rect 7006 11336 7012 11348
rect 6564 11308 7012 11336
rect 5077 11271 5135 11277
rect 5077 11237 5089 11271
rect 5123 11268 5135 11271
rect 5123 11240 5672 11268
rect 5123 11237 5135 11240
rect 5077 11231 5135 11237
rect 4709 11203 4767 11209
rect 4709 11169 4721 11203
rect 4755 11200 4767 11203
rect 4893 11203 4951 11209
rect 4755 11172 4844 11200
rect 4755 11169 4767 11172
rect 4709 11163 4767 11169
rect 4295 11104 4568 11132
rect 4295 11101 4307 11104
rect 4249 11095 4307 11101
rect 4816 11064 4844 11172
rect 4893 11169 4905 11203
rect 4939 11200 4951 11203
rect 4982 11200 4988 11212
rect 4939 11172 4988 11200
rect 4939 11169 4951 11172
rect 4893 11163 4951 11169
rect 4982 11160 4988 11172
rect 5040 11160 5046 11212
rect 5442 11160 5448 11212
rect 5500 11160 5506 11212
rect 5644 11209 5672 11240
rect 5629 11203 5687 11209
rect 5629 11169 5641 11203
rect 5675 11200 5687 11203
rect 5902 11200 5908 11212
rect 5675 11172 5908 11200
rect 5675 11169 5687 11172
rect 5629 11163 5687 11169
rect 5902 11160 5908 11172
rect 5960 11160 5966 11212
rect 6564 11209 6592 11308
rect 7006 11296 7012 11308
rect 7064 11296 7070 11348
rect 7282 11296 7288 11348
rect 7340 11336 7346 11348
rect 8389 11339 8447 11345
rect 8389 11336 8401 11339
rect 7340 11308 8401 11336
rect 7340 11296 7346 11308
rect 8389 11305 8401 11308
rect 8435 11305 8447 11339
rect 8389 11299 8447 11305
rect 8754 11296 8760 11348
rect 8812 11296 8818 11348
rect 9306 11296 9312 11348
rect 9364 11336 9370 11348
rect 10134 11336 10140 11348
rect 9364 11308 10140 11336
rect 9364 11296 9370 11308
rect 10134 11296 10140 11308
rect 10192 11296 10198 11348
rect 11149 11339 11207 11345
rect 11149 11305 11161 11339
rect 11195 11336 11207 11339
rect 11609 11339 11667 11345
rect 11609 11336 11621 11339
rect 11195 11308 11621 11336
rect 11195 11305 11207 11308
rect 11149 11299 11207 11305
rect 11609 11305 11621 11308
rect 11655 11305 11667 11339
rect 11609 11299 11667 11305
rect 12066 11296 12072 11348
rect 12124 11336 12130 11348
rect 12124 11308 13492 11336
rect 12124 11296 12130 11308
rect 6641 11271 6699 11277
rect 6641 11237 6653 11271
rect 6687 11268 6699 11271
rect 6687 11240 7880 11268
rect 6687 11237 6699 11240
rect 6641 11231 6699 11237
rect 5997 11203 6055 11209
rect 5997 11169 6009 11203
rect 6043 11169 6055 11203
rect 5997 11163 6055 11169
rect 6549 11203 6607 11209
rect 6549 11169 6561 11203
rect 6595 11169 6607 11203
rect 6549 11163 6607 11169
rect 6733 11203 6791 11209
rect 6733 11169 6745 11203
rect 6779 11200 6791 11203
rect 6822 11200 6828 11212
rect 6779 11172 6828 11200
rect 6779 11169 6791 11172
rect 6733 11163 6791 11169
rect 5537 11135 5595 11141
rect 5537 11101 5549 11135
rect 5583 11132 5595 11135
rect 6012 11132 6040 11163
rect 5583 11104 6040 11132
rect 5583 11101 5595 11104
rect 5537 11095 5595 11101
rect 6086 11092 6092 11144
rect 6144 11092 6150 11144
rect 6365 11135 6423 11141
rect 6365 11101 6377 11135
rect 6411 11132 6423 11135
rect 6748 11132 6776 11163
rect 6822 11160 6828 11172
rect 6880 11160 6886 11212
rect 7009 11203 7067 11209
rect 7009 11169 7021 11203
rect 7055 11169 7067 11203
rect 7009 11163 7067 11169
rect 6411 11104 6776 11132
rect 6411 11101 6423 11104
rect 6365 11095 6423 11101
rect 6546 11064 6552 11076
rect 4080 11036 6552 11064
rect 6546 11024 6552 11036
rect 6604 11064 6610 11076
rect 7024 11064 7052 11163
rect 7282 11160 7288 11212
rect 7340 11200 7346 11212
rect 7852 11209 7880 11240
rect 11422 11228 11428 11280
rect 11480 11268 11486 11280
rect 11480 11240 11836 11268
rect 11480 11228 11486 11240
rect 7745 11203 7803 11209
rect 7745 11200 7757 11203
rect 7340 11172 7757 11200
rect 7340 11160 7346 11172
rect 7745 11169 7757 11172
rect 7791 11169 7803 11203
rect 7745 11163 7803 11169
rect 7837 11203 7895 11209
rect 7837 11169 7849 11203
rect 7883 11169 7895 11203
rect 7837 11163 7895 11169
rect 8570 11160 8576 11212
rect 8628 11160 8634 11212
rect 8662 11160 8668 11212
rect 8720 11200 8726 11212
rect 8849 11203 8907 11209
rect 8849 11200 8861 11203
rect 8720 11172 8861 11200
rect 8720 11160 8726 11172
rect 8849 11169 8861 11172
rect 8895 11169 8907 11203
rect 8849 11163 8907 11169
rect 9674 11160 9680 11212
rect 9732 11200 9738 11212
rect 10137 11203 10195 11209
rect 10137 11200 10149 11203
rect 9732 11172 10149 11200
rect 9732 11160 9738 11172
rect 10137 11169 10149 11172
rect 10183 11169 10195 11203
rect 10137 11163 10195 11169
rect 11054 11160 11060 11212
rect 11112 11160 11118 11212
rect 11146 11160 11152 11212
rect 11204 11200 11210 11212
rect 11333 11203 11391 11209
rect 11333 11200 11345 11203
rect 11204 11172 11345 11200
rect 11204 11160 11210 11172
rect 11333 11169 11345 11172
rect 11379 11169 11391 11203
rect 11333 11163 11391 11169
rect 7098 11092 7104 11144
rect 7156 11092 7162 11144
rect 7558 11092 7564 11144
rect 7616 11092 7622 11144
rect 7650 11092 7656 11144
rect 7708 11092 7714 11144
rect 8021 11135 8079 11141
rect 8021 11101 8033 11135
rect 8067 11132 8079 11135
rect 8386 11132 8392 11144
rect 8067 11104 8392 11132
rect 8067 11101 8079 11104
rect 8021 11095 8079 11101
rect 8386 11092 8392 11104
rect 8444 11092 8450 11144
rect 11348 11132 11376 11163
rect 11514 11160 11520 11212
rect 11572 11200 11578 11212
rect 11808 11209 11836 11240
rect 12342 11228 12348 11280
rect 12400 11268 12406 11280
rect 12437 11271 12495 11277
rect 12437 11268 12449 11271
rect 12400 11240 12449 11268
rect 12400 11228 12406 11240
rect 12437 11237 12449 11240
rect 12483 11237 12495 11271
rect 13078 11268 13084 11280
rect 12437 11231 12495 11237
rect 12912 11240 13084 11268
rect 11609 11203 11667 11209
rect 11609 11200 11621 11203
rect 11572 11172 11621 11200
rect 11572 11160 11578 11172
rect 11609 11169 11621 11172
rect 11655 11169 11667 11203
rect 11609 11163 11667 11169
rect 11793 11203 11851 11209
rect 11793 11169 11805 11203
rect 11839 11169 11851 11203
rect 11793 11163 11851 11169
rect 12066 11160 12072 11212
rect 12124 11200 12130 11212
rect 12161 11203 12219 11209
rect 12161 11200 12173 11203
rect 12124 11172 12173 11200
rect 12124 11160 12130 11172
rect 12161 11169 12173 11172
rect 12207 11169 12219 11203
rect 12161 11163 12219 11169
rect 12621 11203 12679 11209
rect 12621 11169 12633 11203
rect 12667 11169 12679 11203
rect 12621 11163 12679 11169
rect 12713 11203 12771 11209
rect 12713 11169 12725 11203
rect 12759 11200 12771 11203
rect 12912 11200 12940 11240
rect 13078 11228 13084 11240
rect 13136 11228 13142 11280
rect 13464 11277 13492 11308
rect 13998 11296 14004 11348
rect 14056 11296 14062 11348
rect 14921 11339 14979 11345
rect 14921 11305 14933 11339
rect 14967 11336 14979 11339
rect 15657 11339 15715 11345
rect 15657 11336 15669 11339
rect 14967 11308 15669 11336
rect 14967 11305 14979 11308
rect 14921 11299 14979 11305
rect 15657 11305 15669 11308
rect 15703 11305 15715 11339
rect 15657 11299 15715 11305
rect 16850 11296 16856 11348
rect 16908 11336 16914 11348
rect 17310 11336 17316 11348
rect 16908 11308 17316 11336
rect 16908 11296 16914 11308
rect 17310 11296 17316 11308
rect 17368 11296 17374 11348
rect 17770 11296 17776 11348
rect 17828 11336 17834 11348
rect 18509 11339 18567 11345
rect 18509 11336 18521 11339
rect 17828 11308 18521 11336
rect 17828 11296 17834 11308
rect 18509 11305 18521 11308
rect 18555 11305 18567 11339
rect 18509 11299 18567 11305
rect 18598 11296 18604 11348
rect 18656 11336 18662 11348
rect 20162 11336 20168 11348
rect 18656 11308 20168 11336
rect 18656 11296 18662 11308
rect 20162 11296 20168 11308
rect 20220 11296 20226 11348
rect 13449 11271 13507 11277
rect 13449 11237 13461 11271
rect 13495 11237 13507 11271
rect 13449 11231 13507 11237
rect 13538 11228 13544 11280
rect 13596 11268 13602 11280
rect 13596 11240 14044 11268
rect 13596 11228 13602 11240
rect 12759 11172 12940 11200
rect 12989 11203 13047 11209
rect 12759 11169 12771 11172
rect 12713 11163 12771 11169
rect 12989 11169 13001 11203
rect 13035 11169 13047 11203
rect 12989 11163 13047 11169
rect 11348 11104 12480 11132
rect 6604 11036 7052 11064
rect 7377 11067 7435 11073
rect 6604 11024 6610 11036
rect 7377 11033 7389 11067
rect 7423 11064 7435 11067
rect 8662 11064 8668 11076
rect 7423 11036 8668 11064
rect 7423 11033 7435 11036
rect 7377 11027 7435 11033
rect 8662 11024 8668 11036
rect 8720 11024 8726 11076
rect 11514 11024 11520 11076
rect 11572 11024 11578 11076
rect 11977 11067 12035 11073
rect 11977 11033 11989 11067
rect 12023 11064 12035 11067
rect 12158 11064 12164 11076
rect 12023 11036 12164 11064
rect 12023 11033 12035 11036
rect 11977 11027 12035 11033
rect 12158 11024 12164 11036
rect 12216 11024 12222 11076
rect 3421 10999 3479 11005
rect 3421 10996 3433 10999
rect 3200 10968 3433 10996
rect 3200 10956 3206 10968
rect 3421 10965 3433 10968
rect 3467 10965 3479 10999
rect 3421 10959 3479 10965
rect 7558 10956 7564 11008
rect 7616 10996 7622 11008
rect 8478 10996 8484 11008
rect 7616 10968 8484 10996
rect 7616 10956 7622 10968
rect 8478 10956 8484 10968
rect 8536 10956 8542 11008
rect 10321 10999 10379 11005
rect 10321 10965 10333 10999
rect 10367 10996 10379 10999
rect 10778 10996 10784 11008
rect 10367 10968 10784 10996
rect 10367 10965 10379 10968
rect 10321 10959 10379 10965
rect 10778 10956 10784 10968
rect 10836 10956 10842 11008
rect 12452 11005 12480 11104
rect 12636 11064 12664 11163
rect 12897 11067 12955 11073
rect 12897 11064 12909 11067
rect 12636 11036 12909 11064
rect 12897 11033 12909 11036
rect 12943 11033 12955 11067
rect 12897 11027 12955 11033
rect 12437 10999 12495 11005
rect 12437 10965 12449 10999
rect 12483 10996 12495 10999
rect 12618 10996 12624 11008
rect 12483 10968 12624 10996
rect 12483 10965 12495 10968
rect 12437 10959 12495 10965
rect 12618 10956 12624 10968
rect 12676 10956 12682 11008
rect 12802 10956 12808 11008
rect 12860 10996 12866 11008
rect 13004 10996 13032 11163
rect 13170 11160 13176 11212
rect 13228 11200 13234 11212
rect 13265 11203 13323 11209
rect 13265 11200 13277 11203
rect 13228 11172 13277 11200
rect 13228 11160 13234 11172
rect 13265 11169 13277 11172
rect 13311 11169 13323 11203
rect 13265 11163 13323 11169
rect 13354 11160 13360 11212
rect 13412 11160 13418 11212
rect 14016 11209 14044 11240
rect 14108 11240 15700 11268
rect 13633 11203 13691 11209
rect 13633 11169 13645 11203
rect 13679 11169 13691 11203
rect 13633 11163 13691 11169
rect 13725 11203 13783 11209
rect 13725 11169 13737 11203
rect 13771 11200 13783 11203
rect 13998 11203 14056 11209
rect 13771 11172 13952 11200
rect 13771 11169 13783 11172
rect 13725 11163 13783 11169
rect 13648 11132 13676 11163
rect 13924 11132 13952 11172
rect 13998 11169 14010 11203
rect 14044 11169 14056 11203
rect 13998 11163 14056 11169
rect 14108 11132 14136 11240
rect 15672 11212 15700 11240
rect 15746 11228 15752 11280
rect 15804 11268 15810 11280
rect 15841 11271 15899 11277
rect 15841 11268 15853 11271
rect 15804 11240 15853 11268
rect 15804 11228 15810 11240
rect 15841 11237 15853 11240
rect 15887 11237 15899 11271
rect 15841 11231 15899 11237
rect 17126 11228 17132 11280
rect 17184 11268 17190 11280
rect 20257 11271 20315 11277
rect 20257 11268 20269 11271
rect 17184 11240 20269 11268
rect 17184 11228 17190 11240
rect 14182 11160 14188 11212
rect 14240 11200 14246 11212
rect 14369 11203 14427 11209
rect 14369 11200 14381 11203
rect 14240 11172 14381 11200
rect 14240 11160 14246 11172
rect 14369 11169 14381 11172
rect 14415 11169 14427 11203
rect 14369 11163 14427 11169
rect 14458 11160 14464 11212
rect 14516 11160 14522 11212
rect 14642 11160 14648 11212
rect 14700 11200 14706 11212
rect 14737 11203 14795 11209
rect 14737 11200 14749 11203
rect 14700 11172 14749 11200
rect 14700 11160 14706 11172
rect 14737 11169 14749 11172
rect 14783 11169 14795 11203
rect 14737 11163 14795 11169
rect 14274 11132 14280 11144
rect 13648 11104 13860 11132
rect 13924 11104 14280 11132
rect 13081 11067 13139 11073
rect 13081 11033 13093 11067
rect 13127 11064 13139 11067
rect 13170 11064 13176 11076
rect 13127 11036 13176 11064
rect 13127 11033 13139 11036
rect 13081 11027 13139 11033
rect 13170 11024 13176 11036
rect 13228 11024 13234 11076
rect 13832 11073 13860 11104
rect 14274 11092 14280 11104
rect 14332 11092 14338 11144
rect 14752 11132 14780 11163
rect 14918 11160 14924 11212
rect 14976 11200 14982 11212
rect 15013 11203 15071 11209
rect 15013 11200 15025 11203
rect 14976 11172 15025 11200
rect 14976 11160 14982 11172
rect 15013 11169 15025 11172
rect 15059 11169 15071 11203
rect 15013 11163 15071 11169
rect 15289 11203 15347 11209
rect 15289 11169 15301 11203
rect 15335 11200 15347 11203
rect 15378 11200 15384 11212
rect 15335 11172 15384 11200
rect 15335 11169 15347 11172
rect 15289 11163 15347 11169
rect 15378 11160 15384 11172
rect 15436 11160 15442 11212
rect 15473 11203 15531 11209
rect 15473 11169 15485 11203
rect 15519 11200 15531 11203
rect 15565 11203 15623 11209
rect 15565 11200 15577 11203
rect 15519 11172 15577 11200
rect 15519 11169 15531 11172
rect 15473 11163 15531 11169
rect 15565 11169 15577 11172
rect 15611 11169 15623 11203
rect 15565 11163 15623 11169
rect 15654 11160 15660 11212
rect 15712 11160 15718 11212
rect 16298 11160 16304 11212
rect 16356 11160 16362 11212
rect 15105 11135 15163 11141
rect 15105 11132 15117 11135
rect 14752 11104 15117 11132
rect 15105 11101 15117 11104
rect 15151 11101 15163 11135
rect 15105 11095 15163 11101
rect 15194 11092 15200 11144
rect 15252 11132 15258 11144
rect 15746 11132 15752 11144
rect 15252 11104 15752 11132
rect 15252 11092 15258 11104
rect 15746 11092 15752 11104
rect 15804 11132 15810 11144
rect 16316 11132 16344 11160
rect 17129 11135 17187 11141
rect 17129 11132 17141 11135
rect 15804 11104 16160 11132
rect 16316 11104 17141 11132
rect 15804 11092 15810 11104
rect 16132 11073 16160 11104
rect 17129 11101 17141 11104
rect 17175 11101 17187 11135
rect 17236 11132 17264 11240
rect 20257 11237 20269 11240
rect 20303 11237 20315 11271
rect 21266 11268 21272 11280
rect 20257 11231 20315 11237
rect 20548 11240 21272 11268
rect 17310 11160 17316 11212
rect 17368 11200 17374 11212
rect 17862 11200 17868 11212
rect 17368 11172 17868 11200
rect 17368 11160 17374 11172
rect 17862 11160 17868 11172
rect 17920 11200 17926 11212
rect 18417 11203 18475 11209
rect 18417 11200 18429 11203
rect 17920 11172 18429 11200
rect 17920 11160 17926 11172
rect 18417 11169 18429 11172
rect 18463 11169 18475 11203
rect 18417 11163 18475 11169
rect 18601 11203 18659 11209
rect 18601 11169 18613 11203
rect 18647 11169 18659 11203
rect 18601 11163 18659 11169
rect 17405 11135 17463 11141
rect 17405 11132 17417 11135
rect 17236 11104 17417 11132
rect 17129 11095 17187 11101
rect 17405 11101 17417 11104
rect 17451 11101 17463 11135
rect 17405 11095 17463 11101
rect 17497 11135 17555 11141
rect 17497 11101 17509 11135
rect 17543 11101 17555 11135
rect 17497 11095 17555 11101
rect 13817 11067 13875 11073
rect 13817 11033 13829 11067
rect 13863 11033 13875 11067
rect 16117 11067 16175 11073
rect 13817 11027 13875 11033
rect 13924 11036 15976 11064
rect 13924 10996 13952 11036
rect 12860 10968 13952 10996
rect 12860 10956 12866 10968
rect 15286 10956 15292 11008
rect 15344 10996 15350 11008
rect 15841 10999 15899 11005
rect 15841 10996 15853 10999
rect 15344 10968 15853 10996
rect 15344 10956 15350 10968
rect 15841 10965 15853 10968
rect 15887 10965 15899 10999
rect 15948 10996 15976 11036
rect 16117 11033 16129 11067
rect 16163 11033 16175 11067
rect 17512 11064 17540 11095
rect 17770 11092 17776 11144
rect 17828 11092 17834 11144
rect 17954 11092 17960 11144
rect 18012 11132 18018 11144
rect 18616 11132 18644 11163
rect 18690 11160 18696 11212
rect 18748 11160 18754 11212
rect 18877 11203 18935 11209
rect 18877 11169 18889 11203
rect 18923 11200 18935 11203
rect 19058 11200 19064 11212
rect 18923 11172 19064 11200
rect 18923 11169 18935 11172
rect 18877 11163 18935 11169
rect 19058 11160 19064 11172
rect 19116 11160 19122 11212
rect 19153 11203 19211 11209
rect 19153 11169 19165 11203
rect 19199 11200 19211 11203
rect 19245 11203 19303 11209
rect 19245 11200 19257 11203
rect 19199 11172 19257 11200
rect 19199 11169 19211 11172
rect 19153 11163 19211 11169
rect 19245 11169 19257 11172
rect 19291 11169 19303 11203
rect 19245 11163 19303 11169
rect 19889 11203 19947 11209
rect 19889 11169 19901 11203
rect 19935 11169 19947 11203
rect 19889 11163 19947 11169
rect 18012 11104 18644 11132
rect 18785 11135 18843 11141
rect 18012 11092 18018 11104
rect 18785 11101 18797 11135
rect 18831 11132 18843 11135
rect 19168 11132 19196 11163
rect 18831 11104 19196 11132
rect 18831 11101 18843 11104
rect 18785 11095 18843 11101
rect 18322 11064 18328 11076
rect 17512 11036 18328 11064
rect 16117 11027 16175 11033
rect 18322 11024 18328 11036
rect 18380 11024 18386 11076
rect 18690 11024 18696 11076
rect 18748 11064 18754 11076
rect 18800 11064 18828 11095
rect 19334 11092 19340 11144
rect 19392 11132 19398 11144
rect 19705 11135 19763 11141
rect 19705 11132 19717 11135
rect 19392 11104 19717 11132
rect 19392 11092 19398 11104
rect 19705 11101 19717 11104
rect 19751 11101 19763 11135
rect 19904 11132 19932 11163
rect 20070 11160 20076 11212
rect 20128 11160 20134 11212
rect 20162 11160 20168 11212
rect 20220 11160 20226 11212
rect 20548 11209 20576 11240
rect 21266 11228 21272 11240
rect 21324 11268 21330 11280
rect 21726 11268 21732 11280
rect 21324 11240 21732 11268
rect 21324 11228 21330 11240
rect 21726 11228 21732 11240
rect 21784 11228 21790 11280
rect 21904 11271 21962 11277
rect 21904 11237 21916 11271
rect 21950 11268 21962 11271
rect 22186 11268 22192 11280
rect 21950 11240 22192 11268
rect 21950 11237 21962 11240
rect 21904 11231 21962 11237
rect 22186 11228 22192 11240
rect 22244 11228 22250 11280
rect 20349 11203 20407 11209
rect 20349 11169 20361 11203
rect 20395 11169 20407 11203
rect 20349 11163 20407 11169
rect 20533 11203 20591 11209
rect 20533 11169 20545 11203
rect 20579 11169 20591 11203
rect 20533 11163 20591 11169
rect 20364 11132 20392 11163
rect 20622 11160 20628 11212
rect 20680 11200 20686 11212
rect 20717 11203 20775 11209
rect 20717 11200 20729 11203
rect 20680 11172 20729 11200
rect 20680 11160 20686 11172
rect 20717 11169 20729 11172
rect 20763 11169 20775 11203
rect 20717 11163 20775 11169
rect 20898 11160 20904 11212
rect 20956 11200 20962 11212
rect 21082 11200 21088 11212
rect 20956 11172 21088 11200
rect 20956 11160 20962 11172
rect 21082 11160 21088 11172
rect 21140 11160 21146 11212
rect 21453 11203 21511 11209
rect 21453 11169 21465 11203
rect 21499 11200 21511 11203
rect 21542 11200 21548 11212
rect 21499 11172 21548 11200
rect 21499 11169 21511 11172
rect 21453 11163 21511 11169
rect 21542 11160 21548 11172
rect 21600 11160 21606 11212
rect 21634 11160 21640 11212
rect 21692 11160 21698 11212
rect 20640 11132 20668 11160
rect 19904 11104 20668 11132
rect 19705 11095 19763 11101
rect 18748 11036 18828 11064
rect 18892 11036 19656 11064
rect 18748 11024 18754 11036
rect 18892 10996 18920 11036
rect 15948 10968 18920 10996
rect 18969 10999 19027 11005
rect 15841 10959 15899 10965
rect 18969 10965 18981 10999
rect 19015 10996 19027 10999
rect 19334 10996 19340 11008
rect 19015 10968 19340 10996
rect 19015 10965 19027 10968
rect 18969 10959 19027 10965
rect 19334 10956 19340 10968
rect 19392 10956 19398 11008
rect 19429 10999 19487 11005
rect 19429 10965 19441 10999
rect 19475 10996 19487 10999
rect 19518 10996 19524 11008
rect 19475 10968 19524 10996
rect 19475 10965 19487 10968
rect 19429 10959 19487 10965
rect 19518 10956 19524 10968
rect 19576 10956 19582 11008
rect 19628 10996 19656 11036
rect 20254 11024 20260 11076
rect 20312 11064 20318 11076
rect 21269 11067 21327 11073
rect 21269 11064 21281 11067
rect 20312 11036 21281 11064
rect 20312 11024 20318 11036
rect 21269 11033 21281 11036
rect 21315 11033 21327 11067
rect 21269 11027 21327 11033
rect 20993 10999 21051 11005
rect 20993 10996 21005 10999
rect 19628 10968 21005 10996
rect 20993 10965 21005 10968
rect 21039 10965 21051 10999
rect 20993 10959 21051 10965
rect 23014 10956 23020 11008
rect 23072 10956 23078 11008
rect 552 10906 23368 10928
rect 552 10854 1366 10906
rect 1418 10854 1430 10906
rect 1482 10854 1494 10906
rect 1546 10854 1558 10906
rect 1610 10854 1622 10906
rect 1674 10854 1686 10906
rect 1738 10854 7366 10906
rect 7418 10854 7430 10906
rect 7482 10854 7494 10906
rect 7546 10854 7558 10906
rect 7610 10854 7622 10906
rect 7674 10854 7686 10906
rect 7738 10854 13366 10906
rect 13418 10854 13430 10906
rect 13482 10854 13494 10906
rect 13546 10854 13558 10906
rect 13610 10854 13622 10906
rect 13674 10854 13686 10906
rect 13738 10854 19366 10906
rect 19418 10854 19430 10906
rect 19482 10854 19494 10906
rect 19546 10854 19558 10906
rect 19610 10854 19622 10906
rect 19674 10854 19686 10906
rect 19738 10854 23368 10906
rect 552 10832 23368 10854
rect 1210 10752 1216 10804
rect 1268 10752 1274 10804
rect 1762 10752 1768 10804
rect 1820 10792 1826 10804
rect 1857 10795 1915 10801
rect 1857 10792 1869 10795
rect 1820 10764 1869 10792
rect 1820 10752 1826 10764
rect 1857 10761 1869 10764
rect 1903 10761 1915 10795
rect 1857 10755 1915 10761
rect 5353 10795 5411 10801
rect 5353 10761 5365 10795
rect 5399 10792 5411 10795
rect 5442 10792 5448 10804
rect 5399 10764 5448 10792
rect 5399 10761 5411 10764
rect 5353 10755 5411 10761
rect 5442 10752 5448 10764
rect 5500 10752 5506 10804
rect 6365 10795 6423 10801
rect 6365 10761 6377 10795
rect 6411 10792 6423 10795
rect 6546 10792 6552 10804
rect 6411 10764 6552 10792
rect 6411 10761 6423 10764
rect 6365 10755 6423 10761
rect 6546 10752 6552 10764
rect 6604 10752 6610 10804
rect 6914 10752 6920 10804
rect 6972 10752 6978 10804
rect 7282 10752 7288 10804
rect 7340 10792 7346 10804
rect 7377 10795 7435 10801
rect 7377 10792 7389 10795
rect 7340 10764 7389 10792
rect 7340 10752 7346 10764
rect 7377 10761 7389 10764
rect 7423 10761 7435 10795
rect 7377 10755 7435 10761
rect 7742 10752 7748 10804
rect 7800 10792 7806 10804
rect 8018 10792 8024 10804
rect 7800 10764 8024 10792
rect 7800 10752 7806 10764
rect 8018 10752 8024 10764
rect 8076 10752 8082 10804
rect 10226 10752 10232 10804
rect 10284 10792 10290 10804
rect 11149 10795 11207 10801
rect 10284 10764 11100 10792
rect 10284 10752 10290 10764
rect 1026 10684 1032 10736
rect 1084 10724 1090 10736
rect 1397 10727 1455 10733
rect 1397 10724 1409 10727
rect 1084 10696 1409 10724
rect 1084 10684 1090 10696
rect 1397 10693 1409 10696
rect 1443 10693 1455 10727
rect 1397 10687 1455 10693
rect 1780 10656 1808 10752
rect 3881 10727 3939 10733
rect 3881 10693 3893 10727
rect 3927 10724 3939 10727
rect 3927 10696 4292 10724
rect 3927 10693 3939 10696
rect 3881 10687 3939 10693
rect 1320 10628 1808 10656
rect 2041 10659 2099 10665
rect 934 10548 940 10600
rect 992 10588 998 10600
rect 1320 10597 1348 10628
rect 2041 10625 2053 10659
rect 2087 10656 2099 10659
rect 2406 10656 2412 10668
rect 2087 10628 2412 10656
rect 2087 10625 2099 10628
rect 2041 10619 2099 10625
rect 2406 10616 2412 10628
rect 2464 10616 2470 10668
rect 3326 10616 3332 10668
rect 3384 10656 3390 10668
rect 4264 10665 4292 10696
rect 3421 10659 3479 10665
rect 3421 10656 3433 10659
rect 3384 10628 3433 10656
rect 3384 10616 3390 10628
rect 3421 10625 3433 10628
rect 3467 10625 3479 10659
rect 3421 10619 3479 10625
rect 4249 10659 4307 10665
rect 4249 10625 4261 10659
rect 4295 10625 4307 10659
rect 5460 10656 5488 10752
rect 6086 10684 6092 10736
rect 6144 10724 6150 10736
rect 8294 10724 8300 10736
rect 6144 10696 8300 10724
rect 6144 10684 6150 10696
rect 8294 10684 8300 10696
rect 8352 10684 8358 10736
rect 9033 10727 9091 10733
rect 9033 10693 9045 10727
rect 9079 10724 9091 10727
rect 9079 10696 10088 10724
rect 9079 10693 9091 10696
rect 9033 10687 9091 10693
rect 5537 10659 5595 10665
rect 5537 10656 5549 10659
rect 5460 10628 5549 10656
rect 4249 10619 4307 10625
rect 5537 10625 5549 10628
rect 5583 10625 5595 10659
rect 5537 10619 5595 10625
rect 5902 10616 5908 10668
rect 5960 10616 5966 10668
rect 5994 10616 6000 10668
rect 6052 10616 6058 10668
rect 10060 10665 10088 10696
rect 10134 10684 10140 10736
rect 10192 10724 10198 10736
rect 10505 10727 10563 10733
rect 10505 10724 10517 10727
rect 10192 10696 10517 10724
rect 10192 10684 10198 10696
rect 10505 10693 10517 10696
rect 10551 10693 10563 10727
rect 10796 10724 10824 10764
rect 10505 10687 10563 10693
rect 10704 10696 10824 10724
rect 8757 10659 8815 10665
rect 6196 10628 6776 10656
rect 6196 10600 6224 10628
rect 1029 10591 1087 10597
rect 1029 10588 1041 10591
rect 992 10560 1041 10588
rect 992 10548 998 10560
rect 1029 10557 1041 10560
rect 1075 10557 1087 10591
rect 1029 10551 1087 10557
rect 1305 10591 1363 10597
rect 1305 10557 1317 10591
rect 1351 10557 1363 10591
rect 1305 10551 1363 10557
rect 1489 10591 1547 10597
rect 1489 10557 1501 10591
rect 1535 10557 1547 10591
rect 1489 10551 1547 10557
rect 1673 10591 1731 10597
rect 1673 10557 1685 10591
rect 1719 10588 1731 10591
rect 2222 10588 2228 10600
rect 1719 10560 2228 10588
rect 1719 10557 1731 10560
rect 1673 10551 1731 10557
rect 1504 10520 1532 10551
rect 2222 10548 2228 10560
rect 2280 10588 2286 10600
rect 2317 10591 2375 10597
rect 2317 10588 2329 10591
rect 2280 10560 2329 10588
rect 2280 10548 2286 10560
rect 2317 10557 2329 10560
rect 2363 10557 2375 10591
rect 2317 10551 2375 10557
rect 3513 10591 3571 10597
rect 3513 10557 3525 10591
rect 3559 10588 3571 10591
rect 3602 10588 3608 10600
rect 3559 10560 3608 10588
rect 3559 10557 3571 10560
rect 3513 10551 3571 10557
rect 3602 10548 3608 10560
rect 3660 10548 3666 10600
rect 4338 10548 4344 10600
rect 4396 10548 4402 10600
rect 5258 10548 5264 10600
rect 5316 10548 5322 10600
rect 5445 10591 5503 10597
rect 5445 10557 5457 10591
rect 5491 10588 5503 10591
rect 6178 10588 6184 10600
rect 5491 10560 6184 10588
rect 5491 10557 5503 10560
rect 5445 10551 5503 10557
rect 6178 10548 6184 10560
rect 6236 10548 6242 10600
rect 6546 10548 6552 10600
rect 6604 10548 6610 10600
rect 6748 10597 6776 10628
rect 8757 10625 8769 10659
rect 8803 10656 8815 10659
rect 10045 10659 10103 10665
rect 8803 10628 9352 10656
rect 8803 10625 8815 10628
rect 8757 10619 8815 10625
rect 6733 10591 6791 10597
rect 6733 10557 6745 10591
rect 6779 10557 6791 10591
rect 6733 10551 6791 10557
rect 6822 10548 6828 10600
rect 6880 10588 6886 10600
rect 7193 10591 7251 10597
rect 7193 10588 7205 10591
rect 6880 10560 7205 10588
rect 6880 10548 6886 10560
rect 7193 10557 7205 10560
rect 7239 10557 7251 10591
rect 7193 10551 7251 10557
rect 8662 10548 8668 10600
rect 8720 10588 8726 10600
rect 9324 10597 9352 10628
rect 10045 10625 10057 10659
rect 10091 10656 10103 10659
rect 10091 10628 10548 10656
rect 10091 10625 10103 10628
rect 10045 10619 10103 10625
rect 9125 10591 9183 10597
rect 9125 10588 9137 10591
rect 8720 10560 9137 10588
rect 8720 10548 8726 10560
rect 9125 10557 9137 10560
rect 9171 10557 9183 10591
rect 9125 10551 9183 10557
rect 9309 10591 9367 10597
rect 9309 10557 9321 10591
rect 9355 10588 9367 10591
rect 9398 10588 9404 10600
rect 9355 10560 9404 10588
rect 9355 10557 9367 10560
rect 9309 10551 9367 10557
rect 9398 10548 9404 10560
rect 9456 10548 9462 10600
rect 10137 10591 10195 10597
rect 10137 10557 10149 10591
rect 10183 10557 10195 10591
rect 10137 10551 10195 10557
rect 1946 10520 1952 10532
rect 1504 10492 1952 10520
rect 1946 10480 1952 10492
rect 2004 10480 2010 10532
rect 4724 10492 6960 10520
rect 4724 10461 4752 10492
rect 4709 10455 4767 10461
rect 4709 10421 4721 10455
rect 4755 10421 4767 10455
rect 4709 10415 4767 10421
rect 6181 10455 6239 10461
rect 6181 10421 6193 10455
rect 6227 10452 6239 10455
rect 6454 10452 6460 10464
rect 6227 10424 6460 10452
rect 6227 10421 6239 10424
rect 6181 10415 6239 10421
rect 6454 10412 6460 10424
rect 6512 10412 6518 10464
rect 6932 10452 6960 10492
rect 7006 10480 7012 10532
rect 7064 10480 7070 10532
rect 10152 10520 10180 10551
rect 10226 10548 10232 10600
rect 10284 10548 10290 10600
rect 10318 10548 10324 10600
rect 10376 10548 10382 10600
rect 10520 10597 10548 10628
rect 10704 10597 10732 10696
rect 10870 10684 10876 10736
rect 10928 10684 10934 10736
rect 11072 10724 11100 10764
rect 11149 10761 11161 10795
rect 11195 10792 11207 10795
rect 11195 10764 13952 10792
rect 11195 10761 11207 10764
rect 11149 10755 11207 10761
rect 11974 10724 11980 10736
rect 11072 10696 11980 10724
rect 11974 10684 11980 10696
rect 12032 10684 12038 10736
rect 12161 10727 12219 10733
rect 12161 10693 12173 10727
rect 12207 10724 12219 10727
rect 13814 10724 13820 10736
rect 12207 10696 13820 10724
rect 12207 10693 12219 10696
rect 12161 10687 12219 10693
rect 13814 10684 13820 10696
rect 13872 10684 13878 10736
rect 13924 10724 13952 10764
rect 13998 10752 14004 10804
rect 14056 10792 14062 10804
rect 14185 10795 14243 10801
rect 14185 10792 14197 10795
rect 14056 10764 14197 10792
rect 14056 10752 14062 10764
rect 14185 10761 14197 10764
rect 14231 10761 14243 10795
rect 14185 10755 14243 10761
rect 14829 10795 14887 10801
rect 14829 10761 14841 10795
rect 14875 10792 14887 10795
rect 15194 10792 15200 10804
rect 14875 10764 15200 10792
rect 14875 10761 14887 10764
rect 14829 10755 14887 10761
rect 15194 10752 15200 10764
rect 15252 10752 15258 10804
rect 15838 10752 15844 10804
rect 15896 10792 15902 10804
rect 16577 10795 16635 10801
rect 16577 10792 16589 10795
rect 15896 10764 16589 10792
rect 15896 10752 15902 10764
rect 16577 10761 16589 10764
rect 16623 10761 16635 10795
rect 16577 10755 16635 10761
rect 16758 10752 16764 10804
rect 16816 10792 16822 10804
rect 16942 10792 16948 10804
rect 16816 10764 16948 10792
rect 16816 10752 16822 10764
rect 16942 10752 16948 10764
rect 17000 10752 17006 10804
rect 17586 10752 17592 10804
rect 17644 10792 17650 10804
rect 17773 10795 17831 10801
rect 17773 10792 17785 10795
rect 17644 10764 17785 10792
rect 17644 10752 17650 10764
rect 17773 10761 17785 10764
rect 17819 10761 17831 10795
rect 17773 10755 17831 10761
rect 20073 10795 20131 10801
rect 20073 10761 20085 10795
rect 20119 10792 20131 10795
rect 20162 10792 20168 10804
rect 20119 10764 20168 10792
rect 20119 10761 20131 10764
rect 20073 10755 20131 10761
rect 20162 10752 20168 10764
rect 20220 10752 20226 10804
rect 21361 10795 21419 10801
rect 21361 10761 21373 10795
rect 21407 10792 21419 10795
rect 22094 10792 22100 10804
rect 21407 10764 22100 10792
rect 21407 10761 21419 10764
rect 21361 10755 21419 10761
rect 22094 10752 22100 10764
rect 22152 10752 22158 10804
rect 22278 10752 22284 10804
rect 22336 10792 22342 10804
rect 22465 10795 22523 10801
rect 22465 10792 22477 10795
rect 22336 10764 22477 10792
rect 22336 10752 22342 10764
rect 22465 10761 22477 10764
rect 22511 10761 22523 10795
rect 22465 10755 22523 10761
rect 14366 10724 14372 10736
rect 13924 10696 14372 10724
rect 14366 10684 14372 10696
rect 14424 10684 14430 10736
rect 20717 10727 20775 10733
rect 20717 10724 20729 10727
rect 14660 10696 20729 10724
rect 10888 10656 10916 10684
rect 10796 10628 10916 10656
rect 10796 10597 10824 10628
rect 11606 10616 11612 10668
rect 11664 10616 11670 10668
rect 11701 10659 11759 10665
rect 11701 10625 11713 10659
rect 11747 10656 11759 10659
rect 12066 10656 12072 10668
rect 11747 10628 12072 10656
rect 11747 10625 11759 10628
rect 11701 10619 11759 10625
rect 12066 10616 12072 10628
rect 12124 10616 12130 10668
rect 12526 10616 12532 10668
rect 12584 10656 12590 10668
rect 12805 10659 12863 10665
rect 12805 10656 12817 10659
rect 12584 10628 12817 10656
rect 12584 10616 12590 10628
rect 12805 10625 12817 10628
rect 12851 10625 12863 10659
rect 12805 10619 12863 10625
rect 12894 10616 12900 10668
rect 12952 10656 12958 10668
rect 12952 10628 13400 10656
rect 12952 10616 12958 10628
rect 13372 10600 13400 10628
rect 10505 10591 10563 10597
rect 10505 10557 10517 10591
rect 10551 10557 10563 10591
rect 10505 10551 10563 10557
rect 10689 10591 10747 10597
rect 10689 10557 10701 10591
rect 10735 10557 10747 10591
rect 10689 10551 10747 10557
rect 10781 10591 10839 10597
rect 10781 10557 10793 10591
rect 10827 10557 10839 10591
rect 10781 10551 10839 10557
rect 10796 10520 10824 10551
rect 10870 10548 10876 10600
rect 10928 10548 10934 10600
rect 10965 10591 11023 10597
rect 10965 10557 10977 10591
rect 11011 10588 11023 10591
rect 11330 10588 11336 10600
rect 11011 10560 11336 10588
rect 11011 10557 11023 10560
rect 10965 10551 11023 10557
rect 11330 10548 11336 10560
rect 11388 10548 11394 10600
rect 11422 10548 11428 10600
rect 11480 10548 11486 10600
rect 11974 10548 11980 10600
rect 12032 10548 12038 10600
rect 12161 10591 12219 10597
rect 12161 10557 12173 10591
rect 12207 10588 12219 10591
rect 12250 10588 12256 10600
rect 12207 10560 12256 10588
rect 12207 10557 12219 10560
rect 12161 10551 12219 10557
rect 12250 10548 12256 10560
rect 12308 10548 12314 10600
rect 12618 10548 12624 10600
rect 12676 10548 12682 10600
rect 12713 10591 12771 10597
rect 12713 10557 12725 10591
rect 12759 10557 12771 10591
rect 12713 10551 12771 10557
rect 8128 10492 10088 10520
rect 10152 10492 10824 10520
rect 8128 10452 8156 10492
rect 6932 10424 8156 10452
rect 8202 10412 8208 10464
rect 8260 10452 8266 10464
rect 9217 10455 9275 10461
rect 9217 10452 9229 10455
rect 8260 10424 9229 10452
rect 8260 10412 8266 10424
rect 9217 10421 9229 10424
rect 9263 10421 9275 10455
rect 9217 10415 9275 10421
rect 9861 10455 9919 10461
rect 9861 10421 9873 10455
rect 9907 10452 9919 10455
rect 9950 10452 9956 10464
rect 9907 10424 9956 10452
rect 9907 10421 9919 10424
rect 9861 10415 9919 10421
rect 9950 10412 9956 10424
rect 10008 10412 10014 10464
rect 10060 10452 10088 10492
rect 11146 10480 11152 10532
rect 11204 10520 11210 10532
rect 11241 10523 11299 10529
rect 11241 10520 11253 10523
rect 11204 10492 11253 10520
rect 11204 10480 11210 10492
rect 11241 10489 11253 10492
rect 11287 10489 11299 10523
rect 11241 10483 11299 10489
rect 11793 10523 11851 10529
rect 11793 10489 11805 10523
rect 11839 10489 11851 10523
rect 11793 10483 11851 10489
rect 10870 10452 10876 10464
rect 10060 10424 10876 10452
rect 10870 10412 10876 10424
rect 10928 10412 10934 10464
rect 11808 10452 11836 10483
rect 12728 10464 12756 10551
rect 12986 10548 12992 10600
rect 13044 10588 13050 10600
rect 13081 10591 13139 10597
rect 13081 10588 13093 10591
rect 13044 10560 13093 10588
rect 13044 10548 13050 10560
rect 13081 10557 13093 10560
rect 13127 10557 13139 10591
rect 13081 10551 13139 10557
rect 13354 10548 13360 10600
rect 13412 10588 13418 10600
rect 13633 10591 13691 10597
rect 13633 10588 13645 10591
rect 13412 10560 13645 10588
rect 13412 10548 13418 10560
rect 13633 10557 13645 10560
rect 13679 10557 13691 10591
rect 13633 10551 13691 10557
rect 13906 10548 13912 10600
rect 13964 10588 13970 10600
rect 14660 10597 14688 10696
rect 20717 10693 20729 10696
rect 20763 10693 20775 10727
rect 20717 10687 20775 10693
rect 14734 10616 14740 10668
rect 14792 10656 14798 10668
rect 15013 10659 15071 10665
rect 15013 10656 15025 10659
rect 14792 10628 15025 10656
rect 14792 10616 14798 10628
rect 15013 10625 15025 10628
rect 15059 10625 15071 10659
rect 15013 10619 15071 10625
rect 15102 10616 15108 10668
rect 15160 10616 15166 10668
rect 15286 10616 15292 10668
rect 15344 10616 15350 10668
rect 15746 10616 15752 10668
rect 15804 10656 15810 10668
rect 15804 10628 16160 10656
rect 15804 10616 15810 10628
rect 14093 10591 14151 10597
rect 14093 10588 14105 10591
rect 13964 10560 14105 10588
rect 13964 10548 13970 10560
rect 14093 10557 14105 10560
rect 14139 10557 14151 10591
rect 14093 10551 14151 10557
rect 14277 10591 14335 10597
rect 14277 10557 14289 10591
rect 14323 10588 14335 10591
rect 14645 10591 14703 10597
rect 14645 10588 14657 10591
rect 14323 10560 14657 10588
rect 14323 10557 14335 10560
rect 14277 10551 14335 10557
rect 14645 10557 14657 10560
rect 14691 10557 14703 10591
rect 14645 10551 14703 10557
rect 15197 10591 15255 10597
rect 15197 10557 15209 10591
rect 15243 10557 15255 10591
rect 15197 10551 15255 10557
rect 15102 10480 15108 10532
rect 15160 10480 15166 10532
rect 15212 10520 15240 10551
rect 15654 10548 15660 10600
rect 15712 10588 15718 10600
rect 16132 10597 16160 10628
rect 16206 10616 16212 10668
rect 16264 10616 16270 10668
rect 16666 10616 16672 10668
rect 16724 10656 16730 10668
rect 17037 10659 17095 10665
rect 17037 10656 17049 10659
rect 16724 10628 17049 10656
rect 16724 10616 16730 10628
rect 17037 10625 17049 10628
rect 17083 10625 17095 10659
rect 17770 10656 17776 10668
rect 17037 10619 17095 10625
rect 17512 10628 17776 10656
rect 15841 10591 15899 10597
rect 15841 10588 15853 10591
rect 15712 10560 15853 10588
rect 15712 10548 15718 10560
rect 15841 10557 15853 10560
rect 15887 10557 15899 10591
rect 15841 10551 15899 10557
rect 16117 10591 16175 10597
rect 16117 10557 16129 10591
rect 16163 10557 16175 10591
rect 16224 10588 16252 10616
rect 17512 10600 17540 10628
rect 17770 10616 17776 10628
rect 17828 10616 17834 10668
rect 18690 10616 18696 10668
rect 18748 10616 18754 10668
rect 20993 10659 21051 10665
rect 20993 10656 21005 10659
rect 20272 10628 21005 10656
rect 16301 10591 16359 10597
rect 16301 10588 16313 10591
rect 16224 10560 16313 10588
rect 16117 10551 16175 10557
rect 16301 10557 16313 10560
rect 16347 10557 16359 10591
rect 16301 10551 16359 10557
rect 16761 10591 16819 10597
rect 16761 10557 16773 10591
rect 16807 10557 16819 10591
rect 16761 10551 16819 10557
rect 15286 10520 15292 10532
rect 15212 10492 15292 10520
rect 15286 10480 15292 10492
rect 15344 10480 15350 10532
rect 15746 10480 15752 10532
rect 15804 10520 15810 10532
rect 15979 10523 16037 10529
rect 15979 10520 15991 10523
rect 15804 10492 15991 10520
rect 15804 10480 15810 10492
rect 15979 10489 15991 10492
rect 16025 10489 16037 10523
rect 15979 10483 16037 10489
rect 16206 10480 16212 10532
rect 16264 10480 16270 10532
rect 16776 10520 16804 10551
rect 16942 10548 16948 10600
rect 17000 10548 17006 10600
rect 17310 10548 17316 10600
rect 17368 10548 17374 10600
rect 17405 10591 17463 10597
rect 17405 10557 17417 10591
rect 17451 10588 17463 10591
rect 17494 10588 17500 10600
rect 17451 10560 17500 10588
rect 17451 10557 17463 10560
rect 17405 10551 17463 10557
rect 17494 10548 17500 10560
rect 17552 10548 17558 10600
rect 17586 10548 17592 10600
rect 17644 10548 17650 10600
rect 17678 10548 17684 10600
rect 17736 10588 17742 10600
rect 17865 10591 17923 10597
rect 17865 10588 17877 10591
rect 17736 10560 17877 10588
rect 17736 10548 17742 10560
rect 17865 10557 17877 10560
rect 17911 10557 17923 10591
rect 17865 10551 17923 10557
rect 18325 10591 18383 10597
rect 18325 10557 18337 10591
rect 18371 10557 18383 10591
rect 18325 10551 18383 10557
rect 18340 10520 18368 10551
rect 18414 10548 18420 10600
rect 18472 10588 18478 10600
rect 18509 10591 18567 10597
rect 18509 10588 18521 10591
rect 18472 10560 18521 10588
rect 18472 10548 18478 10560
rect 18509 10557 18521 10560
rect 18555 10557 18567 10591
rect 18509 10551 18567 10557
rect 18598 10548 18604 10600
rect 18656 10588 18662 10600
rect 18969 10591 19027 10597
rect 18969 10588 18981 10591
rect 18656 10560 18981 10588
rect 18656 10548 18662 10560
rect 18969 10557 18981 10560
rect 19015 10557 19027 10591
rect 18969 10551 19027 10557
rect 20070 10548 20076 10600
rect 20128 10588 20134 10600
rect 20272 10597 20300 10628
rect 20993 10625 21005 10628
rect 21039 10625 21051 10659
rect 20993 10619 21051 10625
rect 21818 10616 21824 10668
rect 21876 10616 21882 10668
rect 23382 10656 23388 10668
rect 22112 10628 23388 10656
rect 20257 10591 20315 10597
rect 20257 10588 20269 10591
rect 20128 10560 20269 10588
rect 20128 10548 20134 10560
rect 20257 10557 20269 10560
rect 20303 10557 20315 10591
rect 20257 10551 20315 10557
rect 20530 10548 20536 10600
rect 20588 10548 20594 10600
rect 20625 10591 20683 10597
rect 20625 10557 20637 10591
rect 20671 10588 20683 10591
rect 20714 10588 20720 10600
rect 20671 10560 20720 10588
rect 20671 10557 20683 10560
rect 20625 10551 20683 10557
rect 20714 10548 20720 10560
rect 20772 10548 20778 10600
rect 20809 10591 20867 10597
rect 20809 10557 20821 10591
rect 20855 10588 20867 10591
rect 20855 10560 20944 10588
rect 20855 10557 20867 10560
rect 20809 10551 20867 10557
rect 16309 10492 18368 10520
rect 12066 10452 12072 10464
rect 11808 10424 12072 10452
rect 12066 10412 12072 10424
rect 12124 10412 12130 10464
rect 12434 10412 12440 10464
rect 12492 10412 12498 10464
rect 12710 10412 12716 10464
rect 12768 10412 12774 10464
rect 13262 10412 13268 10464
rect 13320 10412 13326 10464
rect 13817 10455 13875 10461
rect 13817 10421 13829 10455
rect 13863 10452 13875 10455
rect 13906 10452 13912 10464
rect 13863 10424 13912 10452
rect 13863 10421 13875 10424
rect 13817 10415 13875 10421
rect 13906 10412 13912 10424
rect 13964 10452 13970 10464
rect 14274 10452 14280 10464
rect 13964 10424 14280 10452
rect 13964 10412 13970 10424
rect 14274 10412 14280 10424
rect 14332 10412 14338 10464
rect 14458 10412 14464 10464
rect 14516 10412 14522 10464
rect 15120 10452 15148 10480
rect 16309 10452 16337 10492
rect 19058 10480 19064 10532
rect 19116 10520 19122 10532
rect 19797 10523 19855 10529
rect 19797 10520 19809 10523
rect 19116 10492 19809 10520
rect 19116 10480 19122 10492
rect 19797 10489 19809 10492
rect 19843 10489 19855 10523
rect 19797 10483 19855 10489
rect 19981 10523 20039 10529
rect 19981 10489 19993 10523
rect 20027 10520 20039 10523
rect 20162 10520 20168 10532
rect 20027 10492 20168 10520
rect 20027 10489 20039 10492
rect 19981 10483 20039 10489
rect 15120 10424 16337 10452
rect 16390 10412 16396 10464
rect 16448 10452 16454 10464
rect 16485 10455 16543 10461
rect 16485 10452 16497 10455
rect 16448 10424 16497 10452
rect 16448 10412 16454 10424
rect 16485 10421 16497 10424
rect 16531 10421 16543 10455
rect 16485 10415 16543 10421
rect 17034 10412 17040 10464
rect 17092 10452 17098 10464
rect 17310 10452 17316 10464
rect 17092 10424 17316 10452
rect 17092 10412 17098 10424
rect 17310 10412 17316 10424
rect 17368 10412 17374 10464
rect 17954 10412 17960 10464
rect 18012 10452 18018 10464
rect 18049 10455 18107 10461
rect 18049 10452 18061 10455
rect 18012 10424 18061 10452
rect 18012 10412 18018 10424
rect 18049 10421 18061 10424
rect 18095 10421 18107 10455
rect 18049 10415 18107 10421
rect 18322 10412 18328 10464
rect 18380 10452 18386 10464
rect 18417 10455 18475 10461
rect 18417 10452 18429 10455
rect 18380 10424 18429 10452
rect 18380 10412 18386 10424
rect 18417 10421 18429 10424
rect 18463 10421 18475 10455
rect 18417 10415 18475 10421
rect 19426 10412 19432 10464
rect 19484 10452 19490 10464
rect 19613 10455 19671 10461
rect 19613 10452 19625 10455
rect 19484 10424 19625 10452
rect 19484 10412 19490 10424
rect 19613 10421 19625 10424
rect 19659 10421 19671 10455
rect 19812 10452 19840 10483
rect 20162 10480 20168 10492
rect 20220 10480 20226 10532
rect 20916 10464 20944 10560
rect 21082 10548 21088 10600
rect 21140 10588 21146 10600
rect 22112 10597 22140 10628
rect 23382 10616 23388 10628
rect 23440 10616 23446 10668
rect 21453 10591 21511 10597
rect 21453 10588 21465 10591
rect 21140 10560 21465 10588
rect 21140 10548 21146 10560
rect 21453 10557 21465 10560
rect 21499 10557 21511 10591
rect 21453 10551 21511 10557
rect 22097 10591 22155 10597
rect 22097 10557 22109 10591
rect 22143 10557 22155 10591
rect 22097 10551 22155 10557
rect 22741 10591 22799 10597
rect 22741 10557 22753 10591
rect 22787 10588 22799 10591
rect 23014 10588 23020 10600
rect 22787 10560 23020 10588
rect 22787 10557 22799 10560
rect 22741 10551 22799 10557
rect 23014 10548 23020 10560
rect 23072 10548 23078 10600
rect 22005 10523 22063 10529
rect 22005 10489 22017 10523
rect 22051 10520 22063 10523
rect 22051 10492 22600 10520
rect 22051 10489 22063 10492
rect 22005 10483 22063 10489
rect 20070 10452 20076 10464
rect 19812 10424 20076 10452
rect 19613 10415 19671 10421
rect 20070 10412 20076 10424
rect 20128 10412 20134 10464
rect 20349 10455 20407 10461
rect 20349 10421 20361 10455
rect 20395 10452 20407 10455
rect 20898 10452 20904 10464
rect 20395 10424 20904 10452
rect 20395 10421 20407 10424
rect 20349 10415 20407 10421
rect 20898 10412 20904 10424
rect 20956 10412 20962 10464
rect 22572 10461 22600 10492
rect 22557 10455 22615 10461
rect 22557 10421 22569 10455
rect 22603 10452 22615 10455
rect 22830 10452 22836 10464
rect 22603 10424 22836 10452
rect 22603 10421 22615 10424
rect 22557 10415 22615 10421
rect 22830 10412 22836 10424
rect 22888 10412 22894 10464
rect 22922 10412 22928 10464
rect 22980 10412 22986 10464
rect 552 10362 23368 10384
rect 552 10310 4366 10362
rect 4418 10310 4430 10362
rect 4482 10310 4494 10362
rect 4546 10310 4558 10362
rect 4610 10310 4622 10362
rect 4674 10310 4686 10362
rect 4738 10310 10366 10362
rect 10418 10310 10430 10362
rect 10482 10310 10494 10362
rect 10546 10310 10558 10362
rect 10610 10310 10622 10362
rect 10674 10310 10686 10362
rect 10738 10310 16366 10362
rect 16418 10310 16430 10362
rect 16482 10310 16494 10362
rect 16546 10310 16558 10362
rect 16610 10310 16622 10362
rect 16674 10310 16686 10362
rect 16738 10310 22366 10362
rect 22418 10310 22430 10362
rect 22482 10310 22494 10362
rect 22546 10310 22558 10362
rect 22610 10310 22622 10362
rect 22674 10310 22686 10362
rect 22738 10310 23368 10362
rect 552 10288 23368 10310
rect 3602 10208 3608 10260
rect 3660 10208 3666 10260
rect 4617 10251 4675 10257
rect 4617 10217 4629 10251
rect 4663 10248 4675 10251
rect 5258 10248 5264 10260
rect 4663 10220 5264 10248
rect 4663 10217 4675 10220
rect 4617 10211 4675 10217
rect 5258 10208 5264 10220
rect 5316 10248 5322 10260
rect 5442 10248 5448 10260
rect 5316 10220 5448 10248
rect 5316 10208 5322 10220
rect 5442 10208 5448 10220
rect 5500 10208 5506 10260
rect 6733 10251 6791 10257
rect 6733 10248 6745 10251
rect 6472 10220 6745 10248
rect 4062 10140 4068 10192
rect 4120 10180 4126 10192
rect 4157 10183 4215 10189
rect 4157 10180 4169 10183
rect 4120 10152 4169 10180
rect 4120 10140 4126 10152
rect 4157 10149 4169 10152
rect 4203 10149 4215 10183
rect 4157 10143 4215 10149
rect 842 10072 848 10124
rect 900 10072 906 10124
rect 1118 10121 1124 10124
rect 1112 10075 1124 10121
rect 1118 10072 1124 10075
rect 1176 10072 1182 10124
rect 1946 10072 1952 10124
rect 2004 10112 2010 10124
rect 2317 10115 2375 10121
rect 2317 10112 2329 10115
rect 2004 10084 2329 10112
rect 2004 10072 2010 10084
rect 2317 10081 2329 10084
rect 2363 10081 2375 10115
rect 2317 10075 2375 10081
rect 2590 10072 2596 10124
rect 2648 10072 2654 10124
rect 2777 10115 2835 10121
rect 2777 10081 2789 10115
rect 2823 10081 2835 10115
rect 2777 10075 2835 10081
rect 2501 9979 2559 9985
rect 2501 9945 2513 9979
rect 2547 9976 2559 9979
rect 2792 9976 2820 10075
rect 3142 10072 3148 10124
rect 3200 10072 3206 10124
rect 3970 10072 3976 10124
rect 4028 10072 4034 10124
rect 4172 10112 4200 10143
rect 5810 10140 5816 10192
rect 5868 10180 5874 10192
rect 5997 10183 6055 10189
rect 5997 10180 6009 10183
rect 5868 10152 6009 10180
rect 5868 10140 5874 10152
rect 5997 10149 6009 10152
rect 6043 10149 6055 10183
rect 5997 10143 6055 10149
rect 4433 10115 4491 10121
rect 4433 10112 4445 10115
rect 4172 10084 4445 10112
rect 4433 10081 4445 10084
rect 4479 10081 4491 10115
rect 4433 10075 4491 10081
rect 6012 10044 6040 10143
rect 6178 10140 6184 10192
rect 6236 10140 6242 10192
rect 6196 10112 6224 10140
rect 6472 10121 6500 10220
rect 6733 10217 6745 10220
rect 6779 10217 6791 10251
rect 6733 10211 6791 10217
rect 8478 10208 8484 10260
rect 8536 10248 8542 10260
rect 11146 10248 11152 10260
rect 8536 10220 11152 10248
rect 8536 10208 8542 10220
rect 11146 10208 11152 10220
rect 11204 10208 11210 10260
rect 11882 10208 11888 10260
rect 11940 10248 11946 10260
rect 11977 10251 12035 10257
rect 11977 10248 11989 10251
rect 11940 10220 11989 10248
rect 11940 10208 11946 10220
rect 11977 10217 11989 10220
rect 12023 10248 12035 10251
rect 12618 10248 12624 10260
rect 12023 10220 12624 10248
rect 12023 10217 12035 10220
rect 11977 10211 12035 10217
rect 12618 10208 12624 10220
rect 12676 10208 12682 10260
rect 12805 10251 12863 10257
rect 12805 10217 12817 10251
rect 12851 10248 12863 10251
rect 12894 10248 12900 10260
rect 12851 10220 12900 10248
rect 12851 10217 12863 10220
rect 12805 10211 12863 10217
rect 12894 10208 12900 10220
rect 12952 10208 12958 10260
rect 13078 10208 13084 10260
rect 13136 10248 13142 10260
rect 13136 10220 15608 10248
rect 13136 10208 13142 10220
rect 7668 10152 8064 10180
rect 6457 10115 6515 10121
rect 6457 10112 6469 10115
rect 6196 10084 6469 10112
rect 6457 10081 6469 10084
rect 6503 10081 6515 10115
rect 6457 10075 6515 10081
rect 6546 10072 6552 10124
rect 6604 10112 6610 10124
rect 6917 10115 6975 10121
rect 6917 10112 6929 10115
rect 6604 10084 6929 10112
rect 6604 10072 6610 10084
rect 6917 10081 6929 10084
rect 6963 10081 6975 10115
rect 6917 10075 6975 10081
rect 7098 10072 7104 10124
rect 7156 10112 7162 10124
rect 7193 10115 7251 10121
rect 7193 10112 7205 10115
rect 7156 10084 7205 10112
rect 7156 10072 7162 10084
rect 7193 10081 7205 10084
rect 7239 10081 7251 10115
rect 7193 10075 7251 10081
rect 7282 10072 7288 10124
rect 7340 10112 7346 10124
rect 7377 10115 7435 10121
rect 7377 10112 7389 10115
rect 7340 10084 7389 10112
rect 7340 10072 7346 10084
rect 7377 10081 7389 10084
rect 7423 10081 7435 10115
rect 7377 10075 7435 10081
rect 6641 10047 6699 10053
rect 6641 10044 6653 10047
rect 6012 10016 6653 10044
rect 6641 10013 6653 10016
rect 6687 10013 6699 10047
rect 6641 10007 6699 10013
rect 7006 10004 7012 10056
rect 7064 10044 7070 10056
rect 7668 10053 7696 10152
rect 8036 10121 8064 10152
rect 8386 10140 8392 10192
rect 8444 10180 8450 10192
rect 10962 10180 10968 10192
rect 8444 10152 8708 10180
rect 8444 10140 8450 10152
rect 7929 10115 7987 10121
rect 7929 10081 7941 10115
rect 7975 10081 7987 10115
rect 7929 10075 7987 10081
rect 8021 10115 8079 10121
rect 8021 10081 8033 10115
rect 8067 10081 8079 10115
rect 8021 10075 8079 10081
rect 7653 10047 7711 10053
rect 7653 10044 7665 10047
rect 7064 10016 7665 10044
rect 7064 10004 7070 10016
rect 7653 10013 7665 10016
rect 7699 10013 7711 10047
rect 7944 10044 7972 10075
rect 8202 10072 8208 10124
rect 8260 10072 8266 10124
rect 8680 10121 8708 10152
rect 9876 10152 10968 10180
rect 8481 10115 8539 10121
rect 8481 10081 8493 10115
rect 8527 10081 8539 10115
rect 8481 10075 8539 10081
rect 8665 10115 8723 10121
rect 8665 10081 8677 10115
rect 8711 10081 8723 10115
rect 8665 10075 8723 10081
rect 8220 10044 8248 10072
rect 7944 10016 8248 10044
rect 8496 10044 8524 10075
rect 8754 10072 8760 10124
rect 8812 10072 8818 10124
rect 8849 10115 8907 10121
rect 8849 10081 8861 10115
rect 8895 10112 8907 10115
rect 9030 10112 9036 10124
rect 8895 10084 9036 10112
rect 8895 10081 8907 10084
rect 8849 10075 8907 10081
rect 9030 10072 9036 10084
rect 9088 10072 9094 10124
rect 9214 10072 9220 10124
rect 9272 10072 9278 10124
rect 9398 10072 9404 10124
rect 9456 10112 9462 10124
rect 9876 10121 9904 10152
rect 10962 10140 10968 10152
rect 11020 10140 11026 10192
rect 11422 10140 11428 10192
rect 11480 10180 11486 10192
rect 11480 10152 11928 10180
rect 11480 10140 11486 10152
rect 11900 10124 11928 10152
rect 12342 10140 12348 10192
rect 12400 10180 12406 10192
rect 15470 10180 15476 10192
rect 12400 10152 13032 10180
rect 12400 10140 12406 10152
rect 9677 10115 9735 10121
rect 9677 10112 9689 10115
rect 9456 10084 9689 10112
rect 9456 10072 9462 10084
rect 9677 10081 9689 10084
rect 9723 10081 9735 10115
rect 9677 10075 9735 10081
rect 9861 10115 9919 10121
rect 9861 10081 9873 10115
rect 9907 10081 9919 10115
rect 9861 10075 9919 10081
rect 9950 10072 9956 10124
rect 10008 10072 10014 10124
rect 10045 10115 10103 10121
rect 10045 10081 10057 10115
rect 10091 10112 10103 10115
rect 10134 10112 10140 10124
rect 10091 10084 10140 10112
rect 10091 10081 10103 10084
rect 10045 10075 10103 10081
rect 9232 10044 9260 10072
rect 8496 10016 9260 10044
rect 7653 10007 7711 10013
rect 3602 9976 3608 9988
rect 2547 9948 3608 9976
rect 2547 9945 2559 9948
rect 2501 9939 2559 9945
rect 3602 9936 3608 9948
rect 3660 9936 3666 9988
rect 5534 9936 5540 9988
rect 5592 9976 5598 9988
rect 6273 9979 6331 9985
rect 6273 9976 6285 9979
rect 5592 9948 6285 9976
rect 5592 9936 5598 9948
rect 6273 9945 6285 9948
rect 6319 9945 6331 9979
rect 6273 9939 6331 9945
rect 7837 9979 7895 9985
rect 7837 9945 7849 9979
rect 7883 9976 7895 9979
rect 10060 9976 10088 10075
rect 10134 10072 10140 10084
rect 10192 10072 10198 10124
rect 10502 10072 10508 10124
rect 10560 10072 10566 10124
rect 11698 10072 11704 10124
rect 11756 10112 11762 10124
rect 11793 10115 11851 10121
rect 11793 10112 11805 10115
rect 11756 10084 11805 10112
rect 11756 10072 11762 10084
rect 11793 10081 11805 10084
rect 11839 10081 11851 10115
rect 11793 10075 11851 10081
rect 11882 10072 11888 10124
rect 11940 10112 11946 10124
rect 13004 10121 13032 10152
rect 13096 10152 13400 10180
rect 13096 10121 13124 10152
rect 13372 10124 13400 10152
rect 13724 10152 15476 10180
rect 12253 10115 12311 10121
rect 12253 10112 12265 10115
rect 11940 10084 12265 10112
rect 11940 10072 11946 10084
rect 12253 10081 12265 10084
rect 12299 10081 12311 10115
rect 12253 10075 12311 10081
rect 12989 10115 13047 10121
rect 12989 10081 13001 10115
rect 13035 10081 13047 10115
rect 12989 10075 13047 10081
rect 13081 10115 13139 10121
rect 13081 10081 13093 10115
rect 13127 10081 13139 10115
rect 13081 10075 13139 10081
rect 13265 10115 13323 10121
rect 13265 10081 13277 10115
rect 13311 10081 13323 10115
rect 13265 10075 13323 10081
rect 10152 10016 12112 10044
rect 10152 9988 10180 10016
rect 7883 9948 10088 9976
rect 7883 9945 7895 9948
rect 7837 9939 7895 9945
rect 2130 9868 2136 9920
rect 2188 9908 2194 9920
rect 2225 9911 2283 9917
rect 2225 9908 2237 9911
rect 2188 9880 2237 9908
rect 2188 9868 2194 9880
rect 2225 9877 2237 9880
rect 2271 9877 2283 9911
rect 2225 9871 2283 9877
rect 2958 9868 2964 9920
rect 3016 9868 3022 9920
rect 3418 9868 3424 9920
rect 3476 9868 3482 9920
rect 4246 9868 4252 9920
rect 4304 9908 4310 9920
rect 4341 9911 4399 9917
rect 4341 9908 4353 9911
rect 4304 9880 4353 9908
rect 4304 9868 4310 9880
rect 4341 9877 4353 9880
rect 4387 9877 4399 9911
rect 4341 9871 4399 9877
rect 5626 9868 5632 9920
rect 5684 9908 5690 9920
rect 5813 9911 5871 9917
rect 5813 9908 5825 9911
rect 5684 9880 5825 9908
rect 5684 9868 5690 9880
rect 5813 9877 5825 9880
rect 5859 9877 5871 9911
rect 5813 9871 5871 9877
rect 7190 9868 7196 9920
rect 7248 9868 7254 9920
rect 7745 9911 7803 9917
rect 7745 9877 7757 9911
rect 7791 9908 7803 9911
rect 8018 9908 8024 9920
rect 7791 9880 8024 9908
rect 7791 9877 7803 9880
rect 7745 9871 7803 9877
rect 8018 9868 8024 9880
rect 8076 9868 8082 9920
rect 8220 9917 8248 9948
rect 10134 9936 10140 9988
rect 10192 9936 10198 9988
rect 10321 9979 10379 9985
rect 10321 9945 10333 9979
rect 10367 9976 10379 9979
rect 11974 9976 11980 9988
rect 10367 9948 11980 9976
rect 10367 9945 10379 9948
rect 10321 9939 10379 9945
rect 11974 9936 11980 9948
rect 12032 9936 12038 9988
rect 12084 9976 12112 10016
rect 12894 10004 12900 10056
rect 12952 10044 12958 10056
rect 13173 10047 13231 10053
rect 13173 10044 13185 10047
rect 12952 10016 13185 10044
rect 12952 10004 12958 10016
rect 13173 10013 13185 10016
rect 13219 10013 13231 10047
rect 13280 10044 13308 10075
rect 13354 10072 13360 10124
rect 13412 10072 13418 10124
rect 13630 10072 13636 10124
rect 13688 10110 13694 10124
rect 13724 10110 13752 10152
rect 15470 10140 15476 10152
rect 15528 10140 15534 10192
rect 13688 10082 13752 10110
rect 13688 10072 13694 10082
rect 14550 10072 14556 10124
rect 14608 10112 14614 10124
rect 14645 10115 14703 10121
rect 14645 10112 14657 10115
rect 14608 10084 14657 10112
rect 14608 10072 14614 10084
rect 14645 10081 14657 10084
rect 14691 10081 14703 10115
rect 14645 10075 14703 10081
rect 15286 10072 15292 10124
rect 15344 10072 15350 10124
rect 15580 10122 15608 10220
rect 15838 10208 15844 10260
rect 15896 10248 15902 10260
rect 16209 10251 16267 10257
rect 16209 10248 16221 10251
rect 15896 10220 16221 10248
rect 15896 10208 15902 10220
rect 16209 10217 16221 10220
rect 16255 10217 16267 10251
rect 17954 10248 17960 10260
rect 16209 10211 16267 10217
rect 16868 10220 17960 10248
rect 15746 10140 15752 10192
rect 15804 10180 15810 10192
rect 16868 10180 16896 10220
rect 17954 10208 17960 10220
rect 18012 10208 18018 10260
rect 18414 10208 18420 10260
rect 18472 10248 18478 10260
rect 19886 10248 19892 10260
rect 18472 10220 19892 10248
rect 18472 10208 18478 10220
rect 15804 10152 16896 10180
rect 17773 10183 17831 10189
rect 15804 10140 15810 10152
rect 17773 10149 17785 10183
rect 17819 10180 17831 10183
rect 19242 10180 19248 10192
rect 17819 10152 18092 10180
rect 17819 10149 17831 10152
rect 17773 10143 17831 10149
rect 15580 10121 15700 10122
rect 15580 10115 15715 10121
rect 15580 10094 15669 10115
rect 15657 10081 15669 10094
rect 15703 10081 15715 10115
rect 15657 10075 15715 10081
rect 15933 10115 15991 10121
rect 15933 10081 15945 10115
rect 15979 10081 15991 10115
rect 15933 10075 15991 10081
rect 13446 10044 13452 10056
rect 13280 10016 13452 10044
rect 13173 10007 13231 10013
rect 13446 10004 13452 10016
rect 13504 10044 13510 10056
rect 13814 10044 13820 10056
rect 13504 10016 13820 10044
rect 13504 10004 13510 10016
rect 13814 10004 13820 10016
rect 13872 10004 13878 10056
rect 14737 10047 14795 10053
rect 14737 10013 14749 10047
rect 14783 10044 14795 10047
rect 14826 10044 14832 10056
rect 14783 10016 14832 10044
rect 14783 10013 14795 10016
rect 14737 10007 14795 10013
rect 14826 10004 14832 10016
rect 14884 10004 14890 10056
rect 14918 10004 14924 10056
rect 14976 10044 14982 10056
rect 15304 10044 15332 10072
rect 15948 10044 15976 10075
rect 16114 10072 16120 10124
rect 16172 10072 16178 10124
rect 16298 10072 16304 10124
rect 16356 10072 16362 10124
rect 18064 10121 18092 10152
rect 19168 10152 19248 10180
rect 17681 10115 17739 10121
rect 17681 10081 17693 10115
rect 17727 10081 17739 10115
rect 17681 10075 17739 10081
rect 17865 10115 17923 10121
rect 17865 10081 17877 10115
rect 17911 10081 17923 10115
rect 17865 10075 17923 10081
rect 18049 10115 18107 10121
rect 18049 10081 18061 10115
rect 18095 10081 18107 10115
rect 18049 10075 18107 10081
rect 18141 10115 18199 10121
rect 18141 10081 18153 10115
rect 18187 10112 18199 10115
rect 18230 10112 18236 10124
rect 18187 10084 18236 10112
rect 18187 10081 18199 10084
rect 18141 10075 18199 10081
rect 14976 10016 15976 10044
rect 16132 10044 16160 10072
rect 17696 10044 17724 10075
rect 16132 10016 17724 10044
rect 17880 10044 17908 10075
rect 18230 10072 18236 10084
rect 18288 10072 18294 10124
rect 18322 10072 18328 10124
rect 18380 10072 18386 10124
rect 19168 10121 19196 10152
rect 19242 10140 19248 10152
rect 19300 10140 19306 10192
rect 19352 10121 19380 10220
rect 19886 10208 19892 10220
rect 19944 10208 19950 10260
rect 20257 10251 20315 10257
rect 20257 10217 20269 10251
rect 20303 10248 20315 10251
rect 21266 10248 21272 10260
rect 20303 10220 21272 10248
rect 20303 10217 20315 10220
rect 20257 10211 20315 10217
rect 21266 10208 21272 10220
rect 21324 10208 21330 10260
rect 21450 10208 21456 10260
rect 21508 10208 21514 10260
rect 20070 10140 20076 10192
rect 20128 10180 20134 10192
rect 21542 10180 21548 10192
rect 20128 10152 21548 10180
rect 20128 10140 20134 10152
rect 21542 10140 21548 10152
rect 21600 10140 21606 10192
rect 22646 10180 22652 10192
rect 22480 10152 22652 10180
rect 19153 10115 19211 10121
rect 19153 10081 19165 10115
rect 19199 10081 19211 10115
rect 19153 10075 19211 10081
rect 19337 10115 19395 10121
rect 19337 10081 19349 10115
rect 19383 10081 19395 10115
rect 19337 10075 19395 10081
rect 19610 10072 19616 10124
rect 19668 10072 19674 10124
rect 19978 10072 19984 10124
rect 20036 10112 20042 10124
rect 20530 10112 20536 10124
rect 20036 10084 20536 10112
rect 20036 10072 20042 10084
rect 20530 10072 20536 10084
rect 20588 10072 20594 10124
rect 20625 10115 20683 10121
rect 20625 10081 20637 10115
rect 20671 10112 20683 10115
rect 20714 10112 20720 10124
rect 20671 10084 20720 10112
rect 20671 10081 20683 10084
rect 20625 10075 20683 10081
rect 20714 10072 20720 10084
rect 20772 10112 20778 10124
rect 22480 10121 22508 10152
rect 22646 10140 22652 10152
rect 22704 10180 22710 10192
rect 22922 10180 22928 10192
rect 22704 10152 22928 10180
rect 22704 10140 22710 10152
rect 22922 10140 22928 10152
rect 22980 10140 22986 10192
rect 20901 10115 20959 10121
rect 20901 10112 20913 10115
rect 20772 10084 20913 10112
rect 20772 10072 20778 10084
rect 20901 10081 20913 10084
rect 20947 10112 20959 10115
rect 21637 10115 21695 10121
rect 21637 10112 21649 10115
rect 20947 10084 21649 10112
rect 20947 10081 20959 10084
rect 20901 10075 20959 10081
rect 21637 10081 21649 10084
rect 21683 10081 21695 10115
rect 21637 10075 21695 10081
rect 22465 10115 22523 10121
rect 22465 10081 22477 10115
rect 22511 10081 22523 10115
rect 22465 10075 22523 10081
rect 22741 10115 22799 10121
rect 22741 10081 22753 10115
rect 22787 10112 22799 10115
rect 23017 10115 23075 10121
rect 23017 10112 23029 10115
rect 22787 10084 23029 10112
rect 22787 10081 22799 10084
rect 22741 10075 22799 10081
rect 23017 10081 23029 10084
rect 23063 10112 23075 10115
rect 23198 10112 23204 10124
rect 23063 10084 23204 10112
rect 23063 10081 23075 10084
rect 23017 10075 23075 10081
rect 23198 10072 23204 10084
rect 23256 10072 23262 10124
rect 19061 10047 19119 10053
rect 19061 10044 19073 10047
rect 17880 10016 18184 10044
rect 14976 10004 14982 10016
rect 12084 9948 14228 9976
rect 8205 9911 8263 9917
rect 8205 9877 8217 9911
rect 8251 9877 8263 9911
rect 8205 9871 8263 9877
rect 8389 9911 8447 9917
rect 8389 9877 8401 9911
rect 8435 9908 8447 9911
rect 8570 9908 8576 9920
rect 8435 9880 8576 9908
rect 8435 9877 8447 9880
rect 8389 9871 8447 9877
rect 8570 9868 8576 9880
rect 8628 9868 8634 9920
rect 9122 9868 9128 9920
rect 9180 9868 9186 9920
rect 9398 9868 9404 9920
rect 9456 9868 9462 9920
rect 9582 9868 9588 9920
rect 9640 9908 9646 9920
rect 10502 9908 10508 9920
rect 9640 9880 10508 9908
rect 9640 9868 9646 9880
rect 10502 9868 10508 9880
rect 10560 9868 10566 9920
rect 10689 9911 10747 9917
rect 10689 9877 10701 9911
rect 10735 9908 10747 9911
rect 11698 9908 11704 9920
rect 10735 9880 11704 9908
rect 10735 9877 10747 9880
rect 10689 9871 10747 9877
rect 11698 9868 11704 9880
rect 11756 9868 11762 9920
rect 12066 9868 12072 9920
rect 12124 9868 12130 9920
rect 12526 9868 12532 9920
rect 12584 9908 12590 9920
rect 12802 9908 12808 9920
rect 12584 9880 12808 9908
rect 12584 9868 12590 9880
rect 12802 9868 12808 9880
rect 12860 9868 12866 9920
rect 14200 9908 14228 9948
rect 15010 9936 15016 9988
rect 15068 9936 15074 9988
rect 15286 9936 15292 9988
rect 15344 9976 15350 9988
rect 15841 9979 15899 9985
rect 15841 9976 15853 9979
rect 15344 9948 15853 9976
rect 15344 9936 15350 9948
rect 15841 9945 15853 9948
rect 15887 9945 15899 9979
rect 15948 9976 15976 10016
rect 16390 9976 16396 9988
rect 15948 9948 16396 9976
rect 15841 9939 15899 9945
rect 16390 9936 16396 9948
rect 16448 9936 16454 9988
rect 17494 9936 17500 9988
rect 17552 9976 17558 9988
rect 17880 9976 17908 10016
rect 18156 9988 18184 10016
rect 18340 10016 19073 10044
rect 17552 9948 17908 9976
rect 17552 9936 17558 9948
rect 18138 9936 18144 9988
rect 18196 9936 18202 9988
rect 18340 9985 18368 10016
rect 19061 10013 19073 10016
rect 19107 10013 19119 10047
rect 19061 10007 19119 10013
rect 19245 10047 19303 10053
rect 19245 10013 19257 10047
rect 19291 10013 19303 10047
rect 19245 10007 19303 10013
rect 19521 10047 19579 10053
rect 19521 10013 19533 10047
rect 19567 10044 19579 10047
rect 20254 10044 20260 10056
rect 19567 10016 20260 10044
rect 19567 10013 19579 10016
rect 19521 10007 19579 10013
rect 18325 9979 18383 9985
rect 18325 9945 18337 9979
rect 18371 9945 18383 9979
rect 19260 9976 19288 10007
rect 20254 10004 20260 10016
rect 20312 10004 20318 10056
rect 21266 10004 21272 10056
rect 21324 10004 21330 10056
rect 19797 9979 19855 9985
rect 19797 9976 19809 9979
rect 19260 9948 19809 9976
rect 18325 9939 18383 9945
rect 19797 9945 19809 9948
rect 19843 9976 19855 9979
rect 20162 9976 20168 9988
rect 19843 9948 20168 9976
rect 19843 9945 19855 9948
rect 19797 9939 19855 9945
rect 20162 9936 20168 9948
rect 20220 9936 20226 9988
rect 20898 9976 20904 9988
rect 20272 9948 20904 9976
rect 19058 9908 19064 9920
rect 14200 9880 19064 9908
rect 19058 9868 19064 9880
rect 19116 9908 19122 9920
rect 19426 9908 19432 9920
rect 19116 9880 19432 9908
rect 19116 9868 19122 9880
rect 19426 9868 19432 9880
rect 19484 9868 19490 9920
rect 19978 9868 19984 9920
rect 20036 9908 20042 9920
rect 20272 9917 20300 9948
rect 20898 9936 20904 9948
rect 20956 9936 20962 9988
rect 21450 9936 21456 9988
rect 21508 9976 21514 9988
rect 21508 9948 22324 9976
rect 21508 9936 21514 9948
rect 20073 9911 20131 9917
rect 20073 9908 20085 9911
rect 20036 9880 20085 9908
rect 20036 9868 20042 9880
rect 20073 9877 20085 9880
rect 20119 9877 20131 9911
rect 20073 9871 20131 9877
rect 20257 9911 20315 9917
rect 20257 9877 20269 9911
rect 20303 9877 20315 9911
rect 20257 9871 20315 9877
rect 20346 9868 20352 9920
rect 20404 9908 20410 9920
rect 20717 9911 20775 9917
rect 20717 9908 20729 9911
rect 20404 9880 20729 9908
rect 20404 9868 20410 9880
rect 20717 9877 20729 9880
rect 20763 9877 20775 9911
rect 20717 9871 20775 9877
rect 21542 9868 21548 9920
rect 21600 9908 21606 9920
rect 22296 9917 22324 9948
rect 22462 9936 22468 9988
rect 22520 9976 22526 9988
rect 22833 9979 22891 9985
rect 22833 9976 22845 9979
rect 22520 9948 22845 9976
rect 22520 9936 22526 9948
rect 22833 9945 22845 9948
rect 22879 9945 22891 9979
rect 22833 9939 22891 9945
rect 21637 9911 21695 9917
rect 21637 9908 21649 9911
rect 21600 9880 21649 9908
rect 21600 9868 21606 9880
rect 21637 9877 21649 9880
rect 21683 9877 21695 9911
rect 21637 9871 21695 9877
rect 22281 9911 22339 9917
rect 22281 9877 22293 9911
rect 22327 9877 22339 9911
rect 22281 9871 22339 9877
rect 22649 9911 22707 9917
rect 22649 9877 22661 9911
rect 22695 9908 22707 9911
rect 22738 9908 22744 9920
rect 22695 9880 22744 9908
rect 22695 9877 22707 9880
rect 22649 9871 22707 9877
rect 22738 9868 22744 9880
rect 22796 9868 22802 9920
rect 552 9818 23368 9840
rect 552 9766 1366 9818
rect 1418 9766 1430 9818
rect 1482 9766 1494 9818
rect 1546 9766 1558 9818
rect 1610 9766 1622 9818
rect 1674 9766 1686 9818
rect 1738 9766 7366 9818
rect 7418 9766 7430 9818
rect 7482 9766 7494 9818
rect 7546 9766 7558 9818
rect 7610 9766 7622 9818
rect 7674 9766 7686 9818
rect 7738 9766 13366 9818
rect 13418 9766 13430 9818
rect 13482 9766 13494 9818
rect 13546 9766 13558 9818
rect 13610 9766 13622 9818
rect 13674 9766 13686 9818
rect 13738 9766 19366 9818
rect 19418 9766 19430 9818
rect 19482 9766 19494 9818
rect 19546 9766 19558 9818
rect 19610 9766 19622 9818
rect 19674 9766 19686 9818
rect 19738 9766 23368 9818
rect 552 9744 23368 9766
rect 1946 9704 1952 9716
rect 1688 9676 1952 9704
rect 1688 9648 1716 9676
rect 1946 9664 1952 9676
rect 2004 9704 2010 9716
rect 2363 9707 2421 9713
rect 2363 9704 2375 9707
rect 2004 9676 2375 9704
rect 2004 9664 2010 9676
rect 2363 9673 2375 9676
rect 2409 9673 2421 9707
rect 4798 9704 4804 9716
rect 2363 9667 2421 9673
rect 4172 9676 4804 9704
rect 1670 9596 1676 9648
rect 1728 9596 1734 9648
rect 4062 9636 4068 9648
rect 3715 9608 4068 9636
rect 3418 9528 3424 9580
rect 3476 9568 3482 9580
rect 3715 9568 3743 9608
rect 4062 9596 4068 9608
rect 4120 9596 4126 9648
rect 4172 9568 4200 9676
rect 4798 9664 4804 9676
rect 4856 9664 4862 9716
rect 7282 9704 7288 9716
rect 6932 9676 7288 9704
rect 4246 9596 4252 9648
rect 4304 9636 4310 9648
rect 6365 9639 6423 9645
rect 4304 9608 5120 9636
rect 4304 9596 4310 9608
rect 3476 9540 3743 9568
rect 3476 9528 3482 9540
rect 566 9460 572 9512
rect 624 9500 630 9512
rect 1029 9503 1087 9509
rect 1029 9500 1041 9503
rect 624 9472 1041 9500
rect 624 9460 630 9472
rect 1029 9469 1041 9472
rect 1075 9469 1087 9503
rect 1029 9463 1087 9469
rect 1044 9432 1072 9463
rect 1394 9460 1400 9512
rect 1452 9460 1458 9512
rect 2133 9503 2191 9509
rect 2133 9469 2145 9503
rect 2179 9469 2191 9503
rect 2133 9463 2191 9469
rect 2148 9432 2176 9463
rect 2590 9460 2596 9512
rect 2648 9500 2654 9512
rect 3513 9503 3571 9509
rect 3513 9500 3525 9503
rect 2648 9472 3525 9500
rect 2648 9460 2654 9472
rect 3513 9469 3525 9472
rect 3559 9469 3571 9503
rect 3513 9463 3571 9469
rect 3602 9460 3608 9512
rect 3660 9460 3666 9512
rect 3715 9509 3743 9540
rect 3804 9540 4200 9568
rect 3697 9503 3755 9509
rect 3697 9469 3709 9503
rect 3743 9469 3755 9503
rect 3697 9463 3755 9469
rect 1044 9404 2176 9432
rect 2038 9324 2044 9376
rect 2096 9324 2102 9376
rect 3050 9324 3056 9376
rect 3108 9364 3114 9376
rect 3237 9367 3295 9373
rect 3237 9364 3249 9367
rect 3108 9336 3249 9364
rect 3108 9324 3114 9336
rect 3237 9333 3249 9336
rect 3283 9333 3295 9367
rect 3237 9327 3295 9333
rect 3326 9324 3332 9376
rect 3384 9364 3390 9376
rect 3804 9364 3832 9540
rect 4338 9528 4344 9580
rect 4396 9528 4402 9580
rect 4985 9571 5043 9577
rect 4985 9568 4997 9571
rect 4448 9540 4997 9568
rect 3881 9503 3939 9509
rect 3881 9469 3893 9503
rect 3927 9469 3939 9503
rect 3881 9463 3939 9469
rect 3384 9336 3832 9364
rect 3896 9364 3924 9463
rect 3970 9460 3976 9512
rect 4028 9460 4034 9512
rect 4154 9460 4160 9512
rect 4212 9460 4218 9512
rect 4448 9509 4476 9540
rect 4985 9537 4997 9540
rect 5031 9537 5043 9571
rect 4985 9531 5043 9537
rect 5092 9509 5120 9608
rect 6365 9605 6377 9639
rect 6411 9636 6423 9639
rect 6932 9636 6960 9676
rect 7282 9664 7288 9676
rect 7340 9664 7346 9716
rect 7558 9664 7564 9716
rect 7616 9704 7622 9716
rect 8294 9704 8300 9716
rect 7616 9676 8300 9704
rect 7616 9664 7622 9676
rect 8294 9664 8300 9676
rect 8352 9664 8358 9716
rect 8481 9707 8539 9713
rect 8481 9673 8493 9707
rect 8527 9704 8539 9707
rect 8754 9704 8760 9716
rect 8527 9676 8760 9704
rect 8527 9673 8539 9676
rect 8481 9667 8539 9673
rect 8754 9664 8760 9676
rect 8812 9664 8818 9716
rect 8846 9664 8852 9716
rect 8904 9704 8910 9716
rect 9398 9704 9404 9716
rect 8904 9676 9404 9704
rect 8904 9664 8910 9676
rect 9398 9664 9404 9676
rect 9456 9664 9462 9716
rect 12066 9704 12072 9716
rect 9600 9676 12072 9704
rect 6411 9608 6960 9636
rect 7009 9639 7067 9645
rect 6411 9605 6423 9608
rect 6365 9599 6423 9605
rect 7009 9605 7021 9639
rect 7055 9636 7067 9639
rect 8113 9639 8171 9645
rect 8113 9636 8125 9639
rect 7055 9608 8125 9636
rect 7055 9605 7067 9608
rect 7009 9599 7067 9605
rect 8113 9605 8125 9608
rect 8159 9605 8171 9639
rect 8113 9599 8171 9605
rect 8386 9596 8392 9648
rect 8444 9636 8450 9648
rect 9600 9636 9628 9676
rect 12066 9664 12072 9676
rect 12124 9664 12130 9716
rect 12710 9704 12716 9716
rect 12360 9676 12716 9704
rect 8444 9608 9628 9636
rect 9861 9639 9919 9645
rect 8444 9596 8450 9608
rect 9861 9605 9873 9639
rect 9907 9605 9919 9639
rect 9861 9599 9919 9605
rect 6086 9568 6092 9580
rect 5736 9540 6092 9568
rect 4433 9503 4491 9509
rect 4433 9469 4445 9503
rect 4479 9469 4491 9503
rect 4433 9463 4491 9469
rect 4893 9503 4951 9509
rect 4893 9469 4905 9503
rect 4939 9469 4951 9503
rect 4893 9463 4951 9469
rect 5077 9503 5135 9509
rect 5077 9469 5089 9503
rect 5123 9469 5135 9503
rect 5077 9463 5135 9469
rect 5445 9503 5503 9509
rect 5445 9469 5457 9503
rect 5491 9500 5503 9503
rect 5534 9500 5540 9512
rect 5491 9472 5540 9500
rect 5491 9469 5503 9472
rect 5445 9463 5503 9469
rect 4062 9392 4068 9444
rect 4120 9432 4126 9444
rect 4908 9432 4936 9463
rect 5534 9460 5540 9472
rect 5592 9460 5598 9512
rect 5626 9460 5632 9512
rect 5684 9460 5690 9512
rect 5736 9509 5764 9540
rect 6086 9528 6092 9540
rect 6144 9528 6150 9580
rect 6917 9571 6975 9577
rect 6380 9540 6868 9568
rect 6380 9512 6408 9540
rect 5721 9503 5779 9509
rect 5721 9469 5733 9503
rect 5767 9469 5779 9503
rect 5721 9463 5779 9469
rect 5997 9503 6055 9509
rect 5997 9469 6009 9503
rect 6043 9500 6055 9503
rect 6270 9500 6276 9512
rect 6043 9472 6276 9500
rect 6043 9469 6055 9472
rect 5997 9463 6055 9469
rect 6270 9460 6276 9472
rect 6328 9460 6334 9512
rect 6362 9460 6368 9512
rect 6420 9460 6426 9512
rect 6546 9460 6552 9512
rect 6604 9500 6610 9512
rect 6840 9509 6868 9540
rect 6917 9537 6929 9571
rect 6963 9568 6975 9571
rect 7190 9568 7196 9580
rect 6963 9540 7196 9568
rect 6963 9537 6975 9540
rect 6917 9531 6975 9537
rect 7190 9528 7196 9540
rect 7248 9528 7254 9580
rect 8202 9568 8208 9580
rect 7300 9540 7696 9568
rect 6641 9503 6699 9509
rect 6641 9500 6653 9503
rect 6604 9472 6653 9500
rect 6604 9460 6610 9472
rect 6641 9469 6653 9472
rect 6687 9469 6699 9503
rect 6641 9463 6699 9469
rect 6825 9503 6883 9509
rect 6825 9469 6837 9503
rect 6871 9469 6883 9503
rect 7300 9500 7328 9540
rect 6825 9463 6883 9469
rect 7116 9472 7328 9500
rect 7436 9503 7494 9509
rect 7116 9444 7144 9472
rect 7436 9469 7448 9503
rect 7482 9500 7494 9503
rect 7558 9500 7564 9512
rect 7482 9472 7564 9500
rect 7482 9469 7494 9472
rect 7436 9463 7494 9469
rect 7558 9460 7564 9472
rect 7616 9460 7622 9512
rect 7668 9509 7696 9540
rect 7944 9540 8208 9568
rect 7944 9509 7972 9540
rect 8202 9528 8208 9540
rect 8260 9528 8266 9580
rect 8478 9528 8484 9580
rect 8536 9568 8542 9580
rect 8662 9568 8668 9580
rect 8536 9540 8668 9568
rect 8536 9528 8542 9540
rect 8662 9528 8668 9540
rect 8720 9568 8726 9580
rect 8849 9571 8907 9577
rect 8849 9568 8861 9571
rect 8720 9540 8861 9568
rect 8720 9528 8726 9540
rect 8849 9537 8861 9540
rect 8895 9537 8907 9571
rect 8849 9531 8907 9537
rect 8938 9528 8944 9580
rect 8996 9528 9002 9580
rect 9033 9571 9091 9577
rect 9033 9537 9045 9571
rect 9079 9568 9091 9571
rect 9398 9568 9404 9580
rect 9079 9540 9404 9568
rect 9079 9537 9091 9540
rect 9033 9531 9091 9537
rect 9398 9528 9404 9540
rect 9456 9568 9462 9580
rect 9876 9568 9904 9599
rect 10778 9596 10784 9648
rect 10836 9636 10842 9648
rect 12360 9636 12388 9676
rect 12710 9664 12716 9676
rect 12768 9704 12774 9716
rect 14642 9704 14648 9716
rect 12768 9676 12848 9704
rect 12768 9664 12774 9676
rect 10836 9608 12388 9636
rect 12437 9639 12495 9645
rect 10836 9596 10842 9608
rect 9456 9540 9904 9568
rect 10612 9540 11468 9568
rect 9456 9528 9462 9540
rect 7653 9503 7711 9509
rect 7653 9469 7665 9503
rect 7699 9469 7711 9503
rect 7653 9463 7711 9469
rect 7929 9503 7987 9509
rect 7929 9469 7941 9503
rect 7975 9469 7987 9503
rect 7929 9463 7987 9469
rect 8018 9460 8024 9512
rect 8076 9500 8082 9512
rect 8389 9503 8447 9509
rect 8389 9500 8401 9503
rect 8076 9472 8401 9500
rect 8076 9460 8082 9472
rect 8389 9469 8401 9472
rect 8435 9469 8447 9503
rect 8389 9463 8447 9469
rect 8570 9460 8576 9512
rect 8628 9460 8634 9512
rect 9125 9503 9183 9509
rect 9125 9500 9137 9503
rect 8956 9472 9137 9500
rect 7098 9432 7104 9444
rect 4120 9404 4936 9432
rect 5184 9404 7104 9432
rect 4120 9392 4126 9404
rect 3970 9364 3976 9376
rect 3896 9336 3976 9364
rect 3384 9324 3390 9336
rect 3970 9324 3976 9336
rect 4028 9324 4034 9376
rect 4801 9367 4859 9373
rect 4801 9333 4813 9367
rect 4847 9364 4859 9367
rect 5184 9364 5212 9404
rect 7098 9392 7104 9404
rect 7156 9392 7162 9444
rect 7282 9392 7288 9444
rect 7340 9432 7346 9444
rect 7745 9435 7803 9441
rect 7745 9432 7757 9435
rect 7340 9404 7757 9432
rect 7340 9392 7346 9404
rect 7745 9401 7757 9404
rect 7791 9401 7803 9435
rect 7745 9395 7803 9401
rect 8662 9392 8668 9444
rect 8720 9432 8726 9444
rect 8956 9432 8984 9472
rect 9125 9469 9137 9472
rect 9171 9469 9183 9503
rect 9125 9463 9183 9469
rect 9585 9503 9643 9509
rect 9585 9469 9597 9503
rect 9631 9469 9643 9503
rect 9585 9463 9643 9469
rect 8720 9404 8984 9432
rect 8720 9392 8726 9404
rect 9030 9392 9036 9444
rect 9088 9432 9094 9444
rect 9600 9432 9628 9463
rect 9674 9460 9680 9512
rect 9732 9460 9738 9512
rect 10612 9509 10640 9540
rect 11440 9512 11468 9540
rect 11606 9528 11612 9580
rect 11664 9528 11670 9580
rect 9953 9503 10011 9509
rect 9953 9469 9965 9503
rect 9999 9500 10011 9503
rect 10413 9503 10471 9509
rect 10413 9500 10425 9503
rect 9999 9472 10425 9500
rect 9999 9469 10011 9472
rect 9953 9463 10011 9469
rect 10413 9469 10425 9472
rect 10459 9469 10471 9503
rect 10413 9463 10471 9469
rect 10597 9503 10655 9509
rect 10597 9469 10609 9503
rect 10643 9469 10655 9503
rect 10597 9463 10655 9469
rect 10686 9460 10692 9512
rect 10744 9460 10750 9512
rect 10781 9503 10839 9509
rect 10781 9469 10793 9503
rect 10827 9500 10839 9503
rect 10870 9500 10876 9512
rect 10827 9472 10876 9500
rect 10827 9469 10839 9472
rect 10781 9463 10839 9469
rect 10870 9460 10876 9472
rect 10928 9460 10934 9512
rect 10965 9503 11023 9509
rect 10965 9469 10977 9503
rect 11011 9500 11023 9503
rect 11054 9500 11060 9512
rect 11011 9472 11060 9500
rect 11011 9469 11023 9472
rect 10965 9463 11023 9469
rect 11054 9460 11060 9472
rect 11112 9460 11118 9512
rect 11146 9460 11152 9512
rect 11204 9460 11210 9512
rect 11241 9503 11299 9509
rect 11241 9469 11253 9503
rect 11287 9500 11299 9503
rect 11330 9500 11336 9512
rect 11287 9472 11336 9500
rect 11287 9469 11299 9472
rect 11241 9463 11299 9469
rect 11330 9460 11336 9472
rect 11388 9460 11394 9512
rect 11422 9460 11428 9512
rect 11480 9460 11486 9512
rect 11808 9509 11836 9608
rect 12437 9605 12449 9639
rect 12483 9636 12495 9639
rect 12483 9608 12572 9636
rect 12483 9605 12495 9608
rect 12437 9599 12495 9605
rect 11977 9571 12035 9577
rect 11977 9537 11989 9571
rect 12023 9568 12035 9571
rect 12250 9568 12256 9580
rect 12023 9540 12256 9568
rect 12023 9537 12035 9540
rect 11977 9531 12035 9537
rect 12250 9528 12256 9540
rect 12308 9528 12314 9580
rect 12544 9509 12572 9608
rect 12820 9577 12848 9676
rect 13740 9676 14648 9704
rect 13078 9596 13084 9648
rect 13136 9636 13142 9648
rect 13262 9636 13268 9648
rect 13136 9608 13268 9636
rect 13136 9596 13142 9608
rect 13262 9596 13268 9608
rect 13320 9596 13326 9648
rect 12805 9571 12863 9577
rect 12805 9537 12817 9571
rect 12851 9537 12863 9571
rect 12805 9531 12863 9537
rect 12894 9528 12900 9580
rect 12952 9568 12958 9580
rect 13633 9571 13691 9577
rect 12952 9540 13584 9568
rect 12952 9528 12958 9540
rect 11517 9503 11575 9509
rect 11517 9469 11529 9503
rect 11563 9469 11575 9503
rect 11517 9463 11575 9469
rect 11804 9503 11862 9509
rect 11804 9469 11816 9503
rect 11850 9469 11862 9503
rect 11804 9463 11862 9469
rect 12529 9503 12587 9509
rect 12529 9469 12541 9503
rect 12575 9469 12587 9503
rect 12529 9463 12587 9469
rect 10042 9432 10048 9444
rect 9088 9404 9444 9432
rect 9600 9404 10048 9432
rect 9088 9392 9094 9404
rect 4847 9336 5212 9364
rect 4847 9333 4859 9336
rect 4801 9327 4859 9333
rect 5258 9324 5264 9376
rect 5316 9324 5322 9376
rect 6825 9367 6883 9373
rect 6825 9333 6837 9367
rect 6871 9364 6883 9367
rect 7377 9367 7435 9373
rect 7377 9364 7389 9367
rect 6871 9336 7389 9364
rect 6871 9333 6883 9336
rect 6825 9327 6883 9333
rect 7377 9333 7389 9336
rect 7423 9333 7435 9367
rect 7377 9327 7435 9333
rect 7561 9367 7619 9373
rect 7561 9333 7573 9367
rect 7607 9364 7619 9367
rect 8202 9364 8208 9376
rect 7607 9336 8208 9364
rect 7607 9333 7619 9336
rect 7561 9327 7619 9333
rect 8202 9324 8208 9336
rect 8260 9324 8266 9376
rect 8754 9324 8760 9376
rect 8812 9364 8818 9376
rect 9416 9373 9444 9404
rect 10042 9392 10048 9404
rect 10100 9392 10106 9444
rect 10137 9435 10195 9441
rect 10137 9401 10149 9435
rect 10183 9401 10195 9435
rect 10137 9395 10195 9401
rect 9309 9367 9367 9373
rect 9309 9364 9321 9367
rect 8812 9336 9321 9364
rect 8812 9324 8818 9336
rect 9309 9333 9321 9336
rect 9355 9333 9367 9367
rect 9309 9327 9367 9333
rect 9401 9367 9459 9373
rect 9401 9333 9413 9367
rect 9447 9333 9459 9367
rect 10152 9364 10180 9395
rect 10318 9392 10324 9444
rect 10376 9392 10382 9444
rect 11072 9432 11100 9460
rect 11532 9432 11560 9463
rect 12710 9460 12716 9512
rect 12768 9460 12774 9512
rect 13081 9503 13139 9509
rect 13081 9500 13093 9503
rect 12820 9472 13093 9500
rect 12820 9444 12848 9472
rect 13081 9469 13093 9472
rect 13127 9469 13139 9503
rect 13556 9500 13584 9540
rect 13633 9537 13645 9571
rect 13679 9568 13691 9571
rect 13740 9568 13768 9676
rect 14642 9664 14648 9676
rect 14700 9704 14706 9716
rect 19886 9704 19892 9716
rect 14700 9676 19892 9704
rect 14700 9664 14706 9676
rect 19886 9664 19892 9676
rect 19944 9664 19950 9716
rect 20070 9664 20076 9716
rect 20128 9704 20134 9716
rect 20622 9704 20628 9716
rect 20128 9676 20628 9704
rect 20128 9664 20134 9676
rect 20622 9664 20628 9676
rect 20680 9664 20686 9716
rect 21726 9664 21732 9716
rect 21784 9664 21790 9716
rect 14090 9596 14096 9648
rect 14148 9636 14154 9648
rect 14734 9636 14740 9648
rect 14148 9608 14740 9636
rect 14148 9596 14154 9608
rect 14734 9596 14740 9608
rect 14792 9596 14798 9648
rect 15010 9596 15016 9648
rect 15068 9636 15074 9648
rect 16485 9639 16543 9645
rect 16485 9636 16497 9639
rect 15068 9608 16497 9636
rect 15068 9596 15074 9608
rect 16485 9605 16497 9608
rect 16531 9636 16543 9639
rect 16531 9608 17724 9636
rect 16531 9605 16543 9608
rect 16485 9599 16543 9605
rect 13679 9540 13768 9568
rect 13679 9537 13691 9540
rect 13633 9531 13691 9537
rect 15838 9528 15844 9580
rect 15896 9568 15902 9580
rect 16298 9568 16304 9580
rect 15896 9540 16304 9568
rect 15896 9528 15902 9540
rect 16298 9528 16304 9540
rect 16356 9528 16362 9580
rect 16390 9528 16396 9580
rect 16448 9528 16454 9580
rect 17497 9571 17555 9577
rect 17497 9568 17509 9571
rect 16500 9540 17509 9568
rect 13556 9472 13768 9500
rect 13081 9463 13139 9469
rect 12069 9435 12127 9441
rect 12069 9432 12081 9435
rect 11072 9404 11560 9432
rect 11624 9404 12081 9432
rect 11054 9364 11060 9376
rect 10152 9336 11060 9364
rect 9401 9327 9459 9333
rect 11054 9324 11060 9336
rect 11112 9364 11118 9376
rect 11624 9364 11652 9404
rect 12069 9401 12081 9404
rect 12115 9401 12127 9435
rect 12253 9435 12311 9441
rect 12253 9432 12265 9435
rect 12069 9395 12127 9401
rect 12176 9404 12265 9432
rect 11112 9336 11652 9364
rect 11112 9324 11118 9336
rect 11698 9324 11704 9376
rect 11756 9364 11762 9376
rect 12176 9364 12204 9404
rect 12253 9401 12265 9404
rect 12299 9401 12311 9435
rect 12253 9395 12311 9401
rect 12802 9392 12808 9444
rect 12860 9392 12866 9444
rect 13740 9432 13768 9472
rect 13814 9460 13820 9512
rect 13872 9500 13878 9512
rect 14093 9503 14151 9509
rect 14093 9500 14105 9503
rect 13872 9472 14105 9500
rect 13872 9460 13878 9472
rect 14093 9469 14105 9472
rect 14139 9469 14151 9503
rect 14093 9463 14151 9469
rect 14274 9460 14280 9512
rect 14332 9460 14338 9512
rect 14734 9460 14740 9512
rect 14792 9500 14798 9512
rect 16500 9500 16528 9540
rect 17497 9537 17509 9540
rect 17543 9537 17555 9571
rect 17497 9531 17555 9537
rect 14792 9472 16528 9500
rect 14792 9460 14798 9472
rect 16666 9460 16672 9512
rect 16724 9460 16730 9512
rect 17221 9503 17279 9509
rect 17221 9500 17233 9503
rect 16776 9472 17233 9500
rect 14642 9432 14648 9444
rect 13740 9404 14648 9432
rect 14642 9392 14648 9404
rect 14700 9392 14706 9444
rect 15654 9392 15660 9444
rect 15712 9432 15718 9444
rect 16776 9432 16804 9472
rect 17221 9469 17233 9472
rect 17267 9469 17279 9503
rect 17221 9463 17279 9469
rect 17310 9460 17316 9512
rect 17368 9460 17374 9512
rect 17586 9460 17592 9512
rect 17644 9460 17650 9512
rect 17696 9509 17724 9608
rect 19058 9596 19064 9648
rect 19116 9636 19122 9648
rect 20901 9639 20959 9645
rect 19116 9608 19334 9636
rect 19116 9596 19122 9608
rect 19306 9568 19334 9608
rect 20901 9605 20913 9639
rect 20947 9636 20959 9639
rect 20990 9636 20996 9648
rect 20947 9608 20996 9636
rect 20947 9605 20959 9608
rect 20901 9599 20959 9605
rect 19521 9571 19579 9577
rect 19521 9568 19533 9571
rect 19306 9540 19533 9568
rect 19521 9537 19533 9540
rect 19567 9537 19579 9571
rect 19521 9531 19579 9537
rect 19886 9528 19892 9580
rect 19944 9568 19950 9580
rect 20916 9568 20944 9599
rect 20990 9596 20996 9608
rect 21048 9596 21054 9648
rect 21082 9596 21088 9648
rect 21140 9636 21146 9648
rect 21542 9636 21548 9648
rect 21140 9608 21548 9636
rect 21140 9596 21146 9608
rect 21542 9596 21548 9608
rect 21600 9636 21606 9648
rect 22189 9639 22247 9645
rect 22189 9636 22201 9639
rect 21600 9608 22201 9636
rect 21600 9596 21606 9608
rect 22189 9605 22201 9608
rect 22235 9605 22247 9639
rect 22189 9599 22247 9605
rect 22833 9571 22891 9577
rect 22833 9568 22845 9571
rect 19944 9540 20944 9568
rect 22388 9540 22845 9568
rect 19944 9528 19950 9540
rect 17681 9503 17739 9509
rect 17681 9469 17693 9503
rect 17727 9469 17739 9503
rect 17681 9463 17739 9469
rect 17862 9460 17868 9512
rect 17920 9460 17926 9512
rect 19245 9503 19303 9509
rect 19245 9469 19257 9503
rect 19291 9469 19303 9503
rect 19245 9463 19303 9469
rect 15712 9404 16804 9432
rect 16853 9435 16911 9441
rect 15712 9392 15718 9404
rect 16853 9401 16865 9435
rect 16899 9432 16911 9435
rect 18230 9432 18236 9444
rect 16899 9404 18236 9432
rect 16899 9401 16911 9404
rect 16853 9395 16911 9401
rect 18230 9392 18236 9404
rect 18288 9392 18294 9444
rect 19260 9432 19288 9463
rect 19426 9460 19432 9512
rect 19484 9460 19490 9512
rect 19797 9503 19855 9509
rect 19797 9469 19809 9503
rect 19843 9494 19855 9503
rect 20070 9500 20076 9512
rect 19996 9494 20076 9500
rect 19843 9472 20076 9494
rect 19843 9469 20024 9472
rect 19797 9466 20024 9469
rect 19797 9463 19855 9466
rect 20070 9460 20076 9472
rect 20128 9460 20134 9512
rect 20346 9460 20352 9512
rect 20404 9500 20410 9512
rect 20824 9509 20852 9540
rect 20625 9503 20683 9509
rect 20625 9500 20637 9503
rect 20404 9472 20637 9500
rect 20404 9460 20410 9472
rect 20625 9469 20637 9472
rect 20671 9469 20683 9503
rect 20625 9463 20683 9469
rect 20809 9503 20867 9509
rect 20809 9469 20821 9503
rect 20855 9469 20867 9503
rect 20809 9463 20867 9469
rect 21085 9503 21143 9509
rect 21085 9469 21097 9503
rect 21131 9500 21143 9503
rect 21266 9500 21272 9512
rect 21131 9472 21272 9500
rect 21131 9469 21143 9472
rect 21085 9463 21143 9469
rect 21266 9460 21272 9472
rect 21324 9460 21330 9512
rect 22388 9509 22416 9540
rect 22833 9537 22845 9540
rect 22879 9537 22891 9571
rect 22833 9531 22891 9537
rect 21545 9503 21603 9509
rect 21545 9469 21557 9503
rect 21591 9500 21603 9503
rect 21637 9503 21695 9509
rect 21637 9500 21649 9503
rect 21591 9472 21649 9500
rect 21591 9469 21603 9472
rect 21545 9463 21603 9469
rect 21637 9469 21649 9472
rect 21683 9469 21695 9503
rect 21637 9463 21695 9469
rect 21821 9503 21879 9509
rect 21821 9469 21833 9503
rect 21867 9500 21879 9503
rect 22097 9503 22155 9509
rect 22097 9500 22109 9503
rect 21867 9472 22109 9500
rect 21867 9469 21879 9472
rect 21821 9463 21879 9469
rect 22097 9469 22109 9472
rect 22143 9500 22155 9503
rect 22373 9503 22431 9509
rect 22373 9500 22385 9503
rect 22143 9472 22385 9500
rect 22143 9469 22155 9472
rect 22097 9463 22155 9469
rect 22373 9469 22385 9472
rect 22419 9469 22431 9503
rect 22373 9463 22431 9469
rect 20364 9432 20392 9460
rect 18616 9404 19196 9432
rect 19260 9404 20392 9432
rect 21652 9432 21680 9463
rect 22462 9460 22468 9512
rect 22520 9460 22526 9512
rect 22646 9460 22652 9512
rect 22704 9460 22710 9512
rect 22741 9503 22799 9509
rect 22741 9469 22753 9503
rect 22787 9469 22799 9503
rect 22741 9463 22799 9469
rect 22557 9435 22615 9441
rect 22557 9432 22569 9435
rect 21652 9404 22569 9432
rect 11756 9336 12204 9364
rect 11756 9324 11762 9336
rect 13262 9324 13268 9376
rect 13320 9324 13326 9376
rect 13998 9324 14004 9376
rect 14056 9324 14062 9376
rect 14185 9367 14243 9373
rect 14185 9333 14197 9367
rect 14231 9364 14243 9367
rect 14274 9364 14280 9376
rect 14231 9336 14280 9364
rect 14231 9333 14243 9336
rect 14185 9327 14243 9333
rect 14274 9324 14280 9336
rect 14332 9324 14338 9376
rect 17034 9324 17040 9376
rect 17092 9324 17098 9376
rect 17678 9324 17684 9376
rect 17736 9364 17742 9376
rect 17773 9367 17831 9373
rect 17773 9364 17785 9367
rect 17736 9336 17785 9364
rect 17736 9324 17742 9336
rect 17773 9333 17785 9336
rect 17819 9333 17831 9367
rect 17773 9327 17831 9333
rect 18138 9324 18144 9376
rect 18196 9364 18202 9376
rect 18616 9364 18644 9404
rect 18196 9336 18644 9364
rect 19168 9364 19196 9404
rect 22557 9401 22569 9404
rect 22603 9401 22615 9435
rect 22756 9432 22784 9463
rect 22922 9460 22928 9512
rect 22980 9460 22986 9512
rect 22830 9432 22836 9444
rect 22756 9404 22836 9432
rect 22557 9395 22615 9401
rect 22830 9392 22836 9404
rect 22888 9392 22894 9444
rect 19242 9364 19248 9376
rect 19168 9336 19248 9364
rect 18196 9324 18202 9336
rect 19242 9324 19248 9336
rect 19300 9324 19306 9376
rect 19337 9367 19395 9373
rect 19337 9333 19349 9367
rect 19383 9364 19395 9367
rect 20070 9364 20076 9376
rect 19383 9336 20076 9364
rect 19383 9333 19395 9336
rect 19337 9327 19395 9333
rect 20070 9324 20076 9336
rect 20128 9324 20134 9376
rect 20438 9324 20444 9376
rect 20496 9324 20502 9376
rect 21266 9324 21272 9376
rect 21324 9364 21330 9376
rect 21361 9367 21419 9373
rect 21361 9364 21373 9367
rect 21324 9336 21373 9364
rect 21324 9324 21330 9336
rect 21361 9333 21373 9336
rect 21407 9333 21419 9367
rect 21361 9327 21419 9333
rect 21818 9324 21824 9376
rect 21876 9364 21882 9376
rect 21913 9367 21971 9373
rect 21913 9364 21925 9367
rect 21876 9336 21925 9364
rect 21876 9324 21882 9336
rect 21913 9333 21925 9336
rect 21959 9333 21971 9367
rect 21913 9327 21971 9333
rect 552 9274 23368 9296
rect 552 9222 4366 9274
rect 4418 9222 4430 9274
rect 4482 9222 4494 9274
rect 4546 9222 4558 9274
rect 4610 9222 4622 9274
rect 4674 9222 4686 9274
rect 4738 9222 10366 9274
rect 10418 9222 10430 9274
rect 10482 9222 10494 9274
rect 10546 9222 10558 9274
rect 10610 9222 10622 9274
rect 10674 9222 10686 9274
rect 10738 9222 16366 9274
rect 16418 9222 16430 9274
rect 16482 9222 16494 9274
rect 16546 9222 16558 9274
rect 16610 9222 16622 9274
rect 16674 9222 16686 9274
rect 16738 9222 22366 9274
rect 22418 9222 22430 9274
rect 22482 9222 22494 9274
rect 22546 9222 22558 9274
rect 22610 9222 22622 9274
rect 22674 9222 22686 9274
rect 22738 9222 23368 9274
rect 552 9200 23368 9222
rect 1118 9120 1124 9172
rect 1176 9120 1182 9172
rect 1578 9160 1584 9172
rect 1228 9132 1584 9160
rect 1118 8984 1124 9036
rect 1176 9024 1182 9036
rect 1228 9024 1256 9132
rect 1578 9120 1584 9132
rect 1636 9120 1642 9172
rect 2590 9160 2596 9172
rect 2148 9132 2596 9160
rect 1854 9092 1860 9104
rect 1320 9064 1860 9092
rect 1320 9033 1348 9064
rect 1854 9052 1860 9064
rect 1912 9052 1918 9104
rect 2148 9101 2176 9132
rect 2590 9120 2596 9132
rect 2648 9120 2654 9172
rect 3326 9120 3332 9172
rect 3384 9160 3390 9172
rect 3786 9160 3792 9172
rect 3384 9132 3792 9160
rect 3384 9120 3390 9132
rect 3786 9120 3792 9132
rect 3844 9120 3850 9172
rect 4246 9120 4252 9172
rect 4304 9160 4310 9172
rect 4341 9163 4399 9169
rect 4341 9160 4353 9163
rect 4304 9132 4353 9160
rect 4304 9120 4310 9132
rect 4341 9129 4353 9132
rect 4387 9129 4399 9163
rect 4341 9123 4399 9129
rect 6270 9120 6276 9172
rect 6328 9120 6334 9172
rect 7834 9120 7840 9172
rect 7892 9160 7898 9172
rect 8110 9160 8116 9172
rect 7892 9132 8116 9160
rect 7892 9120 7898 9132
rect 8110 9120 8116 9132
rect 8168 9120 8174 9172
rect 8294 9120 8300 9172
rect 8352 9160 8358 9172
rect 8352 9132 11284 9160
rect 8352 9120 8358 9132
rect 2133 9095 2191 9101
rect 2133 9061 2145 9095
rect 2179 9061 2191 9095
rect 2133 9055 2191 9061
rect 2685 9095 2743 9101
rect 2685 9061 2697 9095
rect 2731 9092 2743 9095
rect 2866 9092 2872 9104
rect 2731 9064 2872 9092
rect 2731 9061 2743 9064
rect 2685 9055 2743 9061
rect 2866 9052 2872 9064
rect 2924 9052 2930 9104
rect 4154 9052 4160 9104
rect 4212 9092 4218 9104
rect 4982 9092 4988 9104
rect 4212 9064 4988 9092
rect 4212 9052 4218 9064
rect 4982 9052 4988 9064
rect 5040 9052 5046 9104
rect 6178 9052 6184 9104
rect 6236 9092 6242 9104
rect 8757 9095 8815 9101
rect 8757 9092 8769 9095
rect 6236 9064 8769 9092
rect 6236 9052 6242 9064
rect 8757 9061 8769 9064
rect 8803 9061 8815 9095
rect 8757 9055 8815 9061
rect 8941 9095 8999 9101
rect 8941 9061 8953 9095
rect 8987 9092 8999 9095
rect 11146 9092 11152 9104
rect 8987 9064 11152 9092
rect 8987 9061 8999 9064
rect 8941 9055 8999 9061
rect 1176 8996 1256 9024
rect 1305 9027 1363 9033
rect 1176 8984 1182 8996
rect 1305 8993 1317 9027
rect 1351 8993 1363 9027
rect 1305 8987 1363 8993
rect 1762 8984 1768 9036
rect 1820 8984 1826 9036
rect 1949 9027 2007 9033
rect 1949 8993 1961 9027
rect 1995 8993 2007 9027
rect 1949 8987 2007 8993
rect 2317 9027 2375 9033
rect 2317 8993 2329 9027
rect 2363 9024 2375 9027
rect 2593 9027 2651 9033
rect 2593 9024 2605 9027
rect 2363 8996 2605 9024
rect 2363 8993 2375 8996
rect 2317 8987 2375 8993
rect 2593 8993 2605 8996
rect 2639 8993 2651 9027
rect 2593 8987 2651 8993
rect 1026 8916 1032 8968
rect 1084 8956 1090 8968
rect 1670 8956 1676 8968
rect 1084 8928 1676 8956
rect 1084 8916 1090 8928
rect 1670 8916 1676 8928
rect 1728 8956 1734 8968
rect 1964 8956 1992 8987
rect 2774 8984 2780 9036
rect 2832 8984 2838 9036
rect 2958 8984 2964 9036
rect 3016 8984 3022 9036
rect 3050 8984 3056 9036
rect 3108 8984 3114 9036
rect 3329 9027 3387 9033
rect 3329 8993 3341 9027
rect 3375 9024 3387 9027
rect 3510 9024 3516 9036
rect 3375 8996 3516 9024
rect 3375 8993 3387 8996
rect 3329 8987 3387 8993
rect 3510 8984 3516 8996
rect 3568 8984 3574 9036
rect 3973 9027 4031 9033
rect 3973 8993 3985 9027
rect 4019 9024 4031 9027
rect 4062 9024 4068 9036
rect 4019 8996 4068 9024
rect 4019 8993 4031 8996
rect 3973 8987 4031 8993
rect 4062 8984 4068 8996
rect 4120 8984 4126 9036
rect 4433 9027 4491 9033
rect 4433 8993 4445 9027
rect 4479 9024 4491 9027
rect 4798 9024 4804 9036
rect 4479 8996 4804 9024
rect 4479 8993 4491 8996
rect 4433 8987 4491 8993
rect 4798 8984 4804 8996
rect 4856 8984 4862 9036
rect 5626 8984 5632 9036
rect 5684 9024 5690 9036
rect 5813 9027 5871 9033
rect 5813 9024 5825 9027
rect 5684 8996 5825 9024
rect 5684 8984 5690 8996
rect 5813 8993 5825 8996
rect 5859 8993 5871 9027
rect 5813 8987 5871 8993
rect 5902 8984 5908 9036
rect 5960 9024 5966 9036
rect 6914 9024 6920 9036
rect 5960 8996 6920 9024
rect 5960 8984 5966 8996
rect 6914 8984 6920 8996
rect 6972 8984 6978 9036
rect 7098 8984 7104 9036
rect 7156 9024 7162 9036
rect 7193 9027 7251 9033
rect 7193 9024 7205 9027
rect 7156 8996 7205 9024
rect 7156 8984 7162 8996
rect 7193 8993 7205 8996
rect 7239 8993 7251 9027
rect 7193 8987 7251 8993
rect 7282 8984 7288 9036
rect 7340 9024 7346 9036
rect 7465 9027 7523 9033
rect 7340 9022 7420 9024
rect 7465 9022 7477 9027
rect 7340 8996 7477 9022
rect 7340 8984 7346 8996
rect 7392 8994 7477 8996
rect 7465 8993 7477 8994
rect 7511 9022 7523 9027
rect 8294 9024 8300 9036
rect 7576 9022 8300 9024
rect 7511 8996 8300 9022
rect 7511 8994 7604 8996
rect 7511 8993 7523 8994
rect 7465 8987 7523 8993
rect 8294 8984 8300 8996
rect 8352 8984 8358 9036
rect 8772 9024 8800 9055
rect 11146 9052 11152 9064
rect 11204 9052 11210 9104
rect 11256 9092 11284 9132
rect 11330 9120 11336 9172
rect 11388 9120 11394 9172
rect 11422 9120 11428 9172
rect 11480 9160 11486 9172
rect 11480 9132 12480 9160
rect 11480 9120 11486 9132
rect 12452 9092 12480 9132
rect 12526 9120 12532 9172
rect 12584 9160 12590 9172
rect 17770 9160 17776 9172
rect 12584 9132 17776 9160
rect 12584 9120 12590 9132
rect 13814 9092 13820 9104
rect 11256 9064 11468 9092
rect 12452 9064 13820 9092
rect 9766 9024 9772 9036
rect 8772 8996 9772 9024
rect 9766 8984 9772 8996
rect 9824 8984 9830 9036
rect 10965 9027 11023 9033
rect 10965 9024 10977 9027
rect 10336 8996 10977 9024
rect 3237 8959 3295 8965
rect 3237 8956 3249 8959
rect 1728 8928 1992 8956
rect 2746 8928 3249 8956
rect 1728 8916 1734 8928
rect 2409 8891 2467 8897
rect 2409 8857 2421 8891
rect 2455 8888 2467 8891
rect 2746 8888 2774 8928
rect 3237 8925 3249 8928
rect 3283 8925 3295 8959
rect 3237 8919 3295 8925
rect 3786 8916 3792 8968
rect 3844 8956 3850 8968
rect 5350 8956 5356 8968
rect 3844 8928 5356 8956
rect 3844 8916 3850 8928
rect 5350 8916 5356 8928
rect 5408 8916 5414 8968
rect 6362 8916 6368 8968
rect 6420 8956 6426 8968
rect 6420 8928 7696 8956
rect 6420 8916 6426 8928
rect 7190 8888 7196 8900
rect 2455 8860 2774 8888
rect 3436 8860 7196 8888
rect 2455 8857 2467 8860
rect 2409 8851 2467 8857
rect 2038 8780 2044 8832
rect 2096 8820 2102 8832
rect 3436 8820 3464 8860
rect 7190 8848 7196 8860
rect 7248 8888 7254 8900
rect 7377 8891 7435 8897
rect 7377 8888 7389 8891
rect 7248 8860 7389 8888
rect 7248 8848 7254 8860
rect 7377 8857 7389 8860
rect 7423 8857 7435 8891
rect 7668 8888 7696 8928
rect 7742 8916 7748 8968
rect 7800 8956 7806 8968
rect 7837 8959 7895 8965
rect 7837 8956 7849 8959
rect 7800 8928 7849 8956
rect 7800 8916 7806 8928
rect 7837 8925 7849 8928
rect 7883 8925 7895 8959
rect 7837 8919 7895 8925
rect 8110 8916 8116 8968
rect 8168 8916 8174 8968
rect 10336 8956 10364 8996
rect 10965 8993 10977 8996
rect 11011 9024 11023 9027
rect 11054 9024 11060 9036
rect 11011 8996 11060 9024
rect 11011 8993 11023 8996
rect 10965 8987 11023 8993
rect 11054 8984 11060 8996
rect 11112 8984 11118 9036
rect 11440 9024 11468 9064
rect 13814 9052 13820 9064
rect 13872 9052 13878 9104
rect 14568 9064 15148 9092
rect 12158 9024 12164 9036
rect 11440 8996 12164 9024
rect 12158 8984 12164 8996
rect 12216 8984 12222 9036
rect 14090 8984 14096 9036
rect 14148 8984 14154 9036
rect 14185 9027 14243 9033
rect 14185 8993 14197 9027
rect 14231 8993 14243 9027
rect 14185 8987 14243 8993
rect 14461 9028 14519 9033
rect 14568 9028 14596 9064
rect 15120 9036 15148 9064
rect 14461 9027 14596 9028
rect 14461 8993 14473 9027
rect 14507 9000 14596 9027
rect 14507 8993 14519 9000
rect 14461 8987 14519 8993
rect 8864 8928 10364 8956
rect 8864 8888 8892 8928
rect 10410 8916 10416 8968
rect 10468 8956 10474 8968
rect 14200 8956 14228 8987
rect 14734 8984 14740 9036
rect 14792 8984 14798 9036
rect 14829 9027 14887 9033
rect 14829 8993 14841 9027
rect 14875 9024 14887 9027
rect 15010 9024 15016 9036
rect 14875 8996 15016 9024
rect 14875 8993 14887 8996
rect 14829 8987 14887 8993
rect 15010 8984 15016 8996
rect 15068 8984 15074 9036
rect 15102 8984 15108 9036
rect 15160 8984 15166 9036
rect 15197 9027 15255 9033
rect 15197 8993 15209 9027
rect 15243 9024 15255 9027
rect 15396 9024 15424 9132
rect 17770 9120 17776 9132
rect 17828 9120 17834 9172
rect 18138 9160 18144 9172
rect 17972 9132 18144 9160
rect 16117 9095 16175 9101
rect 16117 9092 16129 9095
rect 15488 9064 16129 9092
rect 15488 9033 15516 9064
rect 16117 9061 16129 9064
rect 16163 9061 16175 9095
rect 16117 9055 16175 9061
rect 16301 9095 16359 9101
rect 16301 9061 16313 9095
rect 16347 9092 16359 9095
rect 17126 9092 17132 9104
rect 16347 9064 17132 9092
rect 16347 9061 16359 9064
rect 16301 9055 16359 9061
rect 17126 9052 17132 9064
rect 17184 9052 17190 9104
rect 17586 9052 17592 9104
rect 17644 9092 17650 9104
rect 17972 9101 18000 9132
rect 18138 9120 18144 9132
rect 18196 9120 18202 9172
rect 19242 9160 19248 9172
rect 18800 9132 19248 9160
rect 17957 9095 18015 9101
rect 17957 9092 17969 9095
rect 17644 9064 17969 9092
rect 17644 9052 17650 9064
rect 17957 9061 17969 9064
rect 18003 9061 18015 9095
rect 18800 9092 18828 9132
rect 19242 9120 19248 9132
rect 19300 9160 19306 9172
rect 21910 9160 21916 9172
rect 19300 9132 21916 9160
rect 19300 9120 19306 9132
rect 21910 9120 21916 9132
rect 21968 9160 21974 9172
rect 22005 9163 22063 9169
rect 22005 9160 22017 9163
rect 21968 9132 22017 9160
rect 21968 9120 21974 9132
rect 22005 9129 22017 9132
rect 22051 9129 22063 9163
rect 22005 9123 22063 9129
rect 22646 9120 22652 9172
rect 22704 9160 22710 9172
rect 22922 9160 22928 9172
rect 22704 9132 22928 9160
rect 22704 9120 22710 9132
rect 22922 9120 22928 9132
rect 22980 9120 22986 9172
rect 19153 9095 19211 9101
rect 18800 9064 18920 9092
rect 17957 9055 18015 9061
rect 15243 8996 15424 9024
rect 15473 9027 15531 9033
rect 15243 8993 15255 8996
rect 15197 8987 15255 8993
rect 15473 8993 15485 9027
rect 15519 8993 15531 9027
rect 15473 8987 15531 8993
rect 15657 9027 15715 9033
rect 15657 8993 15669 9027
rect 15703 9024 15715 9027
rect 15838 9024 15844 9036
rect 15703 8996 15844 9024
rect 15703 8993 15715 8996
rect 15657 8987 15715 8993
rect 15488 8956 15516 8987
rect 15838 8984 15844 8996
rect 15896 9024 15902 9036
rect 17773 9027 17831 9033
rect 17773 9024 17785 9027
rect 15896 8996 17785 9024
rect 15896 8984 15902 8996
rect 17773 8993 17785 8996
rect 17819 8993 17831 9027
rect 17773 8987 17831 8993
rect 10468 8928 15516 8956
rect 10468 8916 10474 8928
rect 7668 8860 8892 8888
rect 7377 8851 7435 8857
rect 8938 8848 8944 8900
rect 8996 8888 9002 8900
rect 10870 8888 10876 8900
rect 8996 8860 10876 8888
rect 8996 8848 9002 8860
rect 10870 8848 10876 8860
rect 10928 8848 10934 8900
rect 11330 8848 11336 8900
rect 11388 8888 11394 8900
rect 15396 8897 15424 8928
rect 15746 8916 15752 8968
rect 15804 8956 15810 8968
rect 16298 8956 16304 8968
rect 15804 8928 16304 8956
rect 15804 8916 15810 8928
rect 16298 8916 16304 8928
rect 16356 8916 16362 8968
rect 16574 8916 16580 8968
rect 16632 8956 16638 8968
rect 17218 8956 17224 8968
rect 16632 8928 17224 8956
rect 16632 8916 16638 8928
rect 17218 8916 17224 8928
rect 17276 8916 17282 8968
rect 17788 8956 17816 8987
rect 18230 8984 18236 9036
rect 18288 9033 18294 9036
rect 18288 9027 18311 9033
rect 18299 8993 18311 9027
rect 18288 8987 18311 8993
rect 18417 9027 18475 9033
rect 18417 8993 18429 9027
rect 18463 8993 18475 9027
rect 18417 8987 18475 8993
rect 18288 8984 18294 8987
rect 18432 8956 18460 8987
rect 18506 8984 18512 9036
rect 18564 8984 18570 9036
rect 18892 9033 18920 9064
rect 19153 9061 19165 9095
rect 19199 9092 19211 9095
rect 21726 9092 21732 9104
rect 19199 9064 21732 9092
rect 19199 9061 19211 9064
rect 19153 9055 19211 9061
rect 21726 9052 21732 9064
rect 21784 9052 21790 9104
rect 22278 9052 22284 9104
rect 22336 9092 22342 9104
rect 22465 9095 22523 9101
rect 22465 9092 22477 9095
rect 22336 9064 22477 9092
rect 22336 9052 22342 9064
rect 22465 9061 22477 9064
rect 22511 9092 22523 9095
rect 22511 9064 22968 9092
rect 22511 9061 22523 9064
rect 22465 9055 22523 9061
rect 18601 9027 18659 9033
rect 18601 8993 18613 9027
rect 18647 8993 18659 9027
rect 18892 9027 18955 9033
rect 18892 8996 18909 9027
rect 18601 8987 18659 8993
rect 18897 8993 18909 8996
rect 18943 8993 18955 9027
rect 18897 8987 18955 8993
rect 17788 8928 18460 8956
rect 18616 8956 18644 8987
rect 19058 8984 19064 9036
rect 19116 8984 19122 9036
rect 19245 9027 19303 9033
rect 19245 9024 19257 9027
rect 19168 8996 19257 9024
rect 19168 8956 19196 8996
rect 19245 8993 19257 8996
rect 19291 8993 19303 9027
rect 19245 8987 19303 8993
rect 19702 8984 19708 9036
rect 19760 9024 19766 9036
rect 19797 9027 19855 9033
rect 19797 9024 19809 9027
rect 19760 8996 19809 9024
rect 19760 8984 19766 8996
rect 19797 8993 19809 8996
rect 19843 8993 19855 9027
rect 19797 8987 19855 8993
rect 19886 8984 19892 9036
rect 19944 9024 19950 9036
rect 20073 9027 20131 9033
rect 20073 9024 20085 9027
rect 19944 8996 20085 9024
rect 19944 8984 19950 8996
rect 20073 8993 20085 8996
rect 20119 8993 20131 9027
rect 20073 8987 20131 8993
rect 21450 8984 21456 9036
rect 21508 9024 21514 9036
rect 22094 9024 22100 9036
rect 21508 8996 22100 9024
rect 21508 8984 21514 8996
rect 22094 8984 22100 8996
rect 22152 8984 22158 9036
rect 22189 9027 22247 9033
rect 22189 8993 22201 9027
rect 22235 9024 22247 9027
rect 22296 9024 22324 9052
rect 22235 8996 22324 9024
rect 22235 8993 22247 8996
rect 22189 8987 22247 8993
rect 22646 8984 22652 9036
rect 22704 9024 22710 9036
rect 22940 9033 22968 9064
rect 22741 9027 22799 9033
rect 22741 9024 22753 9027
rect 22704 8996 22753 9024
rect 22704 8984 22710 8996
rect 22741 8993 22753 8996
rect 22787 8993 22799 9027
rect 22741 8987 22799 8993
rect 22925 9027 22983 9033
rect 22925 8993 22937 9027
rect 22971 8993 22983 9027
rect 22925 8987 22983 8993
rect 22833 8959 22891 8965
rect 22833 8956 22845 8959
rect 18616 8928 22845 8956
rect 22833 8925 22845 8928
rect 22879 8925 22891 8959
rect 22833 8919 22891 8925
rect 14369 8891 14427 8897
rect 14369 8888 14381 8891
rect 11388 8860 14381 8888
rect 11388 8848 11394 8860
rect 14369 8857 14381 8860
rect 14415 8888 14427 8891
rect 15381 8891 15439 8897
rect 14415 8860 15240 8888
rect 14415 8857 14427 8860
rect 14369 8851 14427 8857
rect 2096 8792 3464 8820
rect 2096 8780 2102 8792
rect 3510 8780 3516 8832
rect 3568 8820 3574 8832
rect 3605 8823 3663 8829
rect 3605 8820 3617 8823
rect 3568 8792 3617 8820
rect 3568 8780 3574 8792
rect 3605 8789 3617 8792
rect 3651 8789 3663 8823
rect 3605 8783 3663 8789
rect 4154 8780 4160 8832
rect 4212 8780 4218 8832
rect 5534 8780 5540 8832
rect 5592 8820 5598 8832
rect 5905 8823 5963 8829
rect 5905 8820 5917 8823
rect 5592 8792 5917 8820
rect 5592 8780 5598 8792
rect 5905 8789 5917 8792
rect 5951 8789 5963 8823
rect 5905 8783 5963 8789
rect 6914 8780 6920 8832
rect 6972 8820 6978 8832
rect 7009 8823 7067 8829
rect 7009 8820 7021 8823
rect 6972 8792 7021 8820
rect 6972 8780 6978 8792
rect 7009 8789 7021 8792
rect 7055 8789 7067 8823
rect 7009 8783 7067 8789
rect 7098 8780 7104 8832
rect 7156 8820 7162 8832
rect 7742 8820 7748 8832
rect 7156 8792 7748 8820
rect 7156 8780 7162 8792
rect 7742 8780 7748 8792
rect 7800 8780 7806 8832
rect 8570 8780 8576 8832
rect 8628 8820 8634 8832
rect 9125 8823 9183 8829
rect 9125 8820 9137 8823
rect 8628 8792 9137 8820
rect 8628 8780 8634 8792
rect 9125 8789 9137 8792
rect 9171 8789 9183 8823
rect 9125 8783 9183 8789
rect 9674 8780 9680 8832
rect 9732 8820 9738 8832
rect 11698 8820 11704 8832
rect 9732 8792 11704 8820
rect 9732 8780 9738 8792
rect 11698 8780 11704 8792
rect 11756 8780 11762 8832
rect 11974 8780 11980 8832
rect 12032 8820 12038 8832
rect 12250 8820 12256 8832
rect 12032 8792 12256 8820
rect 12032 8780 12038 8792
rect 12250 8780 12256 8792
rect 12308 8780 12314 8832
rect 12342 8780 12348 8832
rect 12400 8820 12406 8832
rect 12894 8820 12900 8832
rect 12400 8792 12900 8820
rect 12400 8780 12406 8792
rect 12894 8780 12900 8792
rect 12952 8780 12958 8832
rect 13814 8780 13820 8832
rect 13872 8820 13878 8832
rect 13909 8823 13967 8829
rect 13909 8820 13921 8823
rect 13872 8792 13921 8820
rect 13872 8780 13878 8792
rect 13909 8789 13921 8792
rect 13955 8789 13967 8823
rect 13909 8783 13967 8789
rect 14550 8780 14556 8832
rect 14608 8780 14614 8832
rect 14642 8780 14648 8832
rect 14700 8820 14706 8832
rect 15013 8823 15071 8829
rect 15013 8820 15025 8823
rect 14700 8792 15025 8820
rect 14700 8780 14706 8792
rect 15013 8789 15025 8792
rect 15059 8820 15071 8823
rect 15102 8820 15108 8832
rect 15059 8792 15108 8820
rect 15059 8789 15071 8792
rect 15013 8783 15071 8789
rect 15102 8780 15108 8792
rect 15160 8780 15166 8832
rect 15212 8820 15240 8860
rect 15381 8857 15393 8891
rect 15427 8857 15439 8891
rect 16666 8888 16672 8900
rect 15381 8851 15439 8857
rect 15488 8860 16672 8888
rect 15488 8820 15516 8860
rect 16666 8848 16672 8860
rect 16724 8848 16730 8900
rect 17236 8888 17264 8916
rect 18506 8888 18512 8900
rect 17236 8860 18512 8888
rect 18506 8848 18512 8860
rect 18564 8848 18570 8900
rect 19886 8848 19892 8900
rect 19944 8848 19950 8900
rect 19981 8891 20039 8897
rect 19981 8857 19993 8891
rect 20027 8888 20039 8891
rect 20346 8888 20352 8900
rect 20027 8860 20352 8888
rect 20027 8857 20039 8860
rect 19981 8851 20039 8857
rect 20346 8848 20352 8860
rect 20404 8848 20410 8900
rect 20714 8848 20720 8900
rect 20772 8888 20778 8900
rect 22281 8891 22339 8897
rect 22281 8888 22293 8891
rect 20772 8860 22293 8888
rect 20772 8848 20778 8860
rect 22281 8857 22293 8860
rect 22327 8857 22339 8891
rect 22281 8851 22339 8857
rect 15212 8792 15516 8820
rect 15841 8823 15899 8829
rect 15841 8789 15853 8823
rect 15887 8820 15899 8823
rect 16022 8820 16028 8832
rect 15887 8792 16028 8820
rect 15887 8789 15899 8792
rect 15841 8783 15899 8789
rect 16022 8780 16028 8792
rect 16080 8780 16086 8832
rect 16485 8823 16543 8829
rect 16485 8789 16497 8823
rect 16531 8820 16543 8823
rect 16850 8820 16856 8832
rect 16531 8792 16856 8820
rect 16531 8789 16543 8792
rect 16485 8783 16543 8789
rect 16850 8780 16856 8792
rect 16908 8780 16914 8832
rect 18141 8823 18199 8829
rect 18141 8789 18153 8823
rect 18187 8820 18199 8823
rect 18414 8820 18420 8832
rect 18187 8792 18420 8820
rect 18187 8789 18199 8792
rect 18141 8783 18199 8789
rect 18414 8780 18420 8792
rect 18472 8780 18478 8832
rect 18785 8823 18843 8829
rect 18785 8789 18797 8823
rect 18831 8820 18843 8823
rect 18874 8820 18880 8832
rect 18831 8792 18880 8820
rect 18831 8789 18843 8792
rect 18785 8783 18843 8789
rect 18874 8780 18880 8792
rect 18932 8780 18938 8832
rect 19429 8823 19487 8829
rect 19429 8789 19441 8823
rect 19475 8820 19487 8823
rect 19794 8820 19800 8832
rect 19475 8792 19800 8820
rect 19475 8789 19487 8792
rect 19429 8783 19487 8789
rect 19794 8780 19800 8792
rect 19852 8780 19858 8832
rect 20257 8823 20315 8829
rect 20257 8789 20269 8823
rect 20303 8820 20315 8823
rect 20622 8820 20628 8832
rect 20303 8792 20628 8820
rect 20303 8789 20315 8792
rect 20257 8783 20315 8789
rect 20622 8780 20628 8792
rect 20680 8780 20686 8832
rect 21082 8780 21088 8832
rect 21140 8820 21146 8832
rect 21269 8823 21327 8829
rect 21269 8820 21281 8823
rect 21140 8792 21281 8820
rect 21140 8780 21146 8792
rect 21269 8789 21281 8792
rect 21315 8789 21327 8823
rect 21269 8783 21327 8789
rect 552 8730 23368 8752
rect 552 8678 1366 8730
rect 1418 8678 1430 8730
rect 1482 8678 1494 8730
rect 1546 8678 1558 8730
rect 1610 8678 1622 8730
rect 1674 8678 1686 8730
rect 1738 8678 7366 8730
rect 7418 8678 7430 8730
rect 7482 8678 7494 8730
rect 7546 8678 7558 8730
rect 7610 8678 7622 8730
rect 7674 8678 7686 8730
rect 7738 8678 13366 8730
rect 13418 8678 13430 8730
rect 13482 8678 13494 8730
rect 13546 8678 13558 8730
rect 13610 8678 13622 8730
rect 13674 8678 13686 8730
rect 13738 8678 19366 8730
rect 19418 8678 19430 8730
rect 19482 8678 19494 8730
rect 19546 8678 19558 8730
rect 19610 8678 19622 8730
rect 19674 8678 19686 8730
rect 19738 8678 23368 8730
rect 552 8656 23368 8678
rect 1946 8616 1952 8628
rect 1596 8588 1952 8616
rect 1596 8489 1624 8588
rect 1946 8576 1952 8588
rect 2004 8616 2010 8628
rect 2498 8616 2504 8628
rect 2004 8588 2504 8616
rect 2004 8576 2010 8588
rect 2498 8576 2504 8588
rect 2556 8576 2562 8628
rect 3510 8576 3516 8628
rect 3568 8576 3574 8628
rect 4798 8576 4804 8628
rect 4856 8616 4862 8628
rect 5261 8619 5319 8625
rect 5261 8616 5273 8619
rect 4856 8588 5273 8616
rect 4856 8576 4862 8588
rect 5261 8585 5273 8588
rect 5307 8585 5319 8619
rect 5261 8579 5319 8585
rect 1857 8551 1915 8557
rect 1857 8517 1869 8551
rect 1903 8548 1915 8551
rect 2593 8551 2651 8557
rect 1903 8520 2176 8548
rect 1903 8517 1915 8520
rect 1857 8511 1915 8517
rect 2148 8489 2176 8520
rect 2593 8517 2605 8551
rect 2639 8548 2651 8551
rect 4065 8551 4123 8557
rect 4065 8548 4077 8551
rect 2639 8520 2774 8548
rect 2639 8517 2651 8520
rect 2593 8511 2651 8517
rect 1581 8483 1639 8489
rect 1581 8449 1593 8483
rect 1627 8449 1639 8483
rect 1581 8443 1639 8449
rect 2133 8483 2191 8489
rect 2133 8449 2145 8483
rect 2179 8449 2191 8483
rect 2133 8443 2191 8449
rect 1489 8415 1547 8421
rect 1489 8381 1501 8415
rect 1535 8412 1547 8415
rect 2038 8412 2044 8424
rect 1535 8384 2044 8412
rect 1535 8381 1547 8384
rect 1489 8375 1547 8381
rect 2038 8372 2044 8384
rect 2096 8372 2102 8424
rect 2222 8372 2228 8424
rect 2280 8372 2286 8424
rect 2746 8344 2774 8520
rect 3715 8520 4077 8548
rect 3715 8489 3743 8520
rect 4065 8517 4077 8520
rect 4111 8517 4123 8551
rect 5166 8548 5172 8560
rect 4065 8511 4123 8517
rect 4724 8520 5172 8548
rect 3697 8483 3755 8489
rect 3697 8449 3709 8483
rect 3743 8449 3755 8483
rect 3697 8443 3755 8449
rect 4525 8483 4583 8489
rect 4525 8449 4537 8483
rect 4571 8480 4583 8483
rect 4724 8480 4752 8520
rect 5166 8508 5172 8520
rect 5224 8508 5230 8560
rect 5276 8548 5304 8579
rect 5718 8576 5724 8628
rect 5776 8576 5782 8628
rect 6546 8576 6552 8628
rect 6604 8616 6610 8628
rect 8938 8616 8944 8628
rect 6604 8588 8944 8616
rect 6604 8576 6610 8588
rect 8938 8576 8944 8588
rect 8996 8576 9002 8628
rect 9490 8616 9496 8628
rect 9324 8588 9496 8616
rect 9324 8548 9352 8588
rect 9490 8576 9496 8588
rect 9548 8576 9554 8628
rect 9582 8576 9588 8628
rect 9640 8616 9646 8628
rect 9640 8588 10548 8616
rect 9640 8576 9646 8588
rect 5276 8520 9352 8548
rect 9398 8508 9404 8560
rect 9456 8548 9462 8560
rect 9456 8520 9674 8548
rect 9456 8508 9462 8520
rect 4571 8452 4752 8480
rect 4571 8449 4583 8452
rect 4525 8443 4583 8449
rect 4798 8440 4804 8492
rect 4856 8440 4862 8492
rect 5350 8440 5356 8492
rect 5408 8480 5414 8492
rect 6362 8480 6368 8492
rect 5408 8452 5580 8480
rect 5408 8440 5414 8452
rect 3142 8372 3148 8424
rect 3200 8412 3206 8424
rect 3421 8415 3479 8421
rect 3421 8412 3433 8415
rect 3200 8384 3433 8412
rect 3200 8372 3206 8384
rect 3421 8381 3433 8384
rect 3467 8381 3479 8415
rect 3421 8375 3479 8381
rect 3510 8372 3516 8424
rect 3568 8412 3574 8424
rect 3789 8415 3847 8421
rect 3789 8412 3801 8415
rect 3568 8384 3801 8412
rect 3568 8372 3574 8384
rect 3789 8381 3801 8384
rect 3835 8381 3847 8415
rect 3789 8375 3847 8381
rect 4433 8415 4491 8421
rect 4433 8381 4445 8415
rect 4479 8381 4491 8415
rect 4433 8375 4491 8381
rect 2746 8316 4016 8344
rect 3510 8236 3516 8288
rect 3568 8276 3574 8288
rect 3697 8279 3755 8285
rect 3697 8276 3709 8279
rect 3568 8248 3709 8276
rect 3568 8236 3574 8248
rect 3697 8245 3709 8248
rect 3743 8245 3755 8279
rect 3697 8239 3755 8245
rect 3786 8236 3792 8288
rect 3844 8276 3850 8288
rect 3881 8279 3939 8285
rect 3881 8276 3893 8279
rect 3844 8248 3893 8276
rect 3844 8236 3850 8248
rect 3881 8245 3893 8248
rect 3927 8245 3939 8279
rect 3988 8276 4016 8316
rect 4062 8304 4068 8356
rect 4120 8304 4126 8356
rect 4448 8344 4476 8375
rect 4890 8372 4896 8424
rect 4948 8412 4954 8424
rect 5552 8421 5580 8452
rect 6196 8452 6368 8480
rect 5169 8415 5227 8421
rect 5169 8412 5181 8415
rect 4948 8384 5181 8412
rect 4948 8372 4954 8384
rect 5169 8381 5181 8384
rect 5215 8381 5227 8415
rect 5169 8375 5227 8381
rect 5445 8415 5503 8421
rect 5445 8381 5457 8415
rect 5491 8381 5503 8415
rect 5445 8375 5503 8381
rect 5537 8415 5595 8421
rect 5537 8381 5549 8415
rect 5583 8381 5595 8415
rect 5537 8375 5595 8381
rect 5997 8415 6055 8421
rect 5997 8381 6009 8415
rect 6043 8412 6055 8415
rect 6086 8412 6092 8424
rect 6043 8384 6092 8412
rect 6043 8381 6055 8384
rect 5997 8375 6055 8381
rect 5460 8344 5488 8375
rect 6086 8372 6092 8384
rect 6144 8372 6150 8424
rect 6196 8421 6224 8452
rect 6362 8440 6368 8452
rect 6420 8480 6426 8492
rect 6549 8483 6607 8489
rect 6549 8480 6561 8483
rect 6420 8452 6561 8480
rect 6420 8440 6426 8452
rect 6549 8449 6561 8452
rect 6595 8480 6607 8483
rect 6730 8480 6736 8492
rect 6595 8452 6736 8480
rect 6595 8449 6607 8452
rect 6549 8443 6607 8449
rect 6730 8440 6736 8452
rect 6788 8440 6794 8492
rect 7098 8440 7104 8492
rect 7156 8480 7162 8492
rect 8386 8480 8392 8492
rect 7156 8452 8392 8480
rect 7156 8440 7162 8452
rect 8386 8440 8392 8452
rect 8444 8440 8450 8492
rect 8665 8483 8723 8489
rect 8665 8449 8677 8483
rect 8711 8480 8723 8483
rect 8938 8480 8944 8492
rect 8711 8452 8944 8480
rect 8711 8449 8723 8452
rect 8665 8443 8723 8449
rect 8938 8440 8944 8452
rect 8996 8440 9002 8492
rect 9646 8480 9674 8520
rect 9858 8508 9864 8560
rect 9916 8548 9922 8560
rect 10042 8548 10048 8560
rect 9916 8520 10048 8548
rect 9916 8508 9922 8520
rect 10042 8508 10048 8520
rect 10100 8508 10106 8560
rect 9646 8452 9904 8480
rect 6181 8415 6239 8421
rect 6181 8381 6193 8415
rect 6227 8381 6239 8415
rect 6181 8375 6239 8381
rect 6270 8372 6276 8424
rect 6328 8372 6334 8424
rect 7742 8372 7748 8424
rect 7800 8412 7806 8424
rect 7929 8415 7987 8421
rect 7929 8412 7941 8415
rect 7800 8384 7941 8412
rect 7800 8372 7806 8384
rect 7929 8381 7941 8384
rect 7975 8381 7987 8415
rect 7929 8375 7987 8381
rect 8205 8415 8263 8421
rect 8205 8381 8217 8415
rect 8251 8412 8263 8415
rect 8294 8412 8300 8424
rect 8251 8384 8300 8412
rect 8251 8381 8263 8384
rect 8205 8375 8263 8381
rect 8294 8372 8300 8384
rect 8352 8372 8358 8424
rect 8570 8372 8576 8424
rect 8628 8412 8634 8424
rect 9309 8415 9367 8421
rect 9309 8412 9321 8415
rect 8628 8384 9321 8412
rect 8628 8372 8634 8384
rect 9309 8381 9321 8384
rect 9355 8381 9367 8415
rect 9493 8415 9551 8421
rect 9493 8412 9505 8415
rect 9309 8375 9367 8381
rect 9416 8384 9505 8412
rect 9214 8344 9220 8356
rect 4448 8316 9220 8344
rect 4890 8276 4896 8288
rect 3988 8248 4896 8276
rect 3881 8239 3939 8245
rect 4890 8236 4896 8248
rect 4948 8236 4954 8288
rect 5000 8285 5028 8316
rect 9214 8304 9220 8316
rect 9272 8304 9278 8356
rect 4985 8279 5043 8285
rect 4985 8245 4997 8279
rect 5031 8245 5043 8279
rect 4985 8239 5043 8245
rect 6086 8236 6092 8288
rect 6144 8236 6150 8288
rect 8938 8236 8944 8288
rect 8996 8276 9002 8288
rect 9416 8276 9444 8384
rect 9493 8381 9505 8384
rect 9539 8381 9551 8415
rect 9493 8375 9551 8381
rect 9582 8372 9588 8424
rect 9640 8372 9646 8424
rect 9674 8372 9680 8424
rect 9732 8372 9738 8424
rect 9876 8421 9904 8452
rect 9861 8415 9919 8421
rect 9861 8381 9873 8415
rect 9907 8381 9919 8415
rect 9861 8375 9919 8381
rect 10318 8372 10324 8424
rect 10376 8372 10382 8424
rect 10410 8372 10416 8424
rect 10468 8372 10474 8424
rect 10137 8347 10195 8353
rect 10137 8344 10149 8347
rect 9508 8316 10149 8344
rect 9508 8288 9536 8316
rect 10137 8313 10149 8316
rect 10183 8313 10195 8347
rect 10520 8344 10548 8588
rect 11146 8576 11152 8628
rect 11204 8616 11210 8628
rect 12158 8616 12164 8628
rect 11204 8588 12164 8616
rect 11204 8576 11210 8588
rect 12158 8576 12164 8588
rect 12216 8616 12222 8628
rect 12216 8588 18276 8616
rect 12216 8576 12222 8588
rect 11054 8508 11060 8560
rect 11112 8548 11118 8560
rect 11977 8551 12035 8557
rect 11977 8548 11989 8551
rect 11112 8520 11989 8548
rect 11112 8508 11118 8520
rect 11977 8517 11989 8520
rect 12023 8548 12035 8551
rect 12342 8548 12348 8560
rect 12023 8520 12348 8548
rect 12023 8517 12035 8520
rect 11977 8511 12035 8517
rect 12342 8508 12348 8520
rect 12400 8508 12406 8560
rect 12618 8508 12624 8560
rect 12676 8548 12682 8560
rect 13633 8551 13691 8557
rect 12676 8520 12756 8548
rect 12676 8508 12682 8520
rect 10597 8483 10655 8489
rect 10597 8449 10609 8483
rect 10643 8480 10655 8483
rect 11330 8480 11336 8492
rect 10643 8452 11336 8480
rect 10643 8449 10655 8452
rect 10597 8443 10655 8449
rect 11330 8440 11336 8452
rect 11388 8440 11394 8492
rect 10689 8415 10747 8421
rect 10689 8381 10701 8415
rect 10735 8412 10747 8415
rect 10870 8412 10876 8424
rect 10735 8384 10876 8412
rect 10735 8381 10747 8384
rect 10689 8375 10747 8381
rect 10870 8372 10876 8384
rect 10928 8372 10934 8424
rect 11698 8372 11704 8424
rect 11756 8372 11762 8424
rect 11790 8372 11796 8424
rect 11848 8372 11854 8424
rect 11882 8372 11888 8424
rect 11940 8412 11946 8424
rect 12069 8415 12127 8421
rect 12069 8412 12081 8415
rect 11940 8384 12081 8412
rect 11940 8372 11946 8384
rect 12069 8381 12081 8384
rect 12115 8381 12127 8415
rect 12069 8375 12127 8381
rect 12434 8372 12440 8424
rect 12492 8372 12498 8424
rect 12728 8421 12756 8520
rect 13633 8517 13645 8551
rect 13679 8548 13691 8551
rect 13909 8551 13967 8557
rect 13909 8548 13921 8551
rect 13679 8520 13921 8548
rect 13679 8517 13691 8520
rect 13633 8511 13691 8517
rect 13909 8517 13921 8520
rect 13955 8517 13967 8551
rect 13909 8511 13967 8517
rect 13648 8480 13676 8511
rect 15470 8508 15476 8560
rect 15528 8548 15534 8560
rect 15746 8548 15752 8560
rect 15528 8520 15752 8548
rect 15528 8508 15534 8520
rect 15746 8508 15752 8520
rect 15804 8508 15810 8560
rect 16758 8508 16764 8560
rect 16816 8548 16822 8560
rect 17126 8548 17132 8560
rect 16816 8520 17132 8548
rect 16816 8508 16822 8520
rect 17126 8508 17132 8520
rect 17184 8508 17190 8560
rect 17862 8548 17868 8560
rect 17512 8520 17868 8548
rect 12912 8452 13676 8480
rect 12621 8415 12679 8421
rect 12621 8381 12633 8415
rect 12667 8381 12679 8415
rect 12621 8375 12679 8381
rect 12713 8415 12771 8421
rect 12713 8381 12725 8415
rect 12759 8381 12771 8415
rect 12713 8375 12771 8381
rect 12636 8344 12664 8375
rect 12802 8372 12808 8424
rect 12860 8372 12866 8424
rect 12912 8344 12940 8452
rect 13814 8440 13820 8492
rect 13872 8440 13878 8492
rect 15838 8440 15844 8492
rect 15896 8480 15902 8492
rect 16393 8483 16451 8489
rect 16393 8480 16405 8483
rect 15896 8452 16405 8480
rect 15896 8440 15902 8452
rect 16393 8449 16405 8452
rect 16439 8480 16451 8483
rect 17221 8483 17279 8489
rect 17221 8480 17233 8483
rect 16439 8452 17233 8480
rect 16439 8449 16451 8452
rect 16393 8443 16451 8449
rect 17221 8449 17233 8452
rect 17267 8449 17279 8483
rect 17221 8443 17279 8449
rect 12986 8372 12992 8424
rect 13044 8372 13050 8424
rect 13078 8372 13084 8424
rect 13136 8412 13142 8424
rect 13538 8412 13544 8424
rect 13136 8384 13544 8412
rect 13136 8372 13142 8384
rect 13538 8372 13544 8384
rect 13596 8372 13602 8424
rect 14090 8372 14096 8424
rect 14148 8412 14154 8424
rect 15102 8412 15108 8424
rect 14148 8384 15108 8412
rect 14148 8372 14154 8384
rect 15102 8372 15108 8384
rect 15160 8372 15166 8424
rect 16022 8372 16028 8424
rect 16080 8372 16086 8424
rect 16209 8415 16267 8421
rect 16209 8381 16221 8415
rect 16255 8381 16267 8415
rect 16209 8375 16267 8381
rect 15010 8344 15016 8356
rect 10520 8316 12940 8344
rect 13004 8316 15016 8344
rect 10137 8307 10195 8313
rect 8996 8248 9444 8276
rect 8996 8236 9002 8248
rect 9490 8236 9496 8288
rect 9548 8236 9554 8288
rect 9858 8236 9864 8288
rect 9916 8276 9922 8288
rect 10045 8279 10103 8285
rect 10045 8276 10057 8279
rect 9916 8248 10057 8276
rect 9916 8236 9922 8248
rect 10045 8245 10057 8248
rect 10091 8245 10103 8279
rect 10045 8239 10103 8245
rect 11514 8236 11520 8288
rect 11572 8236 11578 8288
rect 11790 8236 11796 8288
rect 11848 8276 11854 8288
rect 13004 8276 13032 8316
rect 15010 8304 15016 8316
rect 15068 8304 15074 8356
rect 15286 8304 15292 8356
rect 15344 8344 15350 8356
rect 16224 8344 16252 8375
rect 16298 8372 16304 8424
rect 16356 8372 16362 8424
rect 16574 8372 16580 8424
rect 16632 8372 16638 8424
rect 16850 8372 16856 8424
rect 16908 8372 16914 8424
rect 17037 8415 17095 8421
rect 17037 8381 17049 8415
rect 17083 8381 17095 8415
rect 17037 8375 17095 8381
rect 15344 8316 16252 8344
rect 15344 8304 15350 8316
rect 11848 8248 13032 8276
rect 11848 8236 11854 8248
rect 13078 8236 13084 8288
rect 13136 8276 13142 8288
rect 13173 8279 13231 8285
rect 13173 8276 13185 8279
rect 13136 8248 13185 8276
rect 13136 8236 13142 8248
rect 13173 8245 13185 8248
rect 13219 8245 13231 8279
rect 13173 8239 13231 8245
rect 13817 8279 13875 8285
rect 13817 8245 13829 8279
rect 13863 8276 13875 8279
rect 14458 8276 14464 8288
rect 13863 8248 14464 8276
rect 13863 8245 13875 8248
rect 13817 8239 13875 8245
rect 14458 8236 14464 8248
rect 14516 8236 14522 8288
rect 14550 8236 14556 8288
rect 14608 8276 14614 8288
rect 14826 8276 14832 8288
rect 14608 8248 14832 8276
rect 14608 8236 14614 8248
rect 14826 8236 14832 8248
rect 14884 8236 14890 8288
rect 16224 8276 16252 8316
rect 16758 8304 16764 8356
rect 16816 8304 16822 8356
rect 17052 8276 17080 8375
rect 17126 8372 17132 8424
rect 17184 8372 17190 8424
rect 17405 8415 17463 8421
rect 17405 8381 17417 8415
rect 17451 8412 17463 8415
rect 17512 8412 17540 8520
rect 17862 8508 17868 8520
rect 17920 8548 17926 8560
rect 17920 8520 18000 8548
rect 17920 8508 17926 8520
rect 17586 8440 17592 8492
rect 17644 8480 17650 8492
rect 17644 8452 17908 8480
rect 17644 8440 17650 8452
rect 17880 8421 17908 8452
rect 17972 8421 18000 8520
rect 18138 8508 18144 8560
rect 18196 8508 18202 8560
rect 18248 8480 18276 8588
rect 18966 8576 18972 8628
rect 19024 8616 19030 8628
rect 19797 8619 19855 8625
rect 19797 8616 19809 8619
rect 19024 8588 19809 8616
rect 19024 8576 19030 8588
rect 19797 8585 19809 8588
rect 19843 8585 19855 8619
rect 19797 8579 19855 8585
rect 20346 8576 20352 8628
rect 20404 8616 20410 8628
rect 21082 8616 21088 8628
rect 20404 8588 21088 8616
rect 20404 8576 20410 8588
rect 21082 8576 21088 8588
rect 21140 8576 21146 8628
rect 21174 8576 21180 8628
rect 21232 8576 21238 8628
rect 18414 8508 18420 8560
rect 18472 8548 18478 8560
rect 22002 8548 22008 8560
rect 18472 8520 22008 8548
rect 18472 8508 18478 8520
rect 22002 8508 22008 8520
rect 22060 8548 22066 8560
rect 22060 8520 22140 8548
rect 22060 8508 22066 8520
rect 20346 8480 20352 8492
rect 18248 8452 20352 8480
rect 20346 8440 20352 8452
rect 20404 8440 20410 8492
rect 22112 8480 22140 8520
rect 22465 8483 22523 8489
rect 22465 8480 22477 8483
rect 22112 8452 22477 8480
rect 17451 8384 17540 8412
rect 17865 8415 17923 8421
rect 17451 8381 17463 8384
rect 17405 8375 17463 8381
rect 17865 8381 17877 8415
rect 17911 8381 17923 8415
rect 17865 8375 17923 8381
rect 17957 8415 18015 8421
rect 17957 8381 17969 8415
rect 18003 8381 18015 8415
rect 17957 8375 18015 8381
rect 18233 8415 18291 8421
rect 18233 8381 18245 8415
rect 18279 8412 18291 8415
rect 18414 8412 18420 8424
rect 18279 8384 18420 8412
rect 18279 8381 18291 8384
rect 18233 8375 18291 8381
rect 17586 8304 17592 8356
rect 17644 8304 17650 8356
rect 17880 8344 17908 8375
rect 18414 8372 18420 8384
rect 18472 8372 18478 8424
rect 19981 8415 20039 8421
rect 19981 8381 19993 8415
rect 20027 8412 20039 8415
rect 20257 8415 20315 8421
rect 20257 8412 20269 8415
rect 20027 8384 20269 8412
rect 20027 8381 20039 8384
rect 19981 8375 20039 8381
rect 20257 8381 20269 8384
rect 20303 8412 20315 8415
rect 20714 8412 20720 8424
rect 20303 8384 20720 8412
rect 20303 8381 20315 8384
rect 20257 8375 20315 8381
rect 20714 8372 20720 8384
rect 20772 8372 20778 8424
rect 20993 8415 21051 8421
rect 20993 8381 21005 8415
rect 21039 8412 21051 8415
rect 21266 8412 21272 8424
rect 21039 8384 21272 8412
rect 21039 8381 21051 8384
rect 20993 8375 21051 8381
rect 21008 8344 21036 8375
rect 21266 8372 21272 8384
rect 21324 8372 21330 8424
rect 21361 8415 21419 8421
rect 21361 8381 21373 8415
rect 21407 8381 21419 8415
rect 21361 8375 21419 8381
rect 17880 8316 21036 8344
rect 21376 8344 21404 8375
rect 21450 8372 21456 8424
rect 21508 8372 21514 8424
rect 21910 8372 21916 8424
rect 21968 8372 21974 8424
rect 22112 8421 22140 8452
rect 22465 8449 22477 8452
rect 22511 8449 22523 8483
rect 22465 8443 22523 8449
rect 22097 8415 22155 8421
rect 22097 8381 22109 8415
rect 22143 8381 22155 8415
rect 22097 8375 22155 8381
rect 22186 8372 22192 8424
rect 22244 8372 22250 8424
rect 21928 8344 21956 8372
rect 21376 8316 21956 8344
rect 16224 8248 17080 8276
rect 17678 8236 17684 8288
rect 17736 8236 17742 8288
rect 17862 8236 17868 8288
rect 17920 8276 17926 8288
rect 19886 8276 19892 8288
rect 17920 8248 19892 8276
rect 17920 8236 17926 8248
rect 19886 8236 19892 8248
rect 19944 8236 19950 8288
rect 20070 8236 20076 8288
rect 20128 8236 20134 8288
rect 20346 8236 20352 8288
rect 20404 8276 20410 8288
rect 20530 8276 20536 8288
rect 20404 8248 20536 8276
rect 20404 8236 20410 8248
rect 20530 8236 20536 8248
rect 20588 8236 20594 8288
rect 20714 8236 20720 8288
rect 20772 8276 20778 8288
rect 20809 8279 20867 8285
rect 20809 8276 20821 8279
rect 20772 8248 20821 8276
rect 20772 8236 20778 8248
rect 20809 8245 20821 8248
rect 20855 8245 20867 8279
rect 20809 8239 20867 8245
rect 21082 8236 21088 8288
rect 21140 8276 21146 8288
rect 21634 8276 21640 8288
rect 21140 8248 21640 8276
rect 21140 8236 21146 8248
rect 21634 8236 21640 8248
rect 21692 8236 21698 8288
rect 21910 8236 21916 8288
rect 21968 8276 21974 8288
rect 22005 8279 22063 8285
rect 22005 8276 22017 8279
rect 21968 8248 22017 8276
rect 21968 8236 21974 8248
rect 22005 8245 22017 8248
rect 22051 8245 22063 8279
rect 22005 8239 22063 8245
rect 552 8186 23368 8208
rect 552 8134 4366 8186
rect 4418 8134 4430 8186
rect 4482 8134 4494 8186
rect 4546 8134 4558 8186
rect 4610 8134 4622 8186
rect 4674 8134 4686 8186
rect 4738 8134 10366 8186
rect 10418 8134 10430 8186
rect 10482 8134 10494 8186
rect 10546 8134 10558 8186
rect 10610 8134 10622 8186
rect 10674 8134 10686 8186
rect 10738 8134 16366 8186
rect 16418 8134 16430 8186
rect 16482 8134 16494 8186
rect 16546 8134 16558 8186
rect 16610 8134 16622 8186
rect 16674 8134 16686 8186
rect 16738 8134 22366 8186
rect 22418 8134 22430 8186
rect 22482 8134 22494 8186
rect 22546 8134 22558 8186
rect 22610 8134 22622 8186
rect 22674 8134 22686 8186
rect 22738 8134 23368 8186
rect 552 8112 23368 8134
rect 1762 8032 1768 8084
rect 1820 8072 1826 8084
rect 1949 8075 2007 8081
rect 1949 8072 1961 8075
rect 1820 8044 1961 8072
rect 1820 8032 1826 8044
rect 1949 8041 1961 8044
rect 1995 8041 2007 8075
rect 1949 8035 2007 8041
rect 2222 8032 2228 8084
rect 2280 8072 2286 8084
rect 2317 8075 2375 8081
rect 2317 8072 2329 8075
rect 2280 8044 2329 8072
rect 2280 8032 2286 8044
rect 2317 8041 2329 8044
rect 2363 8041 2375 8075
rect 8846 8072 8852 8084
rect 2317 8035 2375 8041
rect 2424 8044 4660 8072
rect 1673 8007 1731 8013
rect 1673 7973 1685 8007
rect 1719 8004 1731 8007
rect 1719 7976 2176 8004
rect 1719 7973 1731 7976
rect 1673 7967 1731 7973
rect 2148 7948 2176 7976
rect 1118 7896 1124 7948
rect 1176 7936 1182 7948
rect 1213 7939 1271 7945
rect 1213 7936 1225 7939
rect 1176 7908 1225 7936
rect 1176 7896 1182 7908
rect 1213 7905 1225 7908
rect 1259 7905 1271 7939
rect 1213 7899 1271 7905
rect 1854 7896 1860 7948
rect 1912 7896 1918 7948
rect 2130 7896 2136 7948
rect 2188 7896 2194 7948
rect 1302 7828 1308 7880
rect 1360 7828 1366 7880
rect 1489 7803 1547 7809
rect 1489 7769 1501 7803
rect 1535 7800 1547 7803
rect 2130 7800 2136 7812
rect 1535 7772 2136 7800
rect 1535 7769 1547 7772
rect 1489 7763 1547 7769
rect 2130 7760 2136 7772
rect 2188 7760 2194 7812
rect 842 7692 848 7744
rect 900 7692 906 7744
rect 1026 7692 1032 7744
rect 1084 7732 1090 7744
rect 2424 7732 2452 8044
rect 2516 7976 3096 8004
rect 2516 7948 2544 7976
rect 2498 7896 2504 7948
rect 2556 7896 2562 7948
rect 2682 7896 2688 7948
rect 2740 7896 2746 7948
rect 2774 7896 2780 7948
rect 2832 7896 2838 7948
rect 2866 7896 2872 7948
rect 2924 7896 2930 7948
rect 3068 7945 3096 7976
rect 3418 7964 3424 8016
rect 3476 8004 3482 8016
rect 3970 8004 3976 8016
rect 3476 7976 3976 8004
rect 3476 7964 3482 7976
rect 3970 7964 3976 7976
rect 4028 7964 4034 8016
rect 3053 7939 3111 7945
rect 3053 7905 3065 7939
rect 3099 7905 3111 7939
rect 3053 7899 3111 7905
rect 3142 7896 3148 7948
rect 3200 7896 3206 7948
rect 3326 7896 3332 7948
rect 3384 7936 3390 7948
rect 3602 7936 3608 7948
rect 3384 7908 3608 7936
rect 3384 7896 3390 7908
rect 3602 7896 3608 7908
rect 3660 7896 3666 7948
rect 4632 7945 4660 8044
rect 6748 8044 8852 8072
rect 4890 7964 4896 8016
rect 4948 8004 4954 8016
rect 4948 7976 6500 8004
rect 4948 7964 4954 7976
rect 4617 7939 4675 7945
rect 4617 7905 4629 7939
rect 4663 7905 4675 7939
rect 4617 7899 4675 7905
rect 5810 7896 5816 7948
rect 5868 7936 5874 7948
rect 6181 7939 6239 7945
rect 6181 7936 6193 7939
rect 5868 7908 6193 7936
rect 5868 7896 5874 7908
rect 6181 7905 6193 7908
rect 6227 7936 6239 7939
rect 6270 7936 6276 7948
rect 6227 7908 6276 7936
rect 6227 7905 6239 7908
rect 6181 7899 6239 7905
rect 6270 7896 6276 7908
rect 6328 7896 6334 7948
rect 6362 7896 6368 7948
rect 6420 7896 6426 7948
rect 6472 7945 6500 7976
rect 6546 7964 6552 8016
rect 6604 7964 6610 8016
rect 6457 7939 6515 7945
rect 6457 7905 6469 7939
rect 6503 7905 6515 7939
rect 6564 7936 6592 7964
rect 6748 7945 6776 8044
rect 8846 8032 8852 8044
rect 8904 8032 8910 8084
rect 9030 8032 9036 8084
rect 9088 8032 9094 8084
rect 9214 8032 9220 8084
rect 9272 8072 9278 8084
rect 9272 8044 9720 8072
rect 9272 8032 9278 8044
rect 6822 7964 6828 8016
rect 6880 8004 6886 8016
rect 6880 7976 7972 8004
rect 6880 7964 6886 7976
rect 6641 7939 6699 7945
rect 6641 7936 6653 7939
rect 6564 7908 6653 7936
rect 6457 7899 6515 7905
rect 6641 7905 6653 7908
rect 6687 7905 6699 7939
rect 6641 7899 6699 7905
rect 6733 7939 6791 7945
rect 6733 7905 6745 7939
rect 6779 7905 6791 7939
rect 6733 7899 6791 7905
rect 6914 7896 6920 7948
rect 6972 7896 6978 7948
rect 7190 7896 7196 7948
rect 7248 7896 7254 7948
rect 7285 7939 7343 7945
rect 7285 7905 7297 7939
rect 7331 7936 7343 7939
rect 7331 7908 7512 7936
rect 7331 7905 7343 7908
rect 7285 7899 7343 7905
rect 2792 7800 2820 7896
rect 2958 7828 2964 7880
rect 3016 7868 3022 7880
rect 3513 7871 3571 7877
rect 3513 7868 3525 7871
rect 3016 7840 3525 7868
rect 3016 7828 3022 7840
rect 3513 7837 3525 7840
rect 3559 7837 3571 7871
rect 3513 7831 3571 7837
rect 4709 7871 4767 7877
rect 4709 7837 4721 7871
rect 4755 7868 4767 7871
rect 4798 7868 4804 7880
rect 4755 7840 4804 7868
rect 4755 7837 4767 7840
rect 4709 7831 4767 7837
rect 4798 7828 4804 7840
rect 4856 7828 4862 7880
rect 6549 7871 6607 7877
rect 6549 7837 6561 7871
rect 6595 7868 6607 7871
rect 7009 7871 7067 7877
rect 7009 7868 7021 7871
rect 6595 7840 7021 7868
rect 6595 7837 6607 7840
rect 6549 7831 6607 7837
rect 7009 7837 7021 7840
rect 7055 7837 7067 7871
rect 7009 7831 7067 7837
rect 7101 7871 7159 7877
rect 7101 7837 7113 7871
rect 7147 7837 7159 7871
rect 7208 7868 7236 7896
rect 7484 7868 7512 7908
rect 7558 7896 7564 7948
rect 7616 7896 7622 7948
rect 7834 7896 7840 7948
rect 7892 7896 7898 7948
rect 7944 7945 7972 7976
rect 7929 7939 7987 7945
rect 7929 7905 7941 7939
rect 7975 7905 7987 7939
rect 9048 7936 9076 8032
rect 7929 7899 7987 7905
rect 8036 7908 9076 7936
rect 9125 7939 9183 7945
rect 8036 7868 8064 7908
rect 9125 7905 9137 7939
rect 9171 7905 9183 7939
rect 9125 7899 9183 7905
rect 7208 7840 7328 7868
rect 7484 7840 8064 7868
rect 8849 7871 8907 7877
rect 7101 7831 7159 7837
rect 2869 7803 2927 7809
rect 2869 7800 2881 7803
rect 2792 7772 2881 7800
rect 2869 7769 2881 7772
rect 2915 7800 2927 7803
rect 3050 7800 3056 7812
rect 2915 7772 3056 7800
rect 2915 7769 2927 7772
rect 2869 7763 2927 7769
rect 3050 7760 3056 7772
rect 3108 7760 3114 7812
rect 4985 7803 5043 7809
rect 4985 7769 4997 7803
rect 5031 7800 5043 7803
rect 5074 7800 5080 7812
rect 5031 7772 5080 7800
rect 5031 7769 5043 7772
rect 4985 7763 5043 7769
rect 5074 7760 5080 7772
rect 5132 7760 5138 7812
rect 7116 7800 7144 7831
rect 7190 7800 7196 7812
rect 6196 7772 7196 7800
rect 1084 7704 2452 7732
rect 3329 7735 3387 7741
rect 1084 7692 1090 7704
rect 3329 7701 3341 7735
rect 3375 7732 3387 7735
rect 3418 7732 3424 7744
rect 3375 7704 3424 7732
rect 3375 7701 3387 7704
rect 3329 7695 3387 7701
rect 3418 7692 3424 7704
rect 3476 7692 3482 7744
rect 3881 7735 3939 7741
rect 3881 7701 3893 7735
rect 3927 7732 3939 7735
rect 6196 7732 6224 7772
rect 7190 7760 7196 7772
rect 7248 7760 7254 7812
rect 7300 7800 7328 7840
rect 7944 7812 7972 7840
rect 8849 7837 8861 7871
rect 8895 7868 8907 7871
rect 8938 7868 8944 7880
rect 8895 7840 8944 7868
rect 8895 7837 8907 7840
rect 8849 7831 8907 7837
rect 7653 7803 7711 7809
rect 7653 7800 7665 7803
rect 7300 7772 7665 7800
rect 7653 7769 7665 7772
rect 7699 7769 7711 7803
rect 7653 7763 7711 7769
rect 7926 7760 7932 7812
rect 7984 7760 7990 7812
rect 8864 7800 8892 7831
rect 8938 7828 8944 7840
rect 8996 7828 9002 7880
rect 9140 7812 9168 7899
rect 9214 7896 9220 7948
rect 9272 7936 9278 7948
rect 9398 7936 9404 7948
rect 9272 7908 9404 7936
rect 9272 7896 9278 7908
rect 9398 7896 9404 7908
rect 9456 7896 9462 7948
rect 9490 7828 9496 7880
rect 9548 7828 9554 7880
rect 9692 7868 9720 8044
rect 10502 8032 10508 8084
rect 10560 8072 10566 8084
rect 11698 8072 11704 8084
rect 10560 8044 11704 8072
rect 10560 8032 10566 8044
rect 11698 8032 11704 8044
rect 11756 8072 11762 8084
rect 12345 8075 12403 8081
rect 11756 8044 12020 8072
rect 11756 8032 11762 8044
rect 11790 8004 11796 8016
rect 9968 7976 11796 8004
rect 9766 7896 9772 7948
rect 9824 7936 9830 7948
rect 9968 7945 9996 7976
rect 11790 7964 11796 7976
rect 11848 7964 11854 8016
rect 11992 8013 12020 8044
rect 12345 8041 12357 8075
rect 12391 8072 12403 8075
rect 12434 8072 12440 8084
rect 12391 8044 12440 8072
rect 12391 8041 12403 8044
rect 12345 8035 12403 8041
rect 12434 8032 12440 8044
rect 12492 8032 12498 8084
rect 12802 8032 12808 8084
rect 12860 8072 12866 8084
rect 12860 8044 14780 8072
rect 12860 8032 12866 8044
rect 11977 8007 12035 8013
rect 11977 7973 11989 8007
rect 12023 7973 12035 8007
rect 11977 7967 12035 7973
rect 12158 7964 12164 8016
rect 12216 7964 12222 8016
rect 14752 8004 14780 8044
rect 15286 8032 15292 8084
rect 15344 8072 15350 8084
rect 15473 8075 15531 8081
rect 15473 8072 15485 8075
rect 15344 8044 15485 8072
rect 15344 8032 15350 8044
rect 15473 8041 15485 8044
rect 15519 8041 15531 8075
rect 15473 8035 15531 8041
rect 18616 8044 20116 8072
rect 17862 8004 17868 8016
rect 14752 7976 17868 8004
rect 17862 7964 17868 7976
rect 17920 7964 17926 8016
rect 9861 7939 9919 7945
rect 9861 7936 9873 7939
rect 9824 7908 9873 7936
rect 9824 7896 9830 7908
rect 9861 7905 9873 7908
rect 9907 7905 9919 7939
rect 9861 7899 9919 7905
rect 9953 7939 10011 7945
rect 9953 7905 9965 7939
rect 9999 7905 10011 7939
rect 9953 7899 10011 7905
rect 10229 7939 10287 7945
rect 10229 7905 10241 7939
rect 10275 7905 10287 7939
rect 10229 7899 10287 7905
rect 10244 7868 10272 7899
rect 10318 7896 10324 7948
rect 10376 7896 10382 7948
rect 10502 7896 10508 7948
rect 10560 7896 10566 7948
rect 10689 7939 10747 7945
rect 10689 7905 10701 7939
rect 10735 7936 10747 7939
rect 10965 7939 11023 7945
rect 10965 7936 10977 7939
rect 10735 7908 10977 7936
rect 10735 7905 10747 7908
rect 10689 7899 10747 7905
rect 10965 7905 10977 7908
rect 11011 7905 11023 7939
rect 10965 7899 11023 7905
rect 11149 7939 11207 7945
rect 11149 7905 11161 7939
rect 11195 7905 11207 7939
rect 11149 7899 11207 7905
rect 11241 7939 11299 7945
rect 11241 7905 11253 7939
rect 11287 7936 11299 7939
rect 11517 7939 11575 7945
rect 11287 7908 11468 7936
rect 11287 7905 11299 7908
rect 11241 7899 11299 7905
rect 10870 7868 10876 7880
rect 9692 7840 10876 7868
rect 10870 7828 10876 7840
rect 10928 7828 10934 7880
rect 11054 7828 11060 7880
rect 11112 7828 11118 7880
rect 8036 7772 8892 7800
rect 3927 7704 6224 7732
rect 3927 7701 3939 7704
rect 3881 7695 3939 7701
rect 6270 7692 6276 7744
rect 6328 7692 6334 7744
rect 7466 7692 7472 7744
rect 7524 7692 7530 7744
rect 7558 7692 7564 7744
rect 7616 7732 7622 7744
rect 8036 7732 8064 7772
rect 9122 7760 9128 7812
rect 9180 7760 9186 7812
rect 9309 7803 9367 7809
rect 9309 7769 9321 7803
rect 9355 7800 9367 7803
rect 9582 7800 9588 7812
rect 9355 7772 9588 7800
rect 9355 7769 9367 7772
rect 9309 7763 9367 7769
rect 9582 7760 9588 7772
rect 9640 7760 9646 7812
rect 10137 7803 10195 7809
rect 10137 7769 10149 7803
rect 10183 7800 10195 7803
rect 11072 7800 11100 7828
rect 11164 7812 11192 7899
rect 11330 7828 11336 7880
rect 11388 7828 11394 7880
rect 11440 7868 11468 7908
rect 11517 7905 11529 7939
rect 11563 7936 11575 7939
rect 11882 7936 11888 7948
rect 11563 7908 11888 7936
rect 11563 7905 11575 7908
rect 11517 7899 11575 7905
rect 11882 7896 11888 7908
rect 11940 7896 11946 7948
rect 13538 7896 13544 7948
rect 13596 7936 13602 7948
rect 14277 7939 14335 7945
rect 14277 7936 14289 7939
rect 13596 7908 14289 7936
rect 13596 7896 13602 7908
rect 14277 7905 14289 7908
rect 14323 7936 14335 7939
rect 14645 7939 14703 7945
rect 14645 7936 14657 7939
rect 14323 7908 14657 7936
rect 14323 7905 14335 7908
rect 14277 7899 14335 7905
rect 14645 7905 14657 7908
rect 14691 7905 14703 7939
rect 14645 7899 14703 7905
rect 15654 7896 15660 7948
rect 15712 7896 15718 7948
rect 15749 7939 15807 7945
rect 15749 7905 15761 7939
rect 15795 7936 15807 7939
rect 16022 7936 16028 7948
rect 15795 7908 16028 7936
rect 15795 7905 15807 7908
rect 15749 7899 15807 7905
rect 16022 7896 16028 7908
rect 16080 7936 16086 7948
rect 17218 7936 17224 7948
rect 16080 7908 17224 7936
rect 16080 7896 16086 7908
rect 17218 7896 17224 7908
rect 17276 7896 17282 7948
rect 17954 7896 17960 7948
rect 18012 7936 18018 7948
rect 18141 7939 18199 7945
rect 18141 7936 18153 7939
rect 18012 7908 18153 7936
rect 18012 7896 18018 7908
rect 18141 7905 18153 7908
rect 18187 7905 18199 7939
rect 18509 7939 18567 7945
rect 18509 7936 18521 7939
rect 18141 7899 18199 7905
rect 18248 7908 18521 7936
rect 11698 7868 11704 7880
rect 11440 7840 11704 7868
rect 11698 7828 11704 7840
rect 11756 7828 11762 7880
rect 14553 7871 14611 7877
rect 14553 7837 14565 7871
rect 14599 7860 14611 7871
rect 14826 7868 14832 7880
rect 14660 7860 14832 7868
rect 14599 7840 14832 7860
rect 14599 7837 14688 7840
rect 14553 7832 14688 7837
rect 14553 7831 14611 7832
rect 14826 7828 14832 7840
rect 14884 7828 14890 7880
rect 14921 7871 14979 7877
rect 14921 7837 14933 7871
rect 14967 7868 14979 7871
rect 17034 7868 17040 7880
rect 14967 7840 17040 7868
rect 14967 7837 14979 7840
rect 14921 7831 14979 7837
rect 17034 7828 17040 7840
rect 17092 7828 17098 7880
rect 10183 7772 11100 7800
rect 10183 7769 10195 7772
rect 10137 7763 10195 7769
rect 11146 7760 11152 7812
rect 11204 7800 11210 7812
rect 14090 7800 14096 7812
rect 11204 7772 14096 7800
rect 11204 7760 11210 7772
rect 14090 7760 14096 7772
rect 14148 7760 14154 7812
rect 14461 7803 14519 7809
rect 14461 7769 14473 7803
rect 14507 7800 14519 7803
rect 15102 7800 15108 7812
rect 14507 7772 15108 7800
rect 14507 7769 14519 7772
rect 14461 7763 14519 7769
rect 15102 7760 15108 7772
rect 15160 7760 15166 7812
rect 15654 7760 15660 7812
rect 15712 7800 15718 7812
rect 18248 7800 18276 7908
rect 18509 7905 18521 7908
rect 18555 7936 18567 7939
rect 18616 7936 18644 8044
rect 19150 7964 19156 8016
rect 19208 7964 19214 8016
rect 20088 8004 20116 8044
rect 20162 8032 20168 8084
rect 20220 8072 20226 8084
rect 20530 8072 20536 8084
rect 20220 8044 20536 8072
rect 20220 8032 20226 8044
rect 20530 8032 20536 8044
rect 20588 8072 20594 8084
rect 21469 8075 21527 8081
rect 21469 8072 21481 8075
rect 20588 8044 21481 8072
rect 20588 8032 20594 8044
rect 21469 8041 21481 8044
rect 21515 8041 21527 8075
rect 21469 8035 21527 8041
rect 20714 8004 20720 8016
rect 20088 7976 20720 8004
rect 20714 7964 20720 7976
rect 20772 7964 20778 8016
rect 21174 7964 21180 8016
rect 21232 8004 21238 8016
rect 21269 8007 21327 8013
rect 21269 8004 21281 8007
rect 21232 7976 21281 8004
rect 21232 7964 21238 7976
rect 21269 7973 21281 7976
rect 21315 7973 21327 8007
rect 21269 7967 21327 7973
rect 18555 7908 18644 7936
rect 18555 7905 18567 7908
rect 18509 7899 18567 7905
rect 18690 7896 18696 7948
rect 18748 7896 18754 7948
rect 18874 7896 18880 7948
rect 18932 7936 18938 7948
rect 18969 7939 19027 7945
rect 18969 7936 18981 7939
rect 18932 7908 18981 7936
rect 18932 7896 18938 7908
rect 18969 7905 18981 7908
rect 19015 7905 19027 7939
rect 18969 7899 19027 7905
rect 19245 7939 19303 7945
rect 19245 7905 19257 7939
rect 19291 7905 19303 7939
rect 19245 7899 19303 7905
rect 19521 7939 19579 7945
rect 19521 7905 19533 7939
rect 19567 7936 19579 7939
rect 19610 7936 19616 7948
rect 19567 7908 19616 7936
rect 19567 7905 19579 7908
rect 19521 7899 19579 7905
rect 18325 7871 18383 7877
rect 18325 7837 18337 7871
rect 18371 7837 18383 7871
rect 18325 7831 18383 7837
rect 15712 7772 18276 7800
rect 18340 7800 18368 7831
rect 18414 7828 18420 7880
rect 18472 7828 18478 7880
rect 19260 7868 19288 7899
rect 19610 7896 19616 7908
rect 19668 7896 19674 7948
rect 19702 7896 19708 7948
rect 19760 7896 19766 7948
rect 19797 7939 19855 7945
rect 19797 7905 19809 7939
rect 19843 7936 19855 7939
rect 21910 7936 21916 7948
rect 19843 7908 21916 7936
rect 19843 7905 19855 7908
rect 19797 7899 19855 7905
rect 19812 7868 19840 7899
rect 21910 7896 21916 7908
rect 21968 7896 21974 7948
rect 19260 7840 19840 7868
rect 20070 7800 20076 7812
rect 18340 7772 20076 7800
rect 15712 7760 15718 7772
rect 20070 7760 20076 7772
rect 20128 7760 20134 7812
rect 7616 7704 8064 7732
rect 8113 7735 8171 7741
rect 7616 7692 7622 7704
rect 8113 7701 8125 7735
rect 8159 7732 8171 7735
rect 8202 7732 8208 7744
rect 8159 7704 8208 7732
rect 8159 7701 8171 7704
rect 8113 7695 8171 7701
rect 8202 7692 8208 7704
rect 8260 7692 8266 7744
rect 9398 7692 9404 7744
rect 9456 7692 9462 7744
rect 9674 7692 9680 7744
rect 9732 7692 9738 7744
rect 11054 7692 11060 7744
rect 11112 7732 11118 7744
rect 11701 7735 11759 7741
rect 11701 7732 11713 7735
rect 11112 7704 11713 7732
rect 11112 7692 11118 7704
rect 11701 7701 11713 7704
rect 11747 7701 11759 7735
rect 11701 7695 11759 7701
rect 11790 7692 11796 7744
rect 11848 7732 11854 7744
rect 14369 7735 14427 7741
rect 14369 7732 14381 7735
rect 11848 7704 14381 7732
rect 11848 7692 11854 7704
rect 14369 7701 14381 7704
rect 14415 7732 14427 7735
rect 14550 7732 14556 7744
rect 14415 7704 14556 7732
rect 14415 7701 14427 7704
rect 14369 7695 14427 7701
rect 14550 7692 14556 7704
rect 14608 7692 14614 7744
rect 14734 7692 14740 7744
rect 14792 7692 14798 7744
rect 14826 7692 14832 7744
rect 14884 7692 14890 7744
rect 15286 7692 15292 7744
rect 15344 7732 15350 7744
rect 15746 7732 15752 7744
rect 15344 7704 15752 7732
rect 15344 7692 15350 7704
rect 15746 7692 15752 7704
rect 15804 7692 15810 7744
rect 15838 7692 15844 7744
rect 15896 7732 15902 7744
rect 15933 7735 15991 7741
rect 15933 7732 15945 7735
rect 15896 7704 15945 7732
rect 15896 7692 15902 7704
rect 15933 7701 15945 7704
rect 15979 7701 15991 7735
rect 15933 7695 15991 7701
rect 17954 7692 17960 7744
rect 18012 7692 18018 7744
rect 18782 7692 18788 7744
rect 18840 7692 18846 7744
rect 18874 7692 18880 7744
rect 18932 7732 18938 7744
rect 19337 7735 19395 7741
rect 19337 7732 19349 7735
rect 18932 7704 19349 7732
rect 18932 7692 18938 7704
rect 19337 7701 19349 7704
rect 19383 7701 19395 7735
rect 19337 7695 19395 7701
rect 19886 7692 19892 7744
rect 19944 7732 19950 7744
rect 20162 7732 20168 7744
rect 19944 7704 20168 7732
rect 19944 7692 19950 7704
rect 20162 7692 20168 7704
rect 20220 7692 20226 7744
rect 20990 7692 20996 7744
rect 21048 7732 21054 7744
rect 21453 7735 21511 7741
rect 21453 7732 21465 7735
rect 21048 7704 21465 7732
rect 21048 7692 21054 7704
rect 21453 7701 21465 7704
rect 21499 7701 21511 7735
rect 21453 7695 21511 7701
rect 21637 7735 21695 7741
rect 21637 7701 21649 7735
rect 21683 7732 21695 7735
rect 22278 7732 22284 7744
rect 21683 7704 22284 7732
rect 21683 7701 21695 7704
rect 21637 7695 21695 7701
rect 22278 7692 22284 7704
rect 22336 7692 22342 7744
rect 552 7642 23368 7664
rect 552 7590 1366 7642
rect 1418 7590 1430 7642
rect 1482 7590 1494 7642
rect 1546 7590 1558 7642
rect 1610 7590 1622 7642
rect 1674 7590 1686 7642
rect 1738 7590 7366 7642
rect 7418 7590 7430 7642
rect 7482 7590 7494 7642
rect 7546 7590 7558 7642
rect 7610 7590 7622 7642
rect 7674 7590 7686 7642
rect 7738 7590 13366 7642
rect 13418 7590 13430 7642
rect 13482 7590 13494 7642
rect 13546 7590 13558 7642
rect 13610 7590 13622 7642
rect 13674 7590 13686 7642
rect 13738 7590 19366 7642
rect 19418 7590 19430 7642
rect 19482 7590 19494 7642
rect 19546 7590 19558 7642
rect 19610 7590 19622 7642
rect 19674 7590 19686 7642
rect 19738 7590 23368 7642
rect 552 7568 23368 7590
rect 1305 7531 1363 7537
rect 1305 7497 1317 7531
rect 1351 7528 1363 7531
rect 1946 7528 1952 7540
rect 1351 7500 1952 7528
rect 1351 7497 1363 7500
rect 1305 7491 1363 7497
rect 1946 7488 1952 7500
rect 2004 7488 2010 7540
rect 2133 7531 2191 7537
rect 2133 7497 2145 7531
rect 2179 7528 2191 7531
rect 2498 7528 2504 7540
rect 2179 7500 2504 7528
rect 2179 7497 2191 7500
rect 2133 7491 2191 7497
rect 2498 7488 2504 7500
rect 2556 7488 2562 7540
rect 6730 7488 6736 7540
rect 6788 7528 6794 7540
rect 7101 7531 7159 7537
rect 7101 7528 7113 7531
rect 6788 7500 7113 7528
rect 6788 7488 6794 7500
rect 7101 7497 7113 7500
rect 7147 7497 7159 7531
rect 7101 7491 7159 7497
rect 7190 7488 7196 7540
rect 7248 7488 7254 7540
rect 8386 7488 8392 7540
rect 8444 7528 8450 7540
rect 10502 7528 10508 7540
rect 8444 7500 10508 7528
rect 8444 7488 8450 7500
rect 10502 7488 10508 7500
rect 10560 7488 10566 7540
rect 10870 7488 10876 7540
rect 10928 7528 10934 7540
rect 11606 7528 11612 7540
rect 10928 7500 11612 7528
rect 10928 7488 10934 7500
rect 11606 7488 11612 7500
rect 11664 7488 11670 7540
rect 15838 7528 15844 7540
rect 12406 7500 15844 7528
rect 3326 7420 3332 7472
rect 3384 7460 3390 7472
rect 5166 7460 5172 7472
rect 3384 7432 5172 7460
rect 3384 7420 3390 7432
rect 5166 7420 5172 7432
rect 5224 7420 5230 7472
rect 6914 7420 6920 7472
rect 6972 7420 6978 7472
rect 9122 7420 9128 7472
rect 9180 7420 9186 7472
rect 9217 7463 9275 7469
rect 9217 7429 9229 7463
rect 9263 7460 9275 7463
rect 11333 7463 11391 7469
rect 11333 7460 11345 7463
rect 9263 7432 11345 7460
rect 9263 7429 9275 7432
rect 9217 7423 9275 7429
rect 11333 7429 11345 7432
rect 11379 7460 11391 7463
rect 12406 7460 12434 7500
rect 15838 7488 15844 7500
rect 15896 7488 15902 7540
rect 16666 7488 16672 7540
rect 16724 7528 16730 7540
rect 17126 7528 17132 7540
rect 16724 7500 17132 7528
rect 16724 7488 16730 7500
rect 17126 7488 17132 7500
rect 17184 7528 17190 7540
rect 19794 7528 19800 7540
rect 17184 7500 19800 7528
rect 17184 7488 17190 7500
rect 19794 7488 19800 7500
rect 19852 7488 19858 7540
rect 21450 7528 21456 7540
rect 20088 7500 21456 7528
rect 14734 7460 14740 7472
rect 11379 7432 12434 7460
rect 12912 7432 14740 7460
rect 11379 7429 11391 7432
rect 11333 7423 11391 7429
rect 1762 7352 1768 7404
rect 1820 7352 1826 7404
rect 2777 7395 2835 7401
rect 2777 7361 2789 7395
rect 2823 7392 2835 7395
rect 2958 7392 2964 7404
rect 2823 7364 2964 7392
rect 2823 7361 2835 7364
rect 2777 7355 2835 7361
rect 2958 7352 2964 7364
rect 3016 7352 3022 7404
rect 3053 7395 3111 7401
rect 3053 7361 3065 7395
rect 3099 7392 3111 7395
rect 3142 7392 3148 7404
rect 3099 7364 3148 7392
rect 3099 7361 3111 7364
rect 3053 7355 3111 7361
rect 3142 7352 3148 7364
rect 3200 7352 3206 7404
rect 3418 7392 3424 7404
rect 3252 7364 3424 7392
rect 1029 7327 1087 7333
rect 1029 7293 1041 7327
rect 1075 7324 1087 7327
rect 1118 7324 1124 7336
rect 1075 7296 1124 7324
rect 1075 7293 1087 7296
rect 1029 7287 1087 7293
rect 1118 7284 1124 7296
rect 1176 7284 1182 7336
rect 1486 7284 1492 7336
rect 1544 7284 1550 7336
rect 1949 7327 2007 7333
rect 1949 7293 1961 7327
rect 1995 7324 2007 7327
rect 3252 7324 3280 7364
rect 3418 7352 3424 7364
rect 3476 7352 3482 7404
rect 3602 7352 3608 7404
rect 3660 7352 3666 7404
rect 3878 7352 3884 7404
rect 3936 7392 3942 7404
rect 5905 7395 5963 7401
rect 5905 7392 5917 7395
rect 3936 7364 5917 7392
rect 3936 7352 3942 7364
rect 5905 7361 5917 7364
rect 5951 7361 5963 7395
rect 5905 7355 5963 7361
rect 6086 7352 6092 7404
rect 6144 7392 6150 7404
rect 7009 7395 7067 7401
rect 6144 7364 6224 7392
rect 6144 7352 6150 7364
rect 1995 7296 3280 7324
rect 3329 7327 3387 7333
rect 1995 7293 2007 7296
rect 1949 7287 2007 7293
rect 3329 7293 3341 7327
rect 3375 7293 3387 7327
rect 3329 7287 3387 7293
rect 2130 7256 2136 7268
rect 1136 7228 2136 7256
rect 1136 7197 1164 7228
rect 2130 7216 2136 7228
rect 2188 7216 2194 7268
rect 1121 7191 1179 7197
rect 1121 7157 1133 7191
rect 1167 7157 1179 7191
rect 1121 7151 1179 7157
rect 1854 7148 1860 7200
rect 1912 7188 1918 7200
rect 3344 7188 3372 7287
rect 4246 7284 4252 7336
rect 4304 7324 4310 7336
rect 4433 7327 4491 7333
rect 4433 7324 4445 7327
rect 4304 7296 4445 7324
rect 4304 7284 4310 7296
rect 4433 7293 4445 7296
rect 4479 7293 4491 7327
rect 4433 7287 4491 7293
rect 4617 7327 4675 7333
rect 4617 7293 4629 7327
rect 4663 7324 4675 7327
rect 4890 7324 4896 7336
rect 4663 7296 4896 7324
rect 4663 7293 4675 7296
rect 4617 7287 4675 7293
rect 4890 7284 4896 7296
rect 4948 7284 4954 7336
rect 5261 7327 5319 7333
rect 5261 7293 5273 7327
rect 5307 7324 5319 7327
rect 5350 7324 5356 7336
rect 5307 7296 5356 7324
rect 5307 7293 5319 7296
rect 5261 7287 5319 7293
rect 5350 7284 5356 7296
rect 5408 7284 5414 7336
rect 5537 7327 5595 7333
rect 5537 7293 5549 7327
rect 5583 7324 5595 7327
rect 5810 7324 5816 7336
rect 5583 7296 5816 7324
rect 5583 7293 5595 7296
rect 5537 7287 5595 7293
rect 5810 7284 5816 7296
rect 5868 7284 5874 7336
rect 5994 7284 6000 7336
rect 6052 7284 6058 7336
rect 6196 7321 6224 7364
rect 7009 7361 7021 7395
rect 7055 7392 7067 7395
rect 7190 7392 7196 7404
rect 7055 7364 7196 7392
rect 7055 7361 7067 7364
rect 7009 7355 7067 7361
rect 7190 7352 7196 7364
rect 7248 7352 7254 7404
rect 7742 7352 7748 7404
rect 7800 7392 7806 7404
rect 9140 7392 9168 7420
rect 7800 7364 8708 7392
rect 7800 7352 7806 7364
rect 6368 7327 6426 7333
rect 6368 7324 6380 7327
rect 6347 7321 6380 7324
rect 6196 7293 6380 7321
rect 6414 7293 6426 7327
rect 6368 7287 6426 7293
rect 6730 7284 6736 7336
rect 6788 7284 6794 7336
rect 6917 7327 6975 7333
rect 6917 7293 6929 7327
rect 6963 7293 6975 7327
rect 6917 7287 6975 7293
rect 6822 7256 6828 7268
rect 6380 7228 6828 7256
rect 1912 7160 3372 7188
rect 4525 7191 4583 7197
rect 1912 7148 1918 7160
rect 4525 7157 4537 7191
rect 4571 7188 4583 7191
rect 4798 7188 4804 7200
rect 4571 7160 4804 7188
rect 4571 7157 4583 7160
rect 4525 7151 4583 7157
rect 4798 7148 4804 7160
rect 4856 7148 4862 7200
rect 5166 7148 5172 7200
rect 5224 7188 5230 7200
rect 5353 7191 5411 7197
rect 5353 7188 5365 7191
rect 5224 7160 5365 7188
rect 5224 7148 5230 7160
rect 5353 7157 5365 7160
rect 5399 7157 5411 7191
rect 5353 7151 5411 7157
rect 5718 7148 5724 7200
rect 5776 7148 5782 7200
rect 6380 7197 6408 7228
rect 6822 7216 6828 7228
rect 6880 7216 6886 7268
rect 6932 7256 6960 7287
rect 7282 7284 7288 7336
rect 7340 7284 7346 7336
rect 7561 7327 7619 7333
rect 7561 7293 7573 7327
rect 7607 7293 7619 7327
rect 7561 7287 7619 7293
rect 7098 7256 7104 7268
rect 6932 7228 7104 7256
rect 7098 7216 7104 7228
rect 7156 7216 7162 7268
rect 7576 7256 7604 7287
rect 7650 7284 7656 7336
rect 7708 7324 7714 7336
rect 7837 7327 7895 7333
rect 7837 7324 7849 7327
rect 7708 7296 7849 7324
rect 7708 7284 7714 7296
rect 7837 7293 7849 7296
rect 7883 7293 7895 7327
rect 7837 7287 7895 7293
rect 8386 7284 8392 7336
rect 8444 7284 8450 7336
rect 8680 7333 8708 7364
rect 8772 7364 9168 7392
rect 9401 7395 9459 7401
rect 8772 7333 8800 7364
rect 9401 7361 9413 7395
rect 9447 7392 9459 7395
rect 9674 7392 9680 7404
rect 9447 7364 9680 7392
rect 9447 7361 9459 7364
rect 9401 7355 9459 7361
rect 9674 7352 9680 7364
rect 9732 7352 9738 7404
rect 9766 7352 9772 7404
rect 9824 7392 9830 7404
rect 10962 7392 10968 7404
rect 9824 7364 10968 7392
rect 9824 7352 9830 7364
rect 10962 7352 10968 7364
rect 11020 7392 11026 7404
rect 11020 7364 11376 7392
rect 11020 7352 11026 7364
rect 8573 7327 8631 7333
rect 8573 7293 8585 7327
rect 8619 7293 8631 7327
rect 8573 7287 8631 7293
rect 8665 7327 8723 7333
rect 8665 7293 8677 7327
rect 8711 7293 8723 7327
rect 8665 7287 8723 7293
rect 8757 7327 8815 7333
rect 8757 7293 8769 7327
rect 8803 7293 8815 7327
rect 8757 7287 8815 7293
rect 9125 7327 9183 7333
rect 9125 7293 9137 7327
rect 9171 7324 9183 7327
rect 9214 7324 9220 7336
rect 9171 7296 9220 7324
rect 9171 7293 9183 7296
rect 9125 7287 9183 7293
rect 8110 7256 8116 7268
rect 7576 7228 8116 7256
rect 8110 7216 8116 7228
rect 8168 7216 8174 7268
rect 6365 7191 6423 7197
rect 6365 7157 6377 7191
rect 6411 7157 6423 7191
rect 6365 7151 6423 7157
rect 6546 7148 6552 7200
rect 6604 7148 6610 7200
rect 7190 7148 7196 7200
rect 7248 7188 7254 7200
rect 7377 7191 7435 7197
rect 7377 7188 7389 7191
rect 7248 7160 7389 7188
rect 7248 7148 7254 7160
rect 7377 7157 7389 7160
rect 7423 7157 7435 7191
rect 7377 7151 7435 7157
rect 7466 7148 7472 7200
rect 7524 7188 7530 7200
rect 8588 7188 8616 7287
rect 9214 7284 9220 7296
rect 9272 7284 9278 7336
rect 10042 7284 10048 7336
rect 10100 7324 10106 7336
rect 10229 7327 10287 7333
rect 10229 7324 10241 7327
rect 10100 7296 10241 7324
rect 10100 7284 10106 7296
rect 10229 7293 10241 7296
rect 10275 7293 10287 7327
rect 10229 7287 10287 7293
rect 11241 7327 11299 7333
rect 11241 7293 11253 7327
rect 11287 7293 11299 7327
rect 11348 7324 11376 7364
rect 11514 7352 11520 7404
rect 11572 7352 11578 7404
rect 11606 7352 11612 7404
rect 11664 7392 11670 7404
rect 12912 7392 12940 7432
rect 14734 7420 14740 7432
rect 14792 7460 14798 7472
rect 16853 7463 16911 7469
rect 16853 7460 16865 7463
rect 14792 7432 16865 7460
rect 14792 7420 14798 7432
rect 16853 7429 16865 7432
rect 16899 7460 16911 7463
rect 18233 7463 18291 7469
rect 18233 7460 18245 7463
rect 16899 7432 18245 7460
rect 16899 7429 16911 7432
rect 16853 7423 16911 7429
rect 18233 7429 18245 7432
rect 18279 7429 18291 7463
rect 18233 7423 18291 7429
rect 18690 7420 18696 7472
rect 18748 7460 18754 7472
rect 20088 7460 20116 7500
rect 21450 7488 21456 7500
rect 21508 7488 21514 7540
rect 21542 7488 21548 7540
rect 21600 7528 21606 7540
rect 21637 7531 21695 7537
rect 21637 7528 21649 7531
rect 21600 7500 21649 7528
rect 21600 7488 21606 7500
rect 21637 7497 21649 7500
rect 21683 7497 21695 7531
rect 21637 7491 21695 7497
rect 18748 7432 20116 7460
rect 18748 7420 18754 7432
rect 11664 7364 12940 7392
rect 11664 7352 11670 7364
rect 12986 7352 12992 7404
rect 13044 7392 13050 7404
rect 13817 7395 13875 7401
rect 13817 7392 13829 7395
rect 13044 7364 13829 7392
rect 13044 7352 13050 7364
rect 13817 7361 13829 7364
rect 13863 7361 13875 7395
rect 13817 7355 13875 7361
rect 14458 7352 14464 7404
rect 14516 7392 14522 7404
rect 17037 7395 17095 7401
rect 14516 7364 14596 7392
rect 14516 7352 14522 7364
rect 11790 7324 11796 7336
rect 11348 7296 11796 7324
rect 11241 7287 11299 7293
rect 10134 7256 10140 7268
rect 9048 7228 10140 7256
rect 9048 7197 9076 7228
rect 10134 7216 10140 7228
rect 10192 7216 10198 7268
rect 11256 7256 11284 7287
rect 11790 7284 11796 7296
rect 11848 7284 11854 7336
rect 11698 7256 11704 7268
rect 10428 7228 11704 7256
rect 7524 7160 8616 7188
rect 9033 7191 9091 7197
rect 7524 7148 7530 7160
rect 9033 7157 9045 7191
rect 9079 7157 9091 7191
rect 9033 7151 9091 7157
rect 9122 7148 9128 7200
rect 9180 7188 9186 7200
rect 10428 7197 10456 7228
rect 11698 7216 11704 7228
rect 11756 7256 11762 7268
rect 13004 7256 13032 7352
rect 13630 7284 13636 7336
rect 13688 7284 13694 7336
rect 13725 7327 13783 7333
rect 13725 7293 13737 7327
rect 13771 7293 13783 7327
rect 13725 7287 13783 7293
rect 13909 7327 13967 7333
rect 13909 7293 13921 7327
rect 13955 7293 13967 7327
rect 13909 7287 13967 7293
rect 11756 7228 13032 7256
rect 11756 7216 11762 7228
rect 9401 7191 9459 7197
rect 9401 7188 9413 7191
rect 9180 7160 9413 7188
rect 9180 7148 9186 7160
rect 9401 7157 9413 7160
rect 9447 7157 9459 7191
rect 9401 7151 9459 7157
rect 10413 7191 10471 7197
rect 10413 7157 10425 7191
rect 10459 7157 10471 7191
rect 10413 7151 10471 7157
rect 11517 7191 11575 7197
rect 11517 7157 11529 7191
rect 11563 7188 11575 7191
rect 11790 7188 11796 7200
rect 11563 7160 11796 7188
rect 11563 7157 11575 7160
rect 11517 7151 11575 7157
rect 11790 7148 11796 7160
rect 11848 7148 11854 7200
rect 11882 7148 11888 7200
rect 11940 7188 11946 7200
rect 13740 7188 13768 7287
rect 13924 7256 13952 7287
rect 14182 7284 14188 7336
rect 14240 7324 14246 7336
rect 14568 7333 14596 7364
rect 17037 7361 17049 7395
rect 17083 7392 17095 7395
rect 17678 7392 17684 7404
rect 17083 7364 17684 7392
rect 17083 7361 17095 7364
rect 17037 7355 17095 7361
rect 17678 7352 17684 7364
rect 17736 7352 17742 7404
rect 19444 7401 19472 7432
rect 20162 7420 20168 7472
rect 20220 7420 20226 7472
rect 21468 7460 21496 7488
rect 21726 7460 21732 7472
rect 21468 7432 21732 7460
rect 21726 7420 21732 7432
rect 21784 7420 21790 7472
rect 21821 7463 21879 7469
rect 21821 7429 21833 7463
rect 21867 7460 21879 7463
rect 22189 7463 22247 7469
rect 22189 7460 22201 7463
rect 21867 7432 22201 7460
rect 21867 7429 21879 7432
rect 21821 7423 21879 7429
rect 22189 7429 22201 7432
rect 22235 7429 22247 7463
rect 22189 7423 22247 7429
rect 19429 7395 19487 7401
rect 17788 7364 19380 7392
rect 14369 7327 14427 7333
rect 14369 7324 14381 7327
rect 14240 7296 14381 7324
rect 14240 7284 14246 7296
rect 14369 7293 14381 7296
rect 14415 7293 14427 7327
rect 14369 7287 14427 7293
rect 14553 7327 14611 7333
rect 14553 7293 14565 7327
rect 14599 7293 14611 7327
rect 14553 7287 14611 7293
rect 14737 7327 14795 7333
rect 14737 7293 14749 7327
rect 14783 7324 14795 7327
rect 14918 7324 14924 7336
rect 14783 7296 14924 7324
rect 14783 7293 14795 7296
rect 14737 7287 14795 7293
rect 14918 7284 14924 7296
rect 14976 7284 14982 7336
rect 15470 7284 15476 7336
rect 15528 7284 15534 7336
rect 16666 7284 16672 7336
rect 16724 7324 16730 7336
rect 16761 7327 16819 7333
rect 16761 7324 16773 7327
rect 16724 7296 16773 7324
rect 16724 7284 16730 7296
rect 16761 7293 16773 7296
rect 16807 7293 16819 7327
rect 16761 7287 16819 7293
rect 14461 7259 14519 7265
rect 14461 7256 14473 7259
rect 13924 7228 14473 7256
rect 14461 7225 14473 7228
rect 14507 7225 14519 7259
rect 17788 7256 17816 7364
rect 19352 7333 19380 7364
rect 19429 7361 19441 7395
rect 19475 7361 19487 7395
rect 19429 7355 19487 7361
rect 19981 7395 20039 7401
rect 19981 7361 19993 7395
rect 20027 7392 20039 7395
rect 20070 7392 20076 7404
rect 20027 7364 20076 7392
rect 20027 7361 20039 7364
rect 19981 7355 20039 7361
rect 18417 7327 18475 7333
rect 18417 7293 18429 7327
rect 18463 7293 18475 7327
rect 18417 7287 18475 7293
rect 19337 7327 19395 7333
rect 19337 7293 19349 7327
rect 19383 7293 19395 7327
rect 19337 7287 19395 7293
rect 14461 7219 14519 7225
rect 15856 7228 17816 7256
rect 18432 7256 18460 7287
rect 19610 7284 19616 7336
rect 19668 7284 19674 7336
rect 19705 7327 19763 7333
rect 19705 7293 19717 7327
rect 19751 7324 19763 7327
rect 19996 7324 20024 7355
rect 20070 7352 20076 7364
rect 20128 7352 20134 7404
rect 20180 7392 20208 7420
rect 20257 7395 20315 7401
rect 20257 7392 20269 7395
rect 20180 7364 20269 7392
rect 20257 7361 20269 7364
rect 20303 7361 20315 7395
rect 20257 7355 20315 7361
rect 22278 7352 22284 7404
rect 22336 7352 22342 7404
rect 21818 7324 21824 7336
rect 19751 7296 20024 7324
rect 20180 7296 21824 7324
rect 19751 7293 19763 7296
rect 19705 7287 19763 7293
rect 19720 7256 19748 7287
rect 18432 7228 19748 7256
rect 11940 7160 13768 7188
rect 11940 7148 11946 7160
rect 14090 7148 14096 7200
rect 14148 7148 14154 7200
rect 14182 7148 14188 7200
rect 14240 7148 14246 7200
rect 14476 7188 14504 7219
rect 14642 7188 14648 7200
rect 14476 7160 14648 7188
rect 14642 7148 14648 7160
rect 14700 7148 14706 7200
rect 15010 7148 15016 7200
rect 15068 7188 15074 7200
rect 15657 7191 15715 7197
rect 15657 7188 15669 7191
rect 15068 7160 15669 7188
rect 15068 7148 15074 7160
rect 15657 7157 15669 7160
rect 15703 7188 15715 7191
rect 15856 7188 15884 7228
rect 19794 7216 19800 7268
rect 19852 7256 19858 7268
rect 20180 7256 20208 7296
rect 21818 7284 21824 7296
rect 21876 7284 21882 7336
rect 21910 7284 21916 7336
rect 21968 7284 21974 7336
rect 19852 7228 20208 7256
rect 19852 7216 19858 7228
rect 21450 7216 21456 7268
rect 21508 7216 21514 7268
rect 21634 7216 21640 7268
rect 21692 7265 21698 7268
rect 21692 7259 21711 7265
rect 21699 7225 21711 7259
rect 21692 7219 21711 7225
rect 21692 7216 21698 7219
rect 22094 7216 22100 7268
rect 22152 7256 22158 7268
rect 22373 7259 22431 7265
rect 22373 7256 22385 7259
rect 22152 7228 22385 7256
rect 22152 7216 22158 7228
rect 22373 7225 22385 7228
rect 22419 7225 22431 7259
rect 22373 7219 22431 7225
rect 15703 7160 15884 7188
rect 15703 7157 15715 7160
rect 15657 7151 15715 7157
rect 16850 7148 16856 7200
rect 16908 7188 16914 7200
rect 17037 7191 17095 7197
rect 17037 7188 17049 7191
rect 16908 7160 17049 7188
rect 16908 7148 16914 7160
rect 17037 7157 17049 7160
rect 17083 7157 17095 7191
rect 17037 7151 17095 7157
rect 19889 7191 19947 7197
rect 19889 7157 19901 7191
rect 19935 7188 19947 7191
rect 20162 7188 20168 7200
rect 19935 7160 20168 7188
rect 19935 7157 19947 7160
rect 19889 7151 19947 7157
rect 20162 7148 20168 7160
rect 20220 7148 20226 7200
rect 21542 7148 21548 7200
rect 21600 7188 21606 7200
rect 22005 7191 22063 7197
rect 22005 7188 22017 7191
rect 21600 7160 22017 7188
rect 21600 7148 21606 7160
rect 22005 7157 22017 7160
rect 22051 7157 22063 7191
rect 22005 7151 22063 7157
rect 552 7098 23368 7120
rect 552 7046 4366 7098
rect 4418 7046 4430 7098
rect 4482 7046 4494 7098
rect 4546 7046 4558 7098
rect 4610 7046 4622 7098
rect 4674 7046 4686 7098
rect 4738 7046 10366 7098
rect 10418 7046 10430 7098
rect 10482 7046 10494 7098
rect 10546 7046 10558 7098
rect 10610 7046 10622 7098
rect 10674 7046 10686 7098
rect 10738 7046 16366 7098
rect 16418 7046 16430 7098
rect 16482 7046 16494 7098
rect 16546 7046 16558 7098
rect 16610 7046 16622 7098
rect 16674 7046 16686 7098
rect 16738 7046 22366 7098
rect 22418 7046 22430 7098
rect 22482 7046 22494 7098
rect 22546 7046 22558 7098
rect 22610 7046 22622 7098
rect 22674 7046 22686 7098
rect 22738 7046 23368 7098
rect 552 7024 23368 7046
rect 1486 6944 1492 6996
rect 1544 6984 1550 6996
rect 1673 6987 1731 6993
rect 1673 6984 1685 6987
rect 1544 6956 1685 6984
rect 1544 6944 1550 6956
rect 1673 6953 1685 6956
rect 1719 6953 1731 6987
rect 1673 6947 1731 6953
rect 1688 6916 1716 6947
rect 1762 6944 1768 6996
rect 1820 6984 1826 6996
rect 1820 6956 2360 6984
rect 1820 6944 1826 6956
rect 1688 6888 1992 6916
rect 1213 6851 1271 6857
rect 1213 6817 1225 6851
rect 1259 6817 1271 6851
rect 1213 6811 1271 6817
rect 1673 6851 1731 6857
rect 1673 6817 1685 6851
rect 1719 6848 1731 6851
rect 1762 6848 1768 6860
rect 1719 6820 1768 6848
rect 1719 6817 1731 6820
rect 1673 6811 1731 6817
rect 1118 6740 1124 6792
rect 1176 6740 1182 6792
rect 1228 6780 1256 6811
rect 1762 6808 1768 6820
rect 1820 6808 1826 6860
rect 1854 6808 1860 6860
rect 1912 6808 1918 6860
rect 1964 6857 1992 6888
rect 1949 6851 2007 6857
rect 1949 6817 1961 6851
rect 1995 6817 2007 6851
rect 1949 6811 2007 6817
rect 2130 6808 2136 6860
rect 2188 6808 2194 6860
rect 2332 6857 2360 6956
rect 4062 6944 4068 6996
rect 4120 6984 4126 6996
rect 4430 6984 4436 6996
rect 4120 6956 4436 6984
rect 4120 6944 4126 6956
rect 4430 6944 4436 6956
rect 4488 6984 4494 6996
rect 5810 6984 5816 6996
rect 4488 6956 5816 6984
rect 4488 6944 4494 6956
rect 5810 6944 5816 6956
rect 5868 6984 5874 6996
rect 5994 6984 6000 6996
rect 5868 6956 6000 6984
rect 5868 6944 5874 6956
rect 5994 6944 6000 6956
rect 6052 6944 6058 6996
rect 6270 6944 6276 6996
rect 6328 6944 6334 6996
rect 7742 6944 7748 6996
rect 7800 6984 7806 6996
rect 9125 6987 9183 6993
rect 7800 6956 8984 6984
rect 7800 6944 7806 6956
rect 2958 6916 2964 6928
rect 2608 6888 2964 6916
rect 2317 6851 2375 6857
rect 2317 6817 2329 6851
rect 2363 6817 2375 6851
rect 2498 6848 2504 6860
rect 2459 6820 2504 6848
rect 2317 6811 2375 6817
rect 2498 6808 2504 6820
rect 2556 6848 2562 6860
rect 2608 6848 2636 6888
rect 2958 6876 2964 6888
rect 3016 6876 3022 6928
rect 4890 6916 4896 6928
rect 4172 6888 4896 6916
rect 2556 6820 2636 6848
rect 2556 6808 2562 6820
rect 2682 6808 2688 6860
rect 2740 6848 2746 6860
rect 2777 6851 2835 6857
rect 2777 6848 2789 6851
rect 2740 6820 2789 6848
rect 2740 6808 2746 6820
rect 2777 6817 2789 6820
rect 2823 6817 2835 6851
rect 2777 6811 2835 6817
rect 3510 6808 3516 6860
rect 3568 6808 3574 6860
rect 3694 6808 3700 6860
rect 3752 6808 3758 6860
rect 4172 6857 4200 6888
rect 4157 6851 4215 6857
rect 4157 6817 4169 6851
rect 4203 6817 4215 6851
rect 4157 6811 4215 6817
rect 4246 6808 4252 6860
rect 4304 6808 4310 6860
rect 2041 6783 2099 6789
rect 2041 6780 2053 6783
rect 1228 6752 2053 6780
rect 2041 6749 2053 6752
rect 2087 6749 2099 6783
rect 2041 6743 2099 6749
rect 2869 6783 2927 6789
rect 2869 6749 2881 6783
rect 2915 6780 2927 6783
rect 3050 6780 3056 6792
rect 2915 6752 3056 6780
rect 2915 6749 2927 6752
rect 2869 6743 2927 6749
rect 3050 6740 3056 6752
rect 3108 6740 3114 6792
rect 4264 6780 4292 6808
rect 3160 6752 4292 6780
rect 1581 6715 1639 6721
rect 1581 6681 1593 6715
rect 1627 6712 1639 6715
rect 2501 6715 2559 6721
rect 1627 6684 2176 6712
rect 1627 6681 1639 6684
rect 1581 6675 1639 6681
rect 2148 6644 2176 6684
rect 2501 6681 2513 6715
rect 2547 6712 2559 6715
rect 2774 6712 2780 6724
rect 2547 6684 2780 6712
rect 2547 6681 2559 6684
rect 2501 6675 2559 6681
rect 2774 6672 2780 6684
rect 2832 6672 2838 6724
rect 3160 6721 3188 6752
rect 3145 6715 3203 6721
rect 3145 6681 3157 6715
rect 3191 6681 3203 6715
rect 4356 6712 4384 6888
rect 4890 6876 4896 6888
rect 4948 6876 4954 6928
rect 5077 6919 5135 6925
rect 5077 6885 5089 6919
rect 5123 6916 5135 6919
rect 7466 6916 7472 6928
rect 5123 6888 7472 6916
rect 5123 6885 5135 6888
rect 5077 6879 5135 6885
rect 7466 6876 7472 6888
rect 7524 6876 7530 6928
rect 8846 6916 8852 6928
rect 8312 6888 8852 6916
rect 4430 6808 4436 6860
rect 4488 6808 4494 6860
rect 4798 6808 4804 6860
rect 4856 6808 4862 6860
rect 5353 6851 5411 6857
rect 5353 6817 5365 6851
rect 5399 6848 5411 6851
rect 5399 6820 5488 6848
rect 5399 6817 5411 6820
rect 5353 6811 5411 6817
rect 5077 6783 5135 6789
rect 5077 6749 5089 6783
rect 5123 6780 5135 6783
rect 5460 6780 5488 6820
rect 5534 6808 5540 6860
rect 5592 6808 5598 6860
rect 5629 6851 5687 6857
rect 5629 6817 5641 6851
rect 5675 6848 5687 6851
rect 6178 6848 6184 6860
rect 5675 6820 6184 6848
rect 5675 6817 5687 6820
rect 5629 6811 5687 6817
rect 6178 6808 6184 6820
rect 6236 6808 6242 6860
rect 6332 6851 6390 6857
rect 6332 6817 6344 6851
rect 6378 6848 6390 6851
rect 7190 6848 7196 6860
rect 6378 6820 7196 6848
rect 6378 6817 6390 6820
rect 6332 6811 6390 6817
rect 7190 6808 7196 6820
rect 7248 6808 7254 6860
rect 8110 6848 8116 6860
rect 7300 6820 8116 6848
rect 5123 6752 5488 6780
rect 5123 6749 5135 6752
rect 5077 6743 5135 6749
rect 3145 6675 3203 6681
rect 3804 6684 4384 6712
rect 5460 6712 5488 6752
rect 5813 6783 5871 6789
rect 5813 6749 5825 6783
rect 5859 6780 5871 6783
rect 6914 6780 6920 6792
rect 5859 6752 6920 6780
rect 5859 6749 5871 6752
rect 5813 6743 5871 6749
rect 6914 6740 6920 6752
rect 6972 6740 6978 6792
rect 7101 6783 7159 6789
rect 7101 6749 7113 6783
rect 7147 6780 7159 6783
rect 7300 6780 7328 6820
rect 8110 6808 8116 6820
rect 8168 6808 8174 6860
rect 8312 6857 8340 6888
rect 8846 6876 8852 6888
rect 8904 6876 8910 6928
rect 8956 6916 8984 6956
rect 9125 6953 9137 6987
rect 9171 6984 9183 6987
rect 9858 6984 9864 6996
rect 9171 6956 9864 6984
rect 9171 6953 9183 6956
rect 9125 6947 9183 6953
rect 9858 6944 9864 6956
rect 9916 6944 9922 6996
rect 10226 6944 10232 6996
rect 10284 6984 10290 6996
rect 11606 6984 11612 6996
rect 10284 6956 11612 6984
rect 10284 6944 10290 6956
rect 11606 6944 11612 6956
rect 11664 6944 11670 6996
rect 11698 6944 11704 6996
rect 11756 6984 11762 6996
rect 11756 6956 12020 6984
rect 11756 6944 11762 6956
rect 11882 6916 11888 6928
rect 8956 6888 11888 6916
rect 11882 6876 11888 6888
rect 11940 6876 11946 6928
rect 8297 6851 8355 6857
rect 8297 6817 8309 6851
rect 8343 6817 8355 6851
rect 8297 6811 8355 6817
rect 8389 6851 8447 6857
rect 8389 6817 8401 6851
rect 8435 6848 8447 6851
rect 9030 6848 9036 6860
rect 8435 6820 9036 6848
rect 8435 6817 8447 6820
rect 8389 6811 8447 6817
rect 7147 6752 7328 6780
rect 7377 6783 7435 6789
rect 7147 6749 7159 6752
rect 7101 6743 7159 6749
rect 7377 6749 7389 6783
rect 7423 6780 7435 6783
rect 8312 6780 8340 6811
rect 9030 6808 9036 6820
rect 9088 6808 9094 6860
rect 9184 6851 9242 6857
rect 9184 6817 9196 6851
rect 9230 6848 9242 6851
rect 9306 6848 9312 6860
rect 9230 6820 9312 6848
rect 9230 6817 9242 6820
rect 9184 6811 9242 6817
rect 9306 6808 9312 6820
rect 9364 6808 9370 6860
rect 9582 6808 9588 6860
rect 9640 6808 9646 6860
rect 9766 6808 9772 6860
rect 9824 6808 9830 6860
rect 9861 6851 9919 6857
rect 9861 6817 9873 6851
rect 9907 6848 9919 6851
rect 10137 6851 10195 6857
rect 9907 6820 10106 6848
rect 9907 6817 9919 6820
rect 9861 6811 9919 6817
rect 7423 6752 8340 6780
rect 8665 6783 8723 6789
rect 7423 6749 7435 6752
rect 7377 6743 7435 6749
rect 8665 6749 8677 6783
rect 8711 6749 8723 6783
rect 8665 6743 8723 6749
rect 6362 6712 6368 6724
rect 5460 6684 6368 6712
rect 3804 6644 3832 6684
rect 6362 6672 6368 6684
rect 6420 6672 6426 6724
rect 6454 6672 6460 6724
rect 6512 6672 6518 6724
rect 6546 6672 6552 6724
rect 6604 6712 6610 6724
rect 8680 6712 8708 6743
rect 8754 6740 8760 6792
rect 8812 6740 8818 6792
rect 9876 6712 9904 6811
rect 9953 6783 10011 6789
rect 9953 6749 9965 6783
rect 9999 6749 10011 6783
rect 10078 6780 10106 6820
rect 10137 6817 10149 6851
rect 10183 6848 10195 6851
rect 10318 6848 10324 6860
rect 10183 6820 10324 6848
rect 10183 6817 10195 6820
rect 10137 6811 10195 6817
rect 10318 6808 10324 6820
rect 10376 6808 10382 6860
rect 10410 6808 10416 6860
rect 10468 6808 10474 6860
rect 10597 6851 10655 6857
rect 10597 6817 10609 6851
rect 10643 6848 10655 6851
rect 10686 6848 10692 6860
rect 10643 6820 10692 6848
rect 10643 6817 10655 6820
rect 10597 6811 10655 6817
rect 10686 6808 10692 6820
rect 10744 6808 10750 6860
rect 10781 6851 10839 6857
rect 10781 6817 10793 6851
rect 10827 6848 10839 6851
rect 10965 6851 11023 6857
rect 10965 6848 10977 6851
rect 10827 6820 10977 6848
rect 10827 6817 10839 6820
rect 10781 6811 10839 6817
rect 10965 6817 10977 6820
rect 11011 6817 11023 6851
rect 10965 6811 11023 6817
rect 11146 6808 11152 6860
rect 11204 6808 11210 6860
rect 11238 6808 11244 6860
rect 11296 6808 11302 6860
rect 11517 6851 11575 6857
rect 11517 6817 11529 6851
rect 11563 6817 11575 6851
rect 11517 6811 11575 6817
rect 10502 6780 10508 6792
rect 10078 6752 10508 6780
rect 9953 6743 10011 6749
rect 6604 6684 8708 6712
rect 9232 6684 9904 6712
rect 9968 6712 9996 6743
rect 10502 6740 10508 6752
rect 10560 6740 10566 6792
rect 11333 6783 11391 6789
rect 11333 6749 11345 6783
rect 11379 6780 11391 6783
rect 11422 6780 11428 6792
rect 11379 6752 11428 6780
rect 11379 6749 11391 6752
rect 11333 6743 11391 6749
rect 11422 6740 11428 6752
rect 11480 6740 11486 6792
rect 11532 6780 11560 6811
rect 11606 6808 11612 6860
rect 11664 6848 11670 6860
rect 11992 6857 12020 6956
rect 12526 6944 12532 6996
rect 12584 6984 12590 6996
rect 13078 6984 13084 6996
rect 12584 6956 13084 6984
rect 12584 6944 12590 6956
rect 13078 6944 13084 6956
rect 13136 6984 13142 6996
rect 13449 6987 13507 6993
rect 13449 6984 13461 6987
rect 13136 6956 13461 6984
rect 13136 6944 13142 6956
rect 13449 6953 13461 6956
rect 13495 6953 13507 6987
rect 13449 6947 13507 6953
rect 14734 6944 14740 6996
rect 14792 6984 14798 6996
rect 16577 6987 16635 6993
rect 16577 6984 16589 6987
rect 14792 6956 16589 6984
rect 14792 6944 14798 6956
rect 16577 6953 16589 6956
rect 16623 6953 16635 6987
rect 16577 6947 16635 6953
rect 17218 6944 17224 6996
rect 17276 6984 17282 6996
rect 19794 6984 19800 6996
rect 17276 6956 19800 6984
rect 17276 6944 17282 6956
rect 19794 6944 19800 6956
rect 19852 6944 19858 6996
rect 20254 6944 20260 6996
rect 20312 6984 20318 6996
rect 21542 6984 21548 6996
rect 20312 6956 21548 6984
rect 20312 6944 20318 6956
rect 21542 6944 21548 6956
rect 21600 6944 21606 6996
rect 15654 6916 15660 6928
rect 12636 6888 15660 6916
rect 12636 6857 12664 6888
rect 15654 6876 15660 6888
rect 15712 6876 15718 6928
rect 11793 6851 11851 6857
rect 11793 6848 11805 6851
rect 11664 6820 11805 6848
rect 11664 6808 11670 6820
rect 11793 6817 11805 6820
rect 11839 6817 11851 6851
rect 11793 6811 11851 6817
rect 11977 6851 12035 6857
rect 11977 6817 11989 6851
rect 12023 6817 12035 6851
rect 11977 6811 12035 6817
rect 12161 6851 12219 6857
rect 12161 6817 12173 6851
rect 12207 6848 12219 6851
rect 12437 6851 12495 6857
rect 12437 6848 12449 6851
rect 12207 6820 12449 6848
rect 12207 6817 12219 6820
rect 12161 6811 12219 6817
rect 12437 6817 12449 6820
rect 12483 6817 12495 6851
rect 12437 6811 12495 6817
rect 12621 6851 12679 6857
rect 12621 6817 12633 6851
rect 12667 6817 12679 6851
rect 12621 6811 12679 6817
rect 12989 6851 13047 6857
rect 12989 6817 13001 6851
rect 13035 6817 13047 6851
rect 12989 6811 13047 6817
rect 11698 6780 11704 6792
rect 11532 6752 11704 6780
rect 11698 6740 11704 6752
rect 11756 6780 11762 6792
rect 12713 6783 12771 6789
rect 12713 6780 12725 6783
rect 11756 6752 12725 6780
rect 11756 6740 11762 6752
rect 12713 6749 12725 6752
rect 12759 6749 12771 6783
rect 12713 6743 12771 6749
rect 12802 6740 12808 6792
rect 12860 6740 12866 6792
rect 11440 6712 11468 6740
rect 9968 6684 11468 6712
rect 6604 6672 6610 6684
rect 2148 6616 3832 6644
rect 3881 6647 3939 6653
rect 3881 6613 3893 6647
rect 3927 6644 3939 6647
rect 4522 6644 4528 6656
rect 3927 6616 4528 6644
rect 3927 6613 3939 6616
rect 3881 6607 3939 6613
rect 4522 6604 4528 6616
rect 4580 6604 4586 6656
rect 4617 6647 4675 6653
rect 4617 6613 4629 6647
rect 4663 6644 4675 6647
rect 4893 6647 4951 6653
rect 4893 6644 4905 6647
rect 4663 6616 4905 6644
rect 4663 6613 4675 6616
rect 4617 6607 4675 6613
rect 4893 6613 4905 6616
rect 4939 6613 4951 6647
rect 4893 6607 4951 6613
rect 5169 6647 5227 6653
rect 5169 6613 5181 6647
rect 5215 6644 5227 6647
rect 5442 6644 5448 6656
rect 5215 6616 5448 6644
rect 5215 6613 5227 6616
rect 5169 6607 5227 6613
rect 5442 6604 5448 6616
rect 5500 6604 5506 6656
rect 5902 6604 5908 6656
rect 5960 6604 5966 6656
rect 7190 6604 7196 6656
rect 7248 6644 7254 6656
rect 7742 6644 7748 6656
rect 7248 6616 7748 6644
rect 7248 6604 7254 6616
rect 7742 6604 7748 6616
rect 7800 6604 7806 6656
rect 8067 6647 8125 6653
rect 8067 6613 8079 6647
rect 8113 6644 8125 6647
rect 8386 6644 8392 6656
rect 8113 6616 8392 6644
rect 8113 6613 8125 6616
rect 8067 6607 8125 6613
rect 8386 6604 8392 6616
rect 8444 6604 8450 6656
rect 8573 6647 8631 6653
rect 8573 6613 8585 6647
rect 8619 6644 8631 6647
rect 8662 6644 8668 6656
rect 8619 6616 8668 6644
rect 8619 6613 8631 6616
rect 8573 6607 8631 6613
rect 8662 6604 8668 6616
rect 8720 6644 8726 6656
rect 9232 6644 9260 6684
rect 11514 6672 11520 6724
rect 11572 6712 11578 6724
rect 13004 6712 13032 6811
rect 13078 6808 13084 6860
rect 13136 6848 13142 6860
rect 13390 6851 13448 6857
rect 13390 6848 13402 6851
rect 13136 6820 13402 6848
rect 13136 6808 13142 6820
rect 13390 6817 13402 6820
rect 13436 6817 13448 6851
rect 13390 6811 13448 6817
rect 13817 6851 13875 6857
rect 13817 6817 13829 6851
rect 13863 6848 13875 6851
rect 14090 6848 14096 6860
rect 13863 6820 14096 6848
rect 13863 6817 13875 6820
rect 13817 6811 13875 6817
rect 14090 6808 14096 6820
rect 14148 6808 14154 6860
rect 14182 6808 14188 6860
rect 14240 6808 14246 6860
rect 14366 6808 14372 6860
rect 14424 6808 14430 6860
rect 14458 6808 14464 6860
rect 14516 6808 14522 6860
rect 14642 6808 14648 6860
rect 14700 6808 14706 6860
rect 14936 6820 15148 6848
rect 13906 6740 13912 6792
rect 13964 6740 13970 6792
rect 14476 6780 14504 6808
rect 14936 6789 14964 6820
rect 14737 6783 14795 6789
rect 14737 6780 14749 6783
rect 14476 6752 14749 6780
rect 14737 6749 14749 6752
rect 14783 6749 14795 6783
rect 14737 6743 14795 6749
rect 14921 6783 14979 6789
rect 14921 6749 14933 6783
rect 14967 6749 14979 6783
rect 14921 6743 14979 6749
rect 15010 6740 15016 6792
rect 15068 6740 15074 6792
rect 15120 6780 15148 6820
rect 15194 6808 15200 6860
rect 15252 6808 15258 6860
rect 15286 6808 15292 6860
rect 15344 6808 15350 6860
rect 15378 6808 15384 6860
rect 15436 6808 15442 6860
rect 15470 6808 15476 6860
rect 15528 6848 15534 6860
rect 16485 6851 16543 6857
rect 16485 6848 16497 6851
rect 15528 6820 16497 6848
rect 15528 6808 15534 6820
rect 16485 6817 16497 6820
rect 16531 6848 16543 6851
rect 17034 6848 17040 6860
rect 16531 6820 17040 6848
rect 16531 6817 16543 6820
rect 16485 6811 16543 6817
rect 17034 6808 17040 6820
rect 17092 6808 17098 6860
rect 17310 6808 17316 6860
rect 17368 6808 17374 6860
rect 17402 6808 17408 6860
rect 17460 6808 17466 6860
rect 17494 6808 17500 6860
rect 17552 6808 17558 6860
rect 18230 6808 18236 6860
rect 18288 6808 18294 6860
rect 18322 6808 18328 6860
rect 18380 6808 18386 6860
rect 19702 6848 19708 6860
rect 18432 6820 19708 6848
rect 15120 6752 16528 6780
rect 16500 6724 16528 6752
rect 16758 6740 16764 6792
rect 16816 6740 16822 6792
rect 17221 6783 17279 6789
rect 17221 6749 17233 6783
rect 17267 6749 17279 6783
rect 17221 6743 17279 6749
rect 17681 6783 17739 6789
rect 17681 6749 17693 6783
rect 17727 6780 17739 6783
rect 18432 6780 18460 6820
rect 19702 6808 19708 6820
rect 19760 6808 19766 6860
rect 19812 6848 19840 6944
rect 19886 6876 19892 6928
rect 19944 6916 19950 6928
rect 19944 6888 20668 6916
rect 19944 6876 19950 6888
rect 20027 6851 20085 6857
rect 20027 6848 20039 6851
rect 19812 6820 20039 6848
rect 20027 6817 20039 6820
rect 20073 6817 20085 6851
rect 20027 6811 20085 6817
rect 20254 6808 20260 6860
rect 20312 6848 20318 6860
rect 20441 6851 20499 6857
rect 20312 6820 20392 6848
rect 20312 6808 20318 6820
rect 17727 6752 18460 6780
rect 17727 6749 17739 6752
rect 17681 6743 17739 6749
rect 13265 6715 13323 6721
rect 13265 6712 13277 6715
rect 11572 6684 13032 6712
rect 13096 6684 13277 6712
rect 11572 6672 11578 6684
rect 8720 6616 9260 6644
rect 9309 6647 9367 6653
rect 8720 6604 8726 6616
rect 9309 6613 9321 6647
rect 9355 6644 9367 6647
rect 9490 6644 9496 6656
rect 9355 6616 9496 6644
rect 9355 6613 9367 6616
rect 9309 6607 9367 6613
rect 9490 6604 9496 6616
rect 9548 6604 9554 6656
rect 10226 6604 10232 6656
rect 10284 6644 10290 6656
rect 10321 6647 10379 6653
rect 10321 6644 10333 6647
rect 10284 6616 10333 6644
rect 10284 6604 10290 6616
rect 10321 6613 10333 6616
rect 10367 6613 10379 6647
rect 10321 6607 10379 6613
rect 11146 6604 11152 6656
rect 11204 6644 11210 6656
rect 11701 6647 11759 6653
rect 11701 6644 11713 6647
rect 11204 6616 11713 6644
rect 11204 6604 11210 6616
rect 11701 6613 11713 6616
rect 11747 6613 11759 6647
rect 11701 6607 11759 6613
rect 12802 6604 12808 6656
rect 12860 6644 12866 6656
rect 13096 6644 13124 6684
rect 13265 6681 13277 6684
rect 13311 6681 13323 6715
rect 14829 6715 14887 6721
rect 14829 6712 14841 6715
rect 13265 6675 13323 6681
rect 14384 6684 14841 6712
rect 12860 6616 13124 6644
rect 13173 6647 13231 6653
rect 12860 6604 12866 6616
rect 13173 6613 13185 6647
rect 13219 6644 13231 6647
rect 14090 6644 14096 6656
rect 13219 6616 14096 6644
rect 13219 6613 13231 6616
rect 13173 6607 13231 6613
rect 14090 6604 14096 6616
rect 14148 6604 14154 6656
rect 14384 6653 14412 6684
rect 14829 6681 14841 6684
rect 14875 6681 14887 6715
rect 14829 6675 14887 6681
rect 15105 6715 15163 6721
rect 15105 6681 15117 6715
rect 15151 6712 15163 6715
rect 15286 6712 15292 6724
rect 15151 6684 15292 6712
rect 15151 6681 15163 6684
rect 15105 6675 15163 6681
rect 15286 6672 15292 6684
rect 15344 6672 15350 6724
rect 15396 6684 16252 6712
rect 14369 6647 14427 6653
rect 14369 6613 14381 6647
rect 14415 6613 14427 6647
rect 14369 6607 14427 6613
rect 14550 6604 14556 6656
rect 14608 6604 14614 6656
rect 14918 6604 14924 6656
rect 14976 6644 14982 6656
rect 15396 6644 15424 6684
rect 14976 6616 15424 6644
rect 14976 6604 14982 6616
rect 15470 6604 15476 6656
rect 15528 6644 15534 6656
rect 15565 6647 15623 6653
rect 15565 6644 15577 6647
rect 15528 6616 15577 6644
rect 15528 6604 15534 6616
rect 15565 6613 15577 6616
rect 15611 6613 15623 6647
rect 15565 6607 15623 6613
rect 15746 6604 15752 6656
rect 15804 6644 15810 6656
rect 16117 6647 16175 6653
rect 16117 6644 16129 6647
rect 15804 6616 16129 6644
rect 15804 6604 15810 6616
rect 16117 6613 16129 6616
rect 16163 6613 16175 6647
rect 16224 6644 16252 6684
rect 16482 6672 16488 6724
rect 16540 6672 16546 6724
rect 17236 6712 17264 6743
rect 18506 6740 18512 6792
rect 18564 6740 18570 6792
rect 18966 6740 18972 6792
rect 19024 6780 19030 6792
rect 19794 6780 19800 6792
rect 19024 6752 19800 6780
rect 19024 6740 19030 6752
rect 19794 6740 19800 6752
rect 19852 6740 19858 6792
rect 20162 6740 20168 6792
rect 20220 6740 20226 6792
rect 20364 6789 20392 6820
rect 20441 6817 20453 6851
rect 20487 6848 20499 6851
rect 20530 6848 20536 6860
rect 20487 6820 20536 6848
rect 20487 6817 20499 6820
rect 20441 6811 20499 6817
rect 20530 6808 20536 6820
rect 20588 6808 20594 6860
rect 20640 6857 20668 6888
rect 20714 6876 20720 6928
rect 20772 6916 20778 6928
rect 20772 6888 21496 6916
rect 20772 6876 20778 6888
rect 21468 6857 21496 6888
rect 20625 6851 20683 6857
rect 20625 6817 20637 6851
rect 20671 6817 20683 6851
rect 20625 6811 20683 6817
rect 21453 6851 21511 6857
rect 21453 6817 21465 6851
rect 21499 6817 21511 6851
rect 21453 6811 21511 6817
rect 21545 6851 21603 6857
rect 21545 6817 21557 6851
rect 21591 6848 21603 6851
rect 21634 6848 21640 6860
rect 21591 6820 21640 6848
rect 21591 6817 21603 6820
rect 21545 6811 21603 6817
rect 21634 6808 21640 6820
rect 21692 6808 21698 6860
rect 21821 6851 21879 6857
rect 21821 6817 21833 6851
rect 21867 6848 21879 6851
rect 22002 6848 22008 6860
rect 21867 6820 22008 6848
rect 21867 6817 21879 6820
rect 21821 6811 21879 6817
rect 22002 6808 22008 6820
rect 22060 6808 22066 6860
rect 20349 6783 20407 6789
rect 20349 6749 20361 6783
rect 20395 6749 20407 6783
rect 20349 6743 20407 6749
rect 20809 6783 20867 6789
rect 20809 6749 20821 6783
rect 20855 6780 20867 6783
rect 21269 6783 21327 6789
rect 21269 6780 21281 6783
rect 20855 6752 21281 6780
rect 20855 6749 20867 6752
rect 20809 6743 20867 6749
rect 21269 6749 21281 6752
rect 21315 6749 21327 6783
rect 21269 6743 21327 6749
rect 21910 6712 21916 6724
rect 17236 6684 21916 6712
rect 21910 6672 21916 6684
rect 21968 6672 21974 6724
rect 18138 6644 18144 6656
rect 16224 6616 18144 6644
rect 16117 6607 16175 6613
rect 18138 6604 18144 6616
rect 18196 6604 18202 6656
rect 18414 6604 18420 6656
rect 18472 6604 18478 6656
rect 18506 6604 18512 6656
rect 18564 6644 18570 6656
rect 19886 6644 19892 6656
rect 18564 6616 19892 6644
rect 18564 6604 18570 6616
rect 19886 6604 19892 6616
rect 19944 6604 19950 6656
rect 20257 6647 20315 6653
rect 20257 6613 20269 6647
rect 20303 6644 20315 6647
rect 20530 6644 20536 6656
rect 20303 6616 20536 6644
rect 20303 6613 20315 6616
rect 20257 6607 20315 6613
rect 20530 6604 20536 6616
rect 20588 6604 20594 6656
rect 20717 6647 20775 6653
rect 20717 6613 20729 6647
rect 20763 6644 20775 6647
rect 21450 6644 21456 6656
rect 20763 6616 21456 6644
rect 20763 6613 20775 6616
rect 20717 6607 20775 6613
rect 21450 6604 21456 6616
rect 21508 6604 21514 6656
rect 21729 6647 21787 6653
rect 21729 6613 21741 6647
rect 21775 6644 21787 6647
rect 21818 6644 21824 6656
rect 21775 6616 21824 6644
rect 21775 6613 21787 6616
rect 21729 6607 21787 6613
rect 21818 6604 21824 6616
rect 21876 6604 21882 6656
rect 552 6554 23368 6576
rect 552 6502 1366 6554
rect 1418 6502 1430 6554
rect 1482 6502 1494 6554
rect 1546 6502 1558 6554
rect 1610 6502 1622 6554
rect 1674 6502 1686 6554
rect 1738 6502 7366 6554
rect 7418 6502 7430 6554
rect 7482 6502 7494 6554
rect 7546 6502 7558 6554
rect 7610 6502 7622 6554
rect 7674 6502 7686 6554
rect 7738 6502 13366 6554
rect 13418 6502 13430 6554
rect 13482 6502 13494 6554
rect 13546 6502 13558 6554
rect 13610 6502 13622 6554
rect 13674 6502 13686 6554
rect 13738 6502 19366 6554
rect 19418 6502 19430 6554
rect 19482 6502 19494 6554
rect 19546 6502 19558 6554
rect 19610 6502 19622 6554
rect 19674 6502 19686 6554
rect 19738 6502 23368 6554
rect 552 6480 23368 6502
rect 3694 6440 3700 6452
rect 2884 6412 3700 6440
rect 1762 6196 1768 6248
rect 1820 6236 1826 6248
rect 1857 6239 1915 6245
rect 1857 6236 1869 6239
rect 1820 6208 1869 6236
rect 1820 6196 1826 6208
rect 1857 6205 1869 6208
rect 1903 6205 1915 6239
rect 1857 6199 1915 6205
rect 2038 6196 2044 6248
rect 2096 6196 2102 6248
rect 2130 6196 2136 6248
rect 2188 6236 2194 6248
rect 2317 6239 2375 6245
rect 2317 6236 2329 6239
rect 2188 6208 2329 6236
rect 2188 6196 2194 6208
rect 2317 6205 2329 6208
rect 2363 6236 2375 6239
rect 2406 6236 2412 6248
rect 2363 6208 2412 6236
rect 2363 6205 2375 6208
rect 2317 6199 2375 6205
rect 2406 6196 2412 6208
rect 2464 6196 2470 6248
rect 2884 6245 2912 6412
rect 3694 6400 3700 6412
rect 3752 6400 3758 6452
rect 5629 6443 5687 6449
rect 5629 6409 5641 6443
rect 5675 6440 5687 6443
rect 5718 6440 5724 6452
rect 5675 6412 5724 6440
rect 5675 6409 5687 6412
rect 5629 6403 5687 6409
rect 5718 6400 5724 6412
rect 5776 6400 5782 6452
rect 5810 6400 5816 6452
rect 5868 6400 5874 6452
rect 5902 6400 5908 6452
rect 5960 6440 5966 6452
rect 6457 6443 6515 6449
rect 6457 6440 6469 6443
rect 5960 6412 6469 6440
rect 5960 6400 5966 6412
rect 6457 6409 6469 6412
rect 6503 6409 6515 6443
rect 6457 6403 6515 6409
rect 8846 6400 8852 6452
rect 8904 6440 8910 6452
rect 9214 6440 9220 6452
rect 8904 6412 9220 6440
rect 8904 6400 8910 6412
rect 9214 6400 9220 6412
rect 9272 6400 9278 6452
rect 9582 6400 9588 6452
rect 9640 6400 9646 6452
rect 10318 6400 10324 6452
rect 10376 6440 10382 6452
rect 10873 6443 10931 6449
rect 10873 6440 10885 6443
rect 10376 6412 10885 6440
rect 10376 6400 10382 6412
rect 10873 6409 10885 6412
rect 10919 6440 10931 6443
rect 11238 6440 11244 6452
rect 10919 6412 11244 6440
rect 10919 6409 10931 6412
rect 10873 6403 10931 6409
rect 11238 6400 11244 6412
rect 11296 6400 11302 6452
rect 12161 6443 12219 6449
rect 12161 6409 12173 6443
rect 12207 6440 12219 6443
rect 12434 6440 12440 6452
rect 12207 6412 12440 6440
rect 12207 6409 12219 6412
rect 12161 6403 12219 6409
rect 12434 6400 12440 6412
rect 12492 6400 12498 6452
rect 14093 6443 14151 6449
rect 14093 6409 14105 6443
rect 14139 6440 14151 6443
rect 14921 6443 14979 6449
rect 14139 6412 14872 6440
rect 14139 6409 14151 6412
rect 14093 6403 14151 6409
rect 5261 6375 5319 6381
rect 3620 6344 4292 6372
rect 2961 6307 3019 6313
rect 2961 6273 2973 6307
rect 3007 6304 3019 6307
rect 3620 6304 3648 6344
rect 3007 6276 3648 6304
rect 3007 6273 3019 6276
rect 2961 6267 3019 6273
rect 2869 6239 2927 6245
rect 2869 6205 2881 6239
rect 2915 6205 2927 6239
rect 2869 6199 2927 6205
rect 3053 6239 3111 6245
rect 3053 6205 3065 6239
rect 3099 6236 3111 6239
rect 3510 6236 3516 6248
rect 3099 6208 3516 6236
rect 3099 6205 3111 6208
rect 3053 6199 3111 6205
rect 3510 6196 3516 6208
rect 3568 6196 3574 6248
rect 3620 6245 3648 6276
rect 3789 6307 3847 6313
rect 3789 6273 3801 6307
rect 3835 6304 3847 6307
rect 4062 6304 4068 6316
rect 3835 6276 4068 6304
rect 3835 6273 3847 6276
rect 3789 6267 3847 6273
rect 4062 6264 4068 6276
rect 4120 6264 4126 6316
rect 3605 6239 3663 6245
rect 3605 6205 3617 6239
rect 3651 6205 3663 6239
rect 3605 6199 3663 6205
rect 3881 6239 3939 6245
rect 3881 6205 3893 6239
rect 3927 6236 3939 6239
rect 4157 6239 4215 6245
rect 4157 6236 4169 6239
rect 3927 6208 4169 6236
rect 3927 6205 3939 6208
rect 3881 6199 3939 6205
rect 4157 6205 4169 6208
rect 4203 6205 4215 6239
rect 4264 6236 4292 6344
rect 5261 6341 5273 6375
rect 5307 6372 5319 6375
rect 7561 6375 7619 6381
rect 5307 6344 7512 6372
rect 5307 6341 5319 6344
rect 5261 6335 5319 6341
rect 4522 6264 4528 6316
rect 4580 6304 4586 6316
rect 5721 6307 5779 6313
rect 4580 6276 4844 6304
rect 4580 6264 4586 6276
rect 4816 6245 4844 6276
rect 5721 6273 5733 6307
rect 5767 6304 5779 6307
rect 6181 6307 6239 6313
rect 6181 6304 6193 6307
rect 5767 6276 6193 6304
rect 5767 6273 5779 6276
rect 5721 6267 5779 6273
rect 6181 6273 6193 6276
rect 6227 6273 6239 6307
rect 6181 6267 6239 6273
rect 7285 6307 7343 6313
rect 7285 6273 7297 6307
rect 7331 6273 7343 6307
rect 7484 6304 7512 6344
rect 7561 6341 7573 6375
rect 7607 6372 7619 6375
rect 7834 6372 7840 6384
rect 7607 6344 7840 6372
rect 7607 6341 7619 6344
rect 7561 6335 7619 6341
rect 7834 6332 7840 6344
rect 7892 6332 7898 6384
rect 8294 6332 8300 6384
rect 8352 6372 8358 6384
rect 8352 6344 11284 6372
rect 8352 6332 8358 6344
rect 7484 6276 8984 6304
rect 7285 6267 7343 6273
rect 4617 6239 4675 6245
rect 4617 6236 4629 6239
rect 4264 6208 4629 6236
rect 4157 6199 4215 6205
rect 4617 6205 4629 6208
rect 4663 6205 4675 6239
rect 4617 6199 4675 6205
rect 4801 6239 4859 6245
rect 4801 6205 4813 6239
rect 4847 6205 4859 6239
rect 4801 6199 4859 6205
rect 3421 6171 3479 6177
rect 3421 6168 3433 6171
rect 2746 6140 3433 6168
rect 1946 6060 1952 6112
rect 2004 6060 2010 6112
rect 2133 6103 2191 6109
rect 2133 6069 2145 6103
rect 2179 6100 2191 6103
rect 2222 6100 2228 6112
rect 2179 6072 2228 6100
rect 2179 6069 2191 6072
rect 2133 6063 2191 6069
rect 2222 6060 2228 6072
rect 2280 6060 2286 6112
rect 2406 6060 2412 6112
rect 2464 6100 2470 6112
rect 2746 6100 2774 6140
rect 3421 6137 3433 6140
rect 3467 6137 3479 6171
rect 4172 6168 4200 6199
rect 5442 6196 5448 6248
rect 5500 6196 5506 6248
rect 5994 6196 6000 6248
rect 6052 6196 6058 6248
rect 6086 6196 6092 6248
rect 6144 6196 6150 6248
rect 6270 6196 6276 6248
rect 6328 6196 6334 6248
rect 6641 6239 6699 6245
rect 6641 6205 6653 6239
rect 6687 6236 6699 6239
rect 6822 6236 6828 6248
rect 6687 6208 6828 6236
rect 6687 6205 6699 6208
rect 6641 6199 6699 6205
rect 6822 6196 6828 6208
rect 6880 6196 6886 6248
rect 6917 6239 6975 6245
rect 6917 6205 6929 6239
rect 6963 6236 6975 6239
rect 7098 6236 7104 6248
rect 6963 6208 7104 6236
rect 6963 6205 6975 6208
rect 6917 6199 6975 6205
rect 4709 6171 4767 6177
rect 4709 6168 4721 6171
rect 4172 6140 4721 6168
rect 3421 6131 3479 6137
rect 4709 6137 4721 6140
rect 4755 6137 4767 6171
rect 6932 6168 6960 6199
rect 7098 6196 7104 6208
rect 7156 6196 7162 6248
rect 7190 6196 7196 6248
rect 7248 6196 7254 6248
rect 7300 6236 7328 6267
rect 7742 6236 7748 6248
rect 7300 6208 7748 6236
rect 7742 6196 7748 6208
rect 7800 6196 7806 6248
rect 7834 6196 7840 6248
rect 7892 6236 7898 6248
rect 8386 6236 8392 6248
rect 7892 6208 8392 6236
rect 7892 6196 7898 6208
rect 8386 6196 8392 6208
rect 8444 6196 8450 6248
rect 8570 6196 8576 6248
rect 8628 6196 8634 6248
rect 8662 6196 8668 6248
rect 8720 6196 8726 6248
rect 8757 6239 8815 6245
rect 8757 6205 8769 6239
rect 8803 6236 8815 6239
rect 8846 6236 8852 6248
rect 8803 6208 8852 6236
rect 8803 6205 8815 6208
rect 8757 6199 8815 6205
rect 8846 6196 8852 6208
rect 8904 6196 8910 6248
rect 8956 6245 8984 6276
rect 9306 6264 9312 6316
rect 9364 6304 9370 6316
rect 11256 6304 11284 6344
rect 11330 6332 11336 6384
rect 11388 6372 11394 6384
rect 14461 6375 14519 6381
rect 14461 6372 14473 6375
rect 11388 6344 14473 6372
rect 11388 6332 11394 6344
rect 12452 6316 12480 6344
rect 14461 6341 14473 6344
rect 14507 6372 14519 6375
rect 14734 6372 14740 6384
rect 14507 6344 14740 6372
rect 14507 6341 14519 6344
rect 14461 6335 14519 6341
rect 14734 6332 14740 6344
rect 14792 6332 14798 6384
rect 14844 6372 14872 6412
rect 14921 6409 14933 6443
rect 14967 6440 14979 6443
rect 15010 6440 15016 6452
rect 14967 6412 15016 6440
rect 14967 6409 14979 6412
rect 14921 6403 14979 6409
rect 15010 6400 15016 6412
rect 15068 6400 15074 6452
rect 19797 6443 19855 6449
rect 19797 6440 19809 6443
rect 15120 6412 19809 6440
rect 15120 6372 15148 6412
rect 19797 6409 19809 6412
rect 19843 6409 19855 6443
rect 19797 6403 19855 6409
rect 19886 6400 19892 6452
rect 19944 6440 19950 6452
rect 20073 6443 20131 6449
rect 20073 6440 20085 6443
rect 19944 6412 20085 6440
rect 19944 6400 19950 6412
rect 20073 6409 20085 6412
rect 20119 6409 20131 6443
rect 20073 6403 20131 6409
rect 20530 6400 20536 6452
rect 20588 6440 20594 6452
rect 20993 6443 21051 6449
rect 20993 6440 21005 6443
rect 20588 6412 21005 6440
rect 20588 6400 20594 6412
rect 20993 6409 21005 6412
rect 21039 6440 21051 6443
rect 21039 6412 22094 6440
rect 21039 6409 21051 6412
rect 20993 6403 21051 6409
rect 16761 6375 16819 6381
rect 16761 6372 16773 6375
rect 14844 6344 14964 6372
rect 14936 6316 14964 6344
rect 15028 6344 15148 6372
rect 16408 6344 16773 6372
rect 12253 6307 12311 6313
rect 12253 6304 12265 6307
rect 9364 6276 11192 6304
rect 11256 6276 12265 6304
rect 9364 6264 9370 6276
rect 8941 6239 8999 6245
rect 8941 6205 8953 6239
rect 8987 6205 8999 6239
rect 8941 6199 8999 6205
rect 9030 6196 9036 6248
rect 9088 6196 9094 6248
rect 9214 6196 9220 6248
rect 9272 6236 9278 6248
rect 9401 6239 9459 6245
rect 9272 6208 9352 6236
rect 9272 6196 9278 6208
rect 4709 6131 4767 6137
rect 6472 6140 6960 6168
rect 2464 6072 2774 6100
rect 4525 6103 4583 6109
rect 2464 6060 2470 6072
rect 4525 6069 4537 6103
rect 4571 6100 4583 6103
rect 6472 6100 6500 6140
rect 7374 6128 7380 6180
rect 7432 6168 7438 6180
rect 9324 6168 9352 6208
rect 9401 6205 9413 6239
rect 9447 6236 9459 6239
rect 9582 6236 9588 6248
rect 9447 6208 9588 6236
rect 9447 6205 9459 6208
rect 9401 6199 9459 6205
rect 9582 6196 9588 6208
rect 9640 6196 9646 6248
rect 11057 6239 11115 6245
rect 11057 6205 11069 6239
rect 11103 6205 11115 6239
rect 11164 6236 11192 6276
rect 12253 6273 12265 6276
rect 12299 6273 12311 6307
rect 12253 6267 12311 6273
rect 12434 6264 12440 6316
rect 12492 6264 12498 6316
rect 14277 6307 14335 6313
rect 14277 6273 14289 6307
rect 14323 6304 14335 6307
rect 14323 6276 14688 6304
rect 14323 6273 14335 6276
rect 14277 6267 14335 6273
rect 14660 6248 14688 6276
rect 14918 6264 14924 6316
rect 14976 6264 14982 6316
rect 11734 6239 11792 6245
rect 11734 6236 11746 6239
rect 11164 6208 11746 6236
rect 11057 6199 11115 6205
rect 11734 6205 11746 6208
rect 11780 6236 11792 6239
rect 13909 6239 13967 6245
rect 11780 6208 11928 6236
rect 11780 6205 11792 6208
rect 11734 6199 11792 6205
rect 10410 6168 10416 6180
rect 7432 6140 9227 6168
rect 9324 6140 10416 6168
rect 7432 6128 7438 6140
rect 4571 6072 6500 6100
rect 4571 6069 4583 6072
rect 4525 6063 4583 6069
rect 6546 6060 6552 6112
rect 6604 6100 6610 6112
rect 6730 6100 6736 6112
rect 6604 6072 6736 6100
rect 6604 6060 6610 6072
rect 6730 6060 6736 6072
rect 6788 6100 6794 6112
rect 6825 6103 6883 6109
rect 6825 6100 6837 6103
rect 6788 6072 6837 6100
rect 6788 6060 6794 6072
rect 6825 6069 6837 6072
rect 6871 6069 6883 6103
rect 6825 6063 6883 6069
rect 8386 6060 8392 6112
rect 8444 6060 8450 6112
rect 9199 6100 9227 6140
rect 10410 6128 10416 6140
rect 10468 6128 10474 6180
rect 11072 6168 11100 6199
rect 11072 6140 11192 6168
rect 11164 6100 11192 6140
rect 11238 6128 11244 6180
rect 11296 6168 11302 6180
rect 11900 6168 11928 6208
rect 13909 6205 13921 6239
rect 13955 6236 13967 6239
rect 13998 6236 14004 6248
rect 13955 6208 14004 6236
rect 13955 6205 13967 6208
rect 13909 6199 13967 6205
rect 13998 6196 14004 6208
rect 14056 6196 14062 6248
rect 14182 6196 14188 6248
rect 14240 6196 14246 6248
rect 14366 6196 14372 6248
rect 14424 6236 14430 6248
rect 14424 6208 14596 6236
rect 14424 6196 14430 6208
rect 13078 6168 13084 6180
rect 11296 6140 11836 6168
rect 11900 6140 13084 6168
rect 11296 6128 11302 6140
rect 11422 6100 11428 6112
rect 9199 6072 11428 6100
rect 11422 6060 11428 6072
rect 11480 6060 11486 6112
rect 11514 6060 11520 6112
rect 11572 6100 11578 6112
rect 11808 6109 11836 6140
rect 13078 6128 13084 6140
rect 13136 6128 13142 6180
rect 14568 6168 14596 6208
rect 14642 6196 14648 6248
rect 14700 6196 14706 6248
rect 15028 6168 15056 6344
rect 15102 6264 15108 6316
rect 15160 6304 15166 6316
rect 15160 6276 15700 6304
rect 15160 6264 15166 6276
rect 15194 6196 15200 6248
rect 15252 6196 15258 6248
rect 15304 6245 15332 6276
rect 15289 6239 15347 6245
rect 15289 6205 15301 6239
rect 15335 6205 15347 6239
rect 15289 6199 15347 6205
rect 15381 6239 15439 6245
rect 15381 6205 15393 6239
rect 15427 6205 15439 6239
rect 15381 6199 15439 6205
rect 14568 6140 15056 6168
rect 15396 6168 15424 6199
rect 15562 6196 15568 6248
rect 15620 6196 15626 6248
rect 15672 6245 15700 6276
rect 15930 6264 15936 6316
rect 15988 6304 15994 6316
rect 16117 6307 16175 6313
rect 16117 6304 16129 6307
rect 15988 6276 16129 6304
rect 15988 6264 15994 6276
rect 16117 6273 16129 6276
rect 16163 6273 16175 6307
rect 16117 6267 16175 6273
rect 16206 6264 16212 6316
rect 16264 6264 16270 6316
rect 16408 6313 16436 6344
rect 16761 6341 16773 6344
rect 16807 6341 16819 6375
rect 17954 6372 17960 6384
rect 16761 6335 16819 6341
rect 17420 6344 17960 6372
rect 17420 6313 17448 6344
rect 17954 6332 17960 6344
rect 18012 6332 18018 6384
rect 18138 6332 18144 6384
rect 18196 6372 18202 6384
rect 21174 6372 21180 6384
rect 18196 6344 21180 6372
rect 18196 6332 18202 6344
rect 16393 6307 16451 6313
rect 16393 6273 16405 6307
rect 16439 6273 16451 6307
rect 16393 6267 16451 6273
rect 17405 6307 17463 6313
rect 17405 6273 17417 6307
rect 17451 6273 17463 6307
rect 17405 6267 17463 6273
rect 17865 6307 17923 6313
rect 17865 6273 17877 6307
rect 17911 6304 17923 6307
rect 18322 6304 18328 6316
rect 17911 6276 18328 6304
rect 17911 6273 17923 6276
rect 17865 6267 17923 6273
rect 18322 6264 18328 6276
rect 18380 6304 18386 6316
rect 18874 6304 18880 6316
rect 18380 6276 18880 6304
rect 18380 6264 18386 6276
rect 18874 6264 18880 6276
rect 18932 6264 18938 6316
rect 19168 6313 19196 6344
rect 21174 6332 21180 6344
rect 21232 6332 21238 6384
rect 21821 6375 21879 6381
rect 21821 6341 21833 6375
rect 21867 6341 21879 6375
rect 21821 6335 21879 6341
rect 19153 6307 19211 6313
rect 19153 6273 19165 6307
rect 19199 6273 19211 6307
rect 19153 6267 19211 6273
rect 19245 6307 19303 6313
rect 19245 6273 19257 6307
rect 19291 6273 19303 6307
rect 20530 6304 20536 6316
rect 19245 6267 19303 6273
rect 19812 6276 20536 6304
rect 15657 6239 15715 6245
rect 15657 6205 15669 6239
rect 15703 6205 15715 6239
rect 15657 6199 15715 6205
rect 15838 6196 15844 6248
rect 15896 6196 15902 6248
rect 16298 6196 16304 6248
rect 16356 6196 16362 6248
rect 16482 6196 16488 6248
rect 16540 6236 16546 6248
rect 16540 6208 18276 6236
rect 16540 6196 16546 6208
rect 15749 6171 15807 6177
rect 15749 6168 15761 6171
rect 15396 6140 15761 6168
rect 15749 6137 15761 6140
rect 15795 6137 15807 6171
rect 17221 6171 17279 6177
rect 17221 6168 17233 6171
rect 15749 6131 15807 6137
rect 15856 6140 17233 6168
rect 11609 6103 11667 6109
rect 11609 6100 11621 6103
rect 11572 6072 11621 6100
rect 11572 6060 11578 6072
rect 11609 6069 11621 6072
rect 11655 6069 11667 6103
rect 11609 6063 11667 6069
rect 11793 6103 11851 6109
rect 11793 6069 11805 6103
rect 11839 6100 11851 6103
rect 11974 6100 11980 6112
rect 11839 6072 11980 6100
rect 11839 6069 11851 6072
rect 11793 6063 11851 6069
rect 11974 6060 11980 6072
rect 12032 6060 12038 6112
rect 14642 6060 14648 6112
rect 14700 6100 14706 6112
rect 15856 6100 15884 6140
rect 17221 6137 17233 6140
rect 17267 6168 17279 6171
rect 18141 6171 18199 6177
rect 18141 6168 18153 6171
rect 17267 6140 18153 6168
rect 17267 6137 17279 6140
rect 17221 6131 17279 6137
rect 18141 6137 18153 6140
rect 18187 6137 18199 6171
rect 18248 6168 18276 6208
rect 18782 6196 18788 6248
rect 18840 6236 18846 6248
rect 19260 6236 19288 6267
rect 19812 6245 19840 6276
rect 20272 6245 20300 6276
rect 20530 6264 20536 6276
rect 20588 6264 20594 6316
rect 21836 6304 21864 6335
rect 21192 6276 21864 6304
rect 22066 6304 22094 6412
rect 22373 6307 22431 6313
rect 22373 6304 22385 6307
rect 22066 6276 22385 6304
rect 21192 6245 21220 6276
rect 22373 6273 22385 6276
rect 22419 6273 22431 6307
rect 22373 6267 22431 6273
rect 18840 6208 19288 6236
rect 19797 6239 19855 6245
rect 18840 6196 18846 6208
rect 19797 6205 19809 6239
rect 19843 6205 19855 6239
rect 19797 6199 19855 6205
rect 19981 6239 20039 6245
rect 19981 6205 19993 6239
rect 20027 6236 20039 6239
rect 20257 6239 20315 6245
rect 20027 6208 20116 6236
rect 20027 6205 20039 6208
rect 19981 6199 20039 6205
rect 18248 6140 19840 6168
rect 18141 6131 18199 6137
rect 19812 6112 19840 6140
rect 14700 6072 15884 6100
rect 14700 6060 14706 6072
rect 15930 6060 15936 6112
rect 15988 6060 15994 6112
rect 17126 6060 17132 6112
rect 17184 6100 17190 6112
rect 18049 6103 18107 6109
rect 18049 6100 18061 6103
rect 17184 6072 18061 6100
rect 17184 6060 17190 6072
rect 18049 6069 18061 6072
rect 18095 6069 18107 6103
rect 18049 6063 18107 6069
rect 18506 6060 18512 6112
rect 18564 6060 18570 6112
rect 18690 6060 18696 6112
rect 18748 6060 18754 6112
rect 19058 6060 19064 6112
rect 19116 6060 19122 6112
rect 19794 6060 19800 6112
rect 19852 6060 19858 6112
rect 20088 6100 20116 6208
rect 20257 6205 20269 6239
rect 20303 6205 20315 6239
rect 20901 6239 20959 6245
rect 20901 6236 20913 6239
rect 20257 6199 20315 6205
rect 20548 6208 20913 6236
rect 20162 6128 20168 6180
rect 20220 6168 20226 6180
rect 20548 6168 20576 6208
rect 20901 6205 20913 6208
rect 20947 6205 20959 6239
rect 20901 6199 20959 6205
rect 21177 6239 21235 6245
rect 21177 6205 21189 6239
rect 21223 6205 21235 6239
rect 21177 6199 21235 6205
rect 21269 6239 21327 6245
rect 21269 6205 21281 6239
rect 21315 6205 21327 6239
rect 21269 6199 21327 6205
rect 20220 6140 20576 6168
rect 20220 6128 20226 6140
rect 20622 6128 20628 6180
rect 20680 6168 20686 6180
rect 21284 6168 21312 6199
rect 20680 6140 21312 6168
rect 20680 6128 20686 6140
rect 20898 6100 20904 6112
rect 20088 6072 20904 6100
rect 20898 6060 20904 6072
rect 20956 6060 20962 6112
rect 21266 6060 21272 6112
rect 21324 6100 21330 6112
rect 21453 6103 21511 6109
rect 21453 6100 21465 6103
rect 21324 6072 21465 6100
rect 21324 6060 21330 6072
rect 21453 6069 21465 6072
rect 21499 6069 21511 6103
rect 21453 6063 21511 6069
rect 22186 6060 22192 6112
rect 22244 6060 22250 6112
rect 22278 6060 22284 6112
rect 22336 6060 22342 6112
rect 552 6010 23368 6032
rect 552 5958 4366 6010
rect 4418 5958 4430 6010
rect 4482 5958 4494 6010
rect 4546 5958 4558 6010
rect 4610 5958 4622 6010
rect 4674 5958 4686 6010
rect 4738 5958 10366 6010
rect 10418 5958 10430 6010
rect 10482 5958 10494 6010
rect 10546 5958 10558 6010
rect 10610 5958 10622 6010
rect 10674 5958 10686 6010
rect 10738 5958 16366 6010
rect 16418 5958 16430 6010
rect 16482 5958 16494 6010
rect 16546 5958 16558 6010
rect 16610 5958 16622 6010
rect 16674 5958 16686 6010
rect 16738 5958 22366 6010
rect 22418 5958 22430 6010
rect 22482 5958 22494 6010
rect 22546 5958 22558 6010
rect 22610 5958 22622 6010
rect 22674 5958 22686 6010
rect 22738 5958 23368 6010
rect 552 5936 23368 5958
rect 2685 5899 2743 5905
rect 2685 5865 2697 5899
rect 2731 5865 2743 5899
rect 2685 5859 2743 5865
rect 3467 5899 3525 5905
rect 3467 5865 3479 5899
rect 3513 5896 3525 5899
rect 3970 5896 3976 5908
rect 3513 5868 3976 5896
rect 3513 5865 3525 5868
rect 3467 5859 3525 5865
rect 2700 5828 2728 5859
rect 3970 5856 3976 5868
rect 4028 5856 4034 5908
rect 4154 5856 4160 5908
rect 4212 5896 4218 5908
rect 4433 5899 4491 5905
rect 4433 5896 4445 5899
rect 4212 5868 4445 5896
rect 4212 5856 4218 5868
rect 4433 5865 4445 5868
rect 4479 5865 4491 5899
rect 4433 5859 4491 5865
rect 5166 5856 5172 5908
rect 5224 5896 5230 5908
rect 6270 5896 6276 5908
rect 5224 5868 6276 5896
rect 5224 5856 5230 5868
rect 6270 5856 6276 5868
rect 6328 5856 6334 5908
rect 6730 5856 6736 5908
rect 6788 5896 6794 5908
rect 7742 5896 7748 5908
rect 6788 5868 7748 5896
rect 6788 5856 6794 5868
rect 7742 5856 7748 5868
rect 7800 5856 7806 5908
rect 8389 5899 8447 5905
rect 8389 5865 8401 5899
rect 8435 5896 8447 5899
rect 8846 5896 8852 5908
rect 8435 5868 8852 5896
rect 8435 5865 8447 5868
rect 8389 5859 8447 5865
rect 8846 5856 8852 5868
rect 8904 5856 8910 5908
rect 12986 5896 12992 5908
rect 8956 5868 12992 5896
rect 5350 5828 5356 5840
rect 2700 5800 5356 5828
rect 5350 5788 5356 5800
rect 5408 5828 5414 5840
rect 6086 5828 6092 5840
rect 5408 5800 6092 5828
rect 5408 5788 5414 5800
rect 6086 5788 6092 5800
rect 6144 5788 6150 5840
rect 7190 5788 7196 5840
rect 7248 5828 7254 5840
rect 8110 5828 8116 5840
rect 7248 5800 8116 5828
rect 7248 5788 7254 5800
rect 8110 5788 8116 5800
rect 8168 5788 8174 5840
rect 1029 5763 1087 5769
rect 1029 5729 1041 5763
rect 1075 5760 1087 5763
rect 1489 5763 1547 5769
rect 1489 5760 1501 5763
rect 1075 5732 1501 5760
rect 1075 5729 1087 5732
rect 1029 5723 1087 5729
rect 1489 5729 1501 5732
rect 1535 5729 1547 5763
rect 1489 5723 1547 5729
rect 1673 5763 1731 5769
rect 1673 5729 1685 5763
rect 1719 5760 1731 5763
rect 1762 5760 1768 5772
rect 1719 5732 1768 5760
rect 1719 5729 1731 5732
rect 1673 5723 1731 5729
rect 1762 5720 1768 5732
rect 1820 5720 1826 5772
rect 1946 5720 1952 5772
rect 2004 5760 2010 5772
rect 2317 5763 2375 5769
rect 2317 5760 2329 5763
rect 2004 5732 2329 5760
rect 2004 5720 2010 5732
rect 2317 5729 2329 5732
rect 2363 5729 2375 5763
rect 2317 5723 2375 5729
rect 2498 5720 2504 5772
rect 2556 5760 2562 5772
rect 3697 5763 3755 5769
rect 3697 5760 3709 5763
rect 2556 5732 3709 5760
rect 2556 5720 2562 5732
rect 3697 5729 3709 5732
rect 3743 5729 3755 5763
rect 3697 5723 3755 5729
rect 3786 5720 3792 5772
rect 3844 5720 3850 5772
rect 3970 5720 3976 5772
rect 4028 5760 4034 5772
rect 4157 5763 4215 5769
rect 4157 5760 4169 5763
rect 4028 5732 4169 5760
rect 4028 5720 4034 5732
rect 4157 5729 4169 5732
rect 4203 5729 4215 5763
rect 4157 5723 4215 5729
rect 4341 5763 4399 5769
rect 4341 5729 4353 5763
rect 4387 5729 4399 5763
rect 4341 5723 4399 5729
rect 4433 5763 4491 5769
rect 4433 5729 4445 5763
rect 4479 5760 4491 5763
rect 4522 5760 4528 5772
rect 4479 5732 4528 5760
rect 4479 5729 4491 5732
rect 4433 5723 4491 5729
rect 842 5652 848 5704
rect 900 5692 906 5704
rect 937 5695 995 5701
rect 937 5692 949 5695
rect 900 5664 949 5692
rect 900 5652 906 5664
rect 937 5661 949 5664
rect 983 5661 995 5695
rect 937 5655 995 5661
rect 1857 5695 1915 5701
rect 1857 5661 1869 5695
rect 1903 5692 1915 5695
rect 2406 5692 2412 5704
rect 1903 5664 2412 5692
rect 1903 5661 1915 5664
rect 1857 5655 1915 5661
rect 2406 5652 2412 5664
rect 2464 5652 2470 5704
rect 2866 5652 2872 5704
rect 2924 5692 2930 5704
rect 3804 5692 3832 5720
rect 2924 5664 3832 5692
rect 2924 5652 2930 5664
rect 4356 5636 4384 5723
rect 4522 5720 4528 5732
rect 4580 5720 4586 5772
rect 4614 5720 4620 5772
rect 4672 5720 4678 5772
rect 4798 5720 4804 5772
rect 4856 5760 4862 5772
rect 5169 5763 5227 5769
rect 5169 5760 5181 5763
rect 4856 5732 5181 5760
rect 4856 5720 4862 5732
rect 5169 5729 5181 5732
rect 5215 5729 5227 5763
rect 5169 5723 5227 5729
rect 5534 5720 5540 5772
rect 5592 5760 5598 5772
rect 5813 5763 5871 5769
rect 5813 5760 5825 5763
rect 5592 5732 5825 5760
rect 5592 5720 5598 5732
rect 5813 5729 5825 5732
rect 5859 5729 5871 5763
rect 5813 5723 5871 5729
rect 5902 5720 5908 5772
rect 5960 5760 5966 5772
rect 6273 5763 6331 5769
rect 6273 5760 6285 5763
rect 5960 5732 6285 5760
rect 5960 5720 5966 5732
rect 6273 5729 6285 5732
rect 6319 5729 6331 5763
rect 6273 5723 6331 5729
rect 6454 5720 6460 5772
rect 6512 5760 6518 5772
rect 6825 5763 6883 5769
rect 6825 5760 6837 5763
rect 6512 5732 6837 5760
rect 6512 5720 6518 5732
rect 6825 5729 6837 5732
rect 6871 5729 6883 5763
rect 6825 5723 6883 5729
rect 8021 5763 8079 5769
rect 8021 5729 8033 5763
rect 8067 5760 8079 5763
rect 8128 5760 8156 5788
rect 8067 5732 8156 5760
rect 8067 5729 8079 5732
rect 8021 5723 8079 5729
rect 8202 5720 8208 5772
rect 8260 5720 8266 5772
rect 8478 5720 8484 5772
rect 8536 5720 8542 5772
rect 8956 5769 8984 5868
rect 12986 5856 12992 5868
rect 13044 5856 13050 5908
rect 13078 5856 13084 5908
rect 13136 5896 13142 5908
rect 13357 5899 13415 5905
rect 13357 5896 13369 5899
rect 13136 5868 13369 5896
rect 13136 5856 13142 5868
rect 13357 5865 13369 5868
rect 13403 5865 13415 5899
rect 13357 5859 13415 5865
rect 13909 5899 13967 5905
rect 13909 5865 13921 5899
rect 13955 5896 13967 5899
rect 14642 5896 14648 5908
rect 13955 5868 14648 5896
rect 13955 5865 13967 5868
rect 13909 5859 13967 5865
rect 9033 5831 9091 5837
rect 9033 5797 9045 5831
rect 9079 5828 9091 5831
rect 9079 5800 9720 5828
rect 9079 5797 9091 5800
rect 9033 5791 9091 5797
rect 8941 5763 8999 5769
rect 8941 5729 8953 5763
rect 8987 5729 8999 5763
rect 8941 5723 8999 5729
rect 9125 5763 9183 5769
rect 9125 5729 9137 5763
rect 9171 5760 9183 5763
rect 9398 5760 9404 5772
rect 9171 5732 9404 5760
rect 9171 5729 9183 5732
rect 9125 5723 9183 5729
rect 9398 5720 9404 5732
rect 9456 5720 9462 5772
rect 9692 5769 9720 5800
rect 9493 5763 9551 5769
rect 9493 5729 9505 5763
rect 9539 5729 9551 5763
rect 9493 5723 9551 5729
rect 9677 5763 9735 5769
rect 9677 5729 9689 5763
rect 9723 5729 9735 5763
rect 9677 5723 9735 5729
rect 9769 5763 9827 5769
rect 9769 5729 9781 5763
rect 9815 5729 9827 5763
rect 9769 5723 9827 5729
rect 5074 5652 5080 5704
rect 5132 5652 5138 5704
rect 5552 5692 5580 5720
rect 5184 5664 5580 5692
rect 1397 5627 1455 5633
rect 1397 5593 1409 5627
rect 1443 5624 1455 5627
rect 1946 5624 1952 5636
rect 1443 5596 1952 5624
rect 1443 5593 1455 5596
rect 1397 5587 1455 5593
rect 1946 5584 1952 5596
rect 2004 5584 2010 5636
rect 4338 5584 4344 5636
rect 4396 5624 4402 5636
rect 5184 5624 5212 5664
rect 6362 5652 6368 5704
rect 6420 5692 6426 5704
rect 6549 5695 6607 5701
rect 6549 5692 6561 5695
rect 6420 5664 6561 5692
rect 6420 5652 6426 5664
rect 6549 5661 6561 5664
rect 6595 5661 6607 5695
rect 6549 5655 6607 5661
rect 6638 5652 6644 5704
rect 6696 5692 6702 5704
rect 6733 5695 6791 5701
rect 6733 5692 6745 5695
rect 6696 5664 6745 5692
rect 6696 5652 6702 5664
rect 6733 5661 6745 5664
rect 6779 5661 6791 5695
rect 6733 5655 6791 5661
rect 7006 5652 7012 5704
rect 7064 5692 7070 5704
rect 7193 5695 7251 5701
rect 7193 5692 7205 5695
rect 7064 5664 7205 5692
rect 7064 5652 7070 5664
rect 7193 5661 7205 5664
rect 7239 5661 7251 5695
rect 7193 5655 7251 5661
rect 7929 5695 7987 5701
rect 7929 5661 7941 5695
rect 7975 5661 7987 5695
rect 7929 5655 7987 5661
rect 4396 5596 5212 5624
rect 4396 5584 4402 5596
rect 5534 5584 5540 5636
rect 5592 5584 5598 5636
rect 5994 5584 6000 5636
rect 6052 5624 6058 5636
rect 7374 5624 7380 5636
rect 6052 5596 7380 5624
rect 6052 5584 6058 5596
rect 7374 5584 7380 5596
rect 7432 5584 7438 5636
rect 3970 5516 3976 5568
rect 4028 5516 4034 5568
rect 4246 5516 4252 5568
rect 4304 5556 4310 5568
rect 4522 5556 4528 5568
rect 4304 5528 4528 5556
rect 4304 5516 4310 5528
rect 4522 5516 4528 5528
rect 4580 5516 4586 5568
rect 6362 5516 6368 5568
rect 6420 5516 6426 5568
rect 6457 5559 6515 5565
rect 6457 5525 6469 5559
rect 6503 5556 6515 5559
rect 6914 5556 6920 5568
rect 6503 5528 6920 5556
rect 6503 5525 6515 5528
rect 6457 5519 6515 5525
rect 6914 5516 6920 5528
rect 6972 5516 6978 5568
rect 7944 5556 7972 5655
rect 8110 5652 8116 5704
rect 8168 5652 8174 5704
rect 8573 5695 8631 5701
rect 8573 5661 8585 5695
rect 8619 5692 8631 5695
rect 8662 5692 8668 5704
rect 8619 5664 8668 5692
rect 8619 5661 8631 5664
rect 8573 5655 8631 5661
rect 8662 5652 8668 5664
rect 8720 5652 8726 5704
rect 9217 5627 9275 5633
rect 9217 5624 9229 5627
rect 8220 5596 9229 5624
rect 8220 5556 8248 5596
rect 9217 5593 9229 5596
rect 9263 5593 9275 5627
rect 9508 5624 9536 5723
rect 9784 5692 9812 5723
rect 9950 5720 9956 5772
rect 10008 5720 10014 5772
rect 10410 5720 10416 5772
rect 10468 5720 10474 5772
rect 11149 5763 11207 5769
rect 11149 5729 11161 5763
rect 11195 5760 11207 5763
rect 11330 5760 11336 5772
rect 11195 5732 11336 5760
rect 11195 5729 11207 5732
rect 11149 5723 11207 5729
rect 11330 5720 11336 5732
rect 11388 5720 11394 5772
rect 11422 5720 11428 5772
rect 11480 5720 11486 5772
rect 11514 5720 11520 5772
rect 11572 5720 11578 5772
rect 11882 5720 11888 5772
rect 11940 5760 11946 5772
rect 11977 5763 12035 5769
rect 11977 5760 11989 5763
rect 11940 5732 11989 5760
rect 11940 5720 11946 5732
rect 11977 5729 11989 5732
rect 12023 5729 12035 5763
rect 11977 5723 12035 5729
rect 12066 5720 12072 5772
rect 12124 5720 12130 5772
rect 12253 5763 12311 5769
rect 12253 5729 12265 5763
rect 12299 5760 12311 5763
rect 12710 5760 12716 5772
rect 12299 5732 12716 5760
rect 12299 5729 12311 5732
rect 12253 5723 12311 5729
rect 12710 5720 12716 5732
rect 12768 5720 12774 5772
rect 12897 5763 12955 5769
rect 12897 5729 12909 5763
rect 12943 5729 12955 5763
rect 12897 5723 12955 5729
rect 12989 5763 13047 5769
rect 12989 5729 13001 5763
rect 13035 5760 13047 5763
rect 13541 5763 13599 5769
rect 13541 5760 13553 5763
rect 13035 5732 13553 5760
rect 13035 5729 13047 5732
rect 12989 5723 13047 5729
rect 13541 5729 13553 5732
rect 13587 5760 13599 5763
rect 13924 5760 13952 5859
rect 14642 5856 14648 5868
rect 14700 5856 14706 5908
rect 15102 5856 15108 5908
rect 15160 5856 15166 5908
rect 15565 5899 15623 5905
rect 15565 5865 15577 5899
rect 15611 5896 15623 5899
rect 15838 5896 15844 5908
rect 15611 5868 15844 5896
rect 15611 5865 15623 5868
rect 15565 5859 15623 5865
rect 15838 5856 15844 5868
rect 15896 5896 15902 5908
rect 19058 5896 19064 5908
rect 15896 5868 19064 5896
rect 15896 5856 15902 5868
rect 19058 5856 19064 5868
rect 19116 5896 19122 5908
rect 22278 5896 22284 5908
rect 19116 5868 22284 5896
rect 19116 5856 19122 5868
rect 22278 5856 22284 5868
rect 22336 5896 22342 5908
rect 22373 5899 22431 5905
rect 22373 5896 22385 5899
rect 22336 5868 22385 5896
rect 22336 5856 22342 5868
rect 22373 5865 22385 5868
rect 22419 5865 22431 5899
rect 22373 5859 22431 5865
rect 14921 5831 14979 5837
rect 14921 5797 14933 5831
rect 14967 5828 14979 5831
rect 15120 5828 15148 5856
rect 14967 5800 15148 5828
rect 15304 5800 16528 5828
rect 14967 5797 14979 5800
rect 14921 5791 14979 5797
rect 13587 5732 13952 5760
rect 13587 5729 13599 5732
rect 13541 5723 13599 5729
rect 10045 5695 10103 5701
rect 10045 5692 10057 5695
rect 9784 5664 10057 5692
rect 10045 5661 10057 5664
rect 10091 5692 10103 5695
rect 10505 5695 10563 5701
rect 10505 5692 10517 5695
rect 10091 5664 10517 5692
rect 10091 5661 10103 5664
rect 10045 5655 10103 5661
rect 10505 5661 10517 5664
rect 10551 5692 10563 5695
rect 11900 5692 11928 5720
rect 10551 5664 11928 5692
rect 12912 5692 12940 5723
rect 13998 5720 14004 5772
rect 14056 5760 14062 5772
rect 14093 5763 14151 5769
rect 14093 5760 14105 5763
rect 14056 5732 14105 5760
rect 14056 5720 14062 5732
rect 14093 5729 14105 5732
rect 14139 5729 14151 5763
rect 14093 5723 14151 5729
rect 13173 5695 13231 5701
rect 12912 5664 13124 5692
rect 10551 5661 10563 5664
rect 10505 5655 10563 5661
rect 9766 5624 9772 5636
rect 9508 5596 9772 5624
rect 9217 5587 9275 5593
rect 9766 5584 9772 5596
rect 9824 5584 9830 5636
rect 10321 5627 10379 5633
rect 10321 5593 10333 5627
rect 10367 5624 10379 5627
rect 10962 5624 10968 5636
rect 10367 5596 10968 5624
rect 10367 5593 10379 5596
rect 10321 5587 10379 5593
rect 10962 5584 10968 5596
rect 11020 5584 11026 5636
rect 11238 5584 11244 5636
rect 11296 5584 11302 5636
rect 11606 5584 11612 5636
rect 11664 5624 11670 5636
rect 11793 5627 11851 5633
rect 11793 5624 11805 5627
rect 11664 5596 11805 5624
rect 11664 5584 11670 5596
rect 11793 5593 11805 5596
rect 11839 5593 11851 5627
rect 11793 5587 11851 5593
rect 12161 5627 12219 5633
rect 12161 5593 12173 5627
rect 12207 5624 12219 5627
rect 12529 5627 12587 5633
rect 12529 5624 12541 5627
rect 12207 5596 12541 5624
rect 12207 5593 12219 5596
rect 12161 5587 12219 5593
rect 12529 5593 12541 5596
rect 12575 5593 12587 5627
rect 13096 5624 13124 5664
rect 13173 5661 13185 5695
rect 13219 5692 13231 5695
rect 13262 5692 13268 5704
rect 13219 5664 13268 5692
rect 13219 5661 13231 5664
rect 13173 5655 13231 5661
rect 13262 5652 13268 5664
rect 13320 5652 13326 5704
rect 14108 5692 14136 5723
rect 14366 5720 14372 5772
rect 14424 5720 14430 5772
rect 14461 5763 14519 5769
rect 14461 5729 14473 5763
rect 14507 5729 14519 5763
rect 14461 5723 14519 5729
rect 15105 5763 15163 5769
rect 15105 5729 15117 5763
rect 15151 5760 15163 5763
rect 15304 5760 15332 5800
rect 15151 5732 15332 5760
rect 15381 5763 15439 5769
rect 15151 5729 15163 5732
rect 15105 5723 15163 5729
rect 15381 5729 15393 5763
rect 15427 5729 15439 5763
rect 16500 5760 16528 5800
rect 16574 5788 16580 5840
rect 16632 5828 16638 5840
rect 16850 5828 16856 5840
rect 16632 5800 16856 5828
rect 16632 5788 16638 5800
rect 16850 5788 16856 5800
rect 16908 5788 16914 5840
rect 18690 5828 18696 5840
rect 17972 5800 18696 5828
rect 17972 5769 18000 5800
rect 18690 5788 18696 5800
rect 18748 5788 18754 5840
rect 19978 5828 19984 5840
rect 19352 5800 19984 5828
rect 17037 5763 17095 5769
rect 17037 5760 17049 5763
rect 16500 5732 17049 5760
rect 15381 5723 15439 5729
rect 17037 5729 17049 5732
rect 17083 5760 17095 5763
rect 17773 5763 17831 5769
rect 17773 5760 17785 5763
rect 17083 5732 17785 5760
rect 17083 5729 17095 5732
rect 17037 5723 17095 5729
rect 17773 5729 17785 5732
rect 17819 5729 17831 5763
rect 17773 5723 17831 5729
rect 17957 5763 18015 5769
rect 17957 5729 17969 5763
rect 18003 5729 18015 5763
rect 17957 5723 18015 5729
rect 14476 5692 14504 5723
rect 14108 5664 14504 5692
rect 14734 5652 14740 5704
rect 14792 5692 14798 5704
rect 15396 5692 15424 5723
rect 14792 5664 15424 5692
rect 14792 5652 14798 5664
rect 15562 5652 15568 5704
rect 15620 5692 15626 5704
rect 17788 5692 17816 5723
rect 18046 5720 18052 5772
rect 18104 5720 18110 5772
rect 18414 5720 18420 5772
rect 18472 5760 18478 5772
rect 18509 5763 18567 5769
rect 18509 5760 18521 5763
rect 18472 5732 18521 5760
rect 18472 5720 18478 5732
rect 18509 5729 18521 5732
rect 18555 5729 18567 5763
rect 18509 5723 18567 5729
rect 18598 5720 18604 5772
rect 18656 5720 18662 5772
rect 19150 5720 19156 5772
rect 19208 5720 19214 5772
rect 19352 5769 19380 5800
rect 19978 5788 19984 5800
rect 20036 5828 20042 5840
rect 20036 5800 20668 5828
rect 20036 5788 20042 5800
rect 19337 5763 19395 5769
rect 19337 5729 19349 5763
rect 19383 5729 19395 5763
rect 19337 5723 19395 5729
rect 19426 5720 19432 5772
rect 19484 5720 19490 5772
rect 19518 5720 19524 5772
rect 19576 5720 19582 5772
rect 20162 5760 20168 5772
rect 19628 5732 20168 5760
rect 19628 5692 19656 5732
rect 20162 5720 20168 5732
rect 20220 5720 20226 5772
rect 20640 5769 20668 5800
rect 21174 5788 21180 5840
rect 21232 5828 21238 5840
rect 22186 5828 22192 5840
rect 21232 5800 22192 5828
rect 21232 5788 21238 5800
rect 22186 5788 22192 5800
rect 22244 5828 22250 5840
rect 22465 5831 22523 5837
rect 22465 5828 22477 5831
rect 22244 5800 22477 5828
rect 22244 5788 22250 5800
rect 22465 5797 22477 5800
rect 22511 5797 22523 5831
rect 22465 5791 22523 5797
rect 20625 5763 20683 5769
rect 20625 5729 20637 5763
rect 20671 5760 20683 5763
rect 20717 5763 20775 5769
rect 20717 5760 20729 5763
rect 20671 5732 20729 5760
rect 20671 5729 20683 5732
rect 20625 5723 20683 5729
rect 20717 5729 20729 5732
rect 20763 5729 20775 5763
rect 20717 5723 20775 5729
rect 20898 5720 20904 5772
rect 20956 5720 20962 5772
rect 21450 5720 21456 5772
rect 21508 5760 21514 5772
rect 21634 5760 21640 5772
rect 21508 5732 21640 5760
rect 21508 5720 21514 5732
rect 21634 5720 21640 5732
rect 21692 5760 21698 5772
rect 21692 5732 22094 5760
rect 21692 5720 21698 5732
rect 15620 5664 17724 5692
rect 17788 5664 19656 5692
rect 19705 5695 19763 5701
rect 15620 5652 15626 5664
rect 14366 5624 14372 5636
rect 13096 5596 14372 5624
rect 12529 5587 12587 5593
rect 14366 5584 14372 5596
rect 14424 5624 14430 5636
rect 17126 5624 17132 5636
rect 14424 5596 17132 5624
rect 14424 5584 14430 5596
rect 17126 5584 17132 5596
rect 17184 5584 17190 5636
rect 17696 5624 17724 5664
rect 19705 5661 19717 5695
rect 19751 5661 19763 5695
rect 19705 5655 19763 5661
rect 18598 5624 18604 5636
rect 17696 5596 18604 5624
rect 18598 5584 18604 5596
rect 18656 5624 18662 5636
rect 19245 5627 19303 5633
rect 19245 5624 19257 5627
rect 18656 5596 19257 5624
rect 18656 5584 18662 5596
rect 19245 5593 19257 5596
rect 19291 5593 19303 5627
rect 19720 5624 19748 5655
rect 20254 5652 20260 5704
rect 20312 5692 20318 5704
rect 20349 5695 20407 5701
rect 20349 5692 20361 5695
rect 20312 5664 20361 5692
rect 20312 5652 20318 5664
rect 20349 5661 20361 5664
rect 20395 5661 20407 5695
rect 20349 5655 20407 5661
rect 20714 5624 20720 5636
rect 19720 5596 20720 5624
rect 19245 5587 19303 5593
rect 20714 5584 20720 5596
rect 20772 5584 20778 5636
rect 22066 5624 22094 5732
rect 22557 5695 22615 5701
rect 22557 5661 22569 5695
rect 22603 5661 22615 5695
rect 22557 5655 22615 5661
rect 22572 5624 22600 5655
rect 22066 5596 22600 5624
rect 7944 5528 8248 5556
rect 8570 5516 8576 5568
rect 8628 5516 8634 5568
rect 8846 5516 8852 5568
rect 8904 5516 8910 5568
rect 8938 5516 8944 5568
rect 8996 5556 9002 5568
rect 9953 5559 10011 5565
rect 9953 5556 9965 5559
rect 8996 5528 9965 5556
rect 8996 5516 9002 5528
rect 9953 5525 9965 5528
rect 9999 5525 10011 5559
rect 9953 5519 10011 5525
rect 10134 5516 10140 5568
rect 10192 5556 10198 5568
rect 10413 5559 10471 5565
rect 10413 5556 10425 5559
rect 10192 5528 10425 5556
rect 10192 5516 10198 5528
rect 10413 5525 10425 5528
rect 10459 5525 10471 5559
rect 10413 5519 10471 5525
rect 10778 5516 10784 5568
rect 10836 5516 10842 5568
rect 11698 5516 11704 5568
rect 11756 5516 11762 5568
rect 13906 5516 13912 5568
rect 13964 5556 13970 5568
rect 14185 5559 14243 5565
rect 14185 5556 14197 5559
rect 13964 5528 14197 5556
rect 13964 5516 13970 5528
rect 14185 5525 14197 5528
rect 14231 5525 14243 5559
rect 14185 5519 14243 5525
rect 14458 5516 14464 5568
rect 14516 5556 14522 5568
rect 14645 5559 14703 5565
rect 14645 5556 14657 5559
rect 14516 5528 14657 5556
rect 14516 5516 14522 5528
rect 14645 5525 14657 5528
rect 14691 5525 14703 5559
rect 14645 5519 14703 5525
rect 15194 5516 15200 5568
rect 15252 5556 15258 5568
rect 15289 5559 15347 5565
rect 15289 5556 15301 5559
rect 15252 5528 15301 5556
rect 15252 5516 15258 5528
rect 15289 5525 15301 5528
rect 15335 5525 15347 5559
rect 15289 5519 15347 5525
rect 17218 5516 17224 5568
rect 17276 5516 17282 5568
rect 17310 5516 17316 5568
rect 17368 5556 17374 5568
rect 17589 5559 17647 5565
rect 17589 5556 17601 5559
rect 17368 5528 17601 5556
rect 17368 5516 17374 5528
rect 17589 5525 17601 5528
rect 17635 5525 17647 5559
rect 17589 5519 17647 5525
rect 18506 5516 18512 5568
rect 18564 5516 18570 5568
rect 18874 5516 18880 5568
rect 18932 5516 18938 5568
rect 19613 5559 19671 5565
rect 19613 5525 19625 5559
rect 19659 5556 19671 5559
rect 20346 5556 20352 5568
rect 19659 5528 20352 5556
rect 19659 5525 19671 5528
rect 19613 5519 19671 5525
rect 20346 5516 20352 5528
rect 20404 5516 20410 5568
rect 20809 5559 20867 5565
rect 20809 5525 20821 5559
rect 20855 5556 20867 5559
rect 21174 5556 21180 5568
rect 20855 5528 21180 5556
rect 20855 5525 20867 5528
rect 20809 5519 20867 5525
rect 21174 5516 21180 5528
rect 21232 5516 21238 5568
rect 22002 5516 22008 5568
rect 22060 5516 22066 5568
rect 552 5466 23368 5488
rect 552 5414 1366 5466
rect 1418 5414 1430 5466
rect 1482 5414 1494 5466
rect 1546 5414 1558 5466
rect 1610 5414 1622 5466
rect 1674 5414 1686 5466
rect 1738 5414 7366 5466
rect 7418 5414 7430 5466
rect 7482 5414 7494 5466
rect 7546 5414 7558 5466
rect 7610 5414 7622 5466
rect 7674 5414 7686 5466
rect 7738 5414 13366 5466
rect 13418 5414 13430 5466
rect 13482 5414 13494 5466
rect 13546 5414 13558 5466
rect 13610 5414 13622 5466
rect 13674 5414 13686 5466
rect 13738 5414 19366 5466
rect 19418 5414 19430 5466
rect 19482 5414 19494 5466
rect 19546 5414 19558 5466
rect 19610 5414 19622 5466
rect 19674 5414 19686 5466
rect 19738 5414 23368 5466
rect 552 5392 23368 5414
rect 1581 5355 1639 5361
rect 1581 5321 1593 5355
rect 1627 5352 1639 5355
rect 1762 5352 1768 5364
rect 1627 5324 1768 5352
rect 1627 5321 1639 5324
rect 1581 5315 1639 5321
rect 1762 5312 1768 5324
rect 1820 5312 1826 5364
rect 1854 5312 1860 5364
rect 1912 5312 1918 5364
rect 1949 5355 2007 5361
rect 1949 5321 1961 5355
rect 1995 5352 2007 5355
rect 2038 5352 2044 5364
rect 1995 5324 2044 5352
rect 1995 5321 2007 5324
rect 1949 5315 2007 5321
rect 2038 5312 2044 5324
rect 2096 5312 2102 5364
rect 3789 5355 3847 5361
rect 3789 5321 3801 5355
rect 3835 5352 3847 5355
rect 4614 5352 4620 5364
rect 3835 5324 4620 5352
rect 3835 5321 3847 5324
rect 3789 5315 3847 5321
rect 4614 5312 4620 5324
rect 4672 5312 4678 5364
rect 8478 5312 8484 5364
rect 8536 5352 8542 5364
rect 8573 5355 8631 5361
rect 8573 5352 8585 5355
rect 8536 5324 8585 5352
rect 8536 5312 8542 5324
rect 8573 5321 8585 5324
rect 8619 5321 8631 5355
rect 8573 5315 8631 5321
rect 9950 5312 9956 5364
rect 10008 5352 10014 5364
rect 10321 5355 10379 5361
rect 10321 5352 10333 5355
rect 10008 5324 10333 5352
rect 10008 5312 10014 5324
rect 10321 5321 10333 5324
rect 10367 5321 10379 5355
rect 10321 5315 10379 5321
rect 10410 5312 10416 5364
rect 10468 5312 10474 5364
rect 11514 5312 11520 5364
rect 11572 5352 11578 5364
rect 11793 5355 11851 5361
rect 11793 5352 11805 5355
rect 11572 5324 11805 5352
rect 11572 5312 11578 5324
rect 11793 5321 11805 5324
rect 11839 5321 11851 5355
rect 11793 5315 11851 5321
rect 11882 5312 11888 5364
rect 11940 5312 11946 5364
rect 12437 5355 12495 5361
rect 12437 5352 12449 5355
rect 11992 5324 12449 5352
rect 1670 5244 1676 5296
rect 1728 5284 1734 5296
rect 1872 5284 1900 5312
rect 1728 5256 1900 5284
rect 1728 5244 1734 5256
rect 3326 5244 3332 5296
rect 3384 5284 3390 5296
rect 3602 5284 3608 5296
rect 3384 5256 3608 5284
rect 3384 5244 3390 5256
rect 3602 5244 3608 5256
rect 3660 5284 3666 5296
rect 5905 5287 5963 5293
rect 3660 5256 4200 5284
rect 3660 5244 3666 5256
rect 1854 5216 1860 5228
rect 1412 5188 1860 5216
rect 1412 5157 1440 5188
rect 1854 5176 1860 5188
rect 1912 5216 1918 5228
rect 3786 5216 3792 5228
rect 1912 5188 3792 5216
rect 1912 5176 1918 5188
rect 3786 5176 3792 5188
rect 3844 5176 3850 5228
rect 4172 5225 4200 5256
rect 5905 5253 5917 5287
rect 5951 5253 5963 5287
rect 5905 5247 5963 5253
rect 6273 5287 6331 5293
rect 6273 5253 6285 5287
rect 6319 5284 6331 5287
rect 6822 5284 6828 5296
rect 6319 5256 6828 5284
rect 6319 5253 6331 5256
rect 6273 5247 6331 5253
rect 4157 5219 4215 5225
rect 4157 5185 4169 5219
rect 4203 5185 4215 5219
rect 5920 5216 5948 5247
rect 6822 5244 6828 5256
rect 6880 5244 6886 5296
rect 8205 5287 8263 5293
rect 8205 5253 8217 5287
rect 8251 5284 8263 5287
rect 8938 5284 8944 5296
rect 8251 5256 8944 5284
rect 8251 5253 8263 5256
rect 8205 5247 8263 5253
rect 8938 5244 8944 5256
rect 8996 5244 9002 5296
rect 10134 5284 10140 5296
rect 9048 5256 10140 5284
rect 7377 5219 7435 5225
rect 5920 5188 7144 5216
rect 4157 5179 4215 5185
rect 1213 5151 1271 5157
rect 1213 5117 1225 5151
rect 1259 5117 1271 5151
rect 1213 5111 1271 5117
rect 1397 5151 1455 5157
rect 1397 5117 1409 5151
rect 1443 5117 1455 5151
rect 1397 5111 1455 5117
rect 1228 5080 1256 5111
rect 1486 5108 1492 5160
rect 1544 5148 1550 5160
rect 1544 5120 1624 5148
rect 1544 5108 1550 5120
rect 1596 5080 1624 5120
rect 1670 5108 1676 5160
rect 1728 5108 1734 5160
rect 2130 5108 2136 5160
rect 2188 5108 2194 5160
rect 2866 5108 2872 5160
rect 2924 5108 2930 5160
rect 3881 5151 3939 5157
rect 3881 5148 3893 5151
rect 3436 5120 3893 5148
rect 2222 5080 2228 5092
rect 1228 5052 2228 5080
rect 2222 5040 2228 5052
rect 2280 5040 2286 5092
rect 3436 5089 3464 5120
rect 3881 5117 3893 5120
rect 3927 5148 3939 5151
rect 3970 5148 3976 5160
rect 3927 5120 3976 5148
rect 3927 5117 3939 5120
rect 3881 5111 3939 5117
rect 3970 5108 3976 5120
rect 4028 5108 4034 5160
rect 4982 5148 4988 5160
rect 4448 5120 4988 5148
rect 2317 5083 2375 5089
rect 2317 5049 2329 5083
rect 2363 5080 2375 5083
rect 3421 5083 3479 5089
rect 3421 5080 3433 5083
rect 2363 5052 3433 5080
rect 2363 5049 2375 5052
rect 2317 5043 2375 5049
rect 3421 5049 3433 5052
rect 3467 5049 3479 5083
rect 3421 5043 3479 5049
rect 3605 5083 3663 5089
rect 3605 5049 3617 5083
rect 3651 5080 3663 5083
rect 4448 5080 4476 5120
rect 4982 5108 4988 5120
rect 5040 5108 5046 5160
rect 5258 5108 5264 5160
rect 5316 5108 5322 5160
rect 5350 5108 5356 5160
rect 5408 5108 5414 5160
rect 5442 5108 5448 5160
rect 5500 5108 5506 5160
rect 5534 5108 5540 5160
rect 5592 5148 5598 5160
rect 5902 5148 5908 5160
rect 5592 5120 5908 5148
rect 5592 5108 5598 5120
rect 5902 5108 5908 5120
rect 5960 5108 5966 5160
rect 6181 5151 6239 5157
rect 6181 5117 6193 5151
rect 6227 5148 6239 5151
rect 6227 5120 6592 5148
rect 6227 5117 6239 5120
rect 6181 5111 6239 5117
rect 3651 5052 4476 5080
rect 4801 5083 4859 5089
rect 3651 5049 3663 5052
rect 3605 5043 3663 5049
rect 4801 5049 4813 5083
rect 4847 5049 4859 5083
rect 5368 5080 5396 5108
rect 5368 5052 5488 5080
rect 4801 5043 4859 5049
rect 1302 4972 1308 5024
rect 1360 4972 1366 5024
rect 1670 4972 1676 5024
rect 1728 5012 1734 5024
rect 2685 5015 2743 5021
rect 2685 5012 2697 5015
rect 1728 4984 2697 5012
rect 1728 4972 1734 4984
rect 2685 4981 2697 4984
rect 2731 4981 2743 5015
rect 2685 4975 2743 4981
rect 3510 4972 3516 5024
rect 3568 5012 3574 5024
rect 4816 5012 4844 5043
rect 4890 5012 4896 5024
rect 3568 4984 4896 5012
rect 3568 4972 3574 4984
rect 4890 4972 4896 4984
rect 4948 4972 4954 5024
rect 5166 4972 5172 5024
rect 5224 4972 5230 5024
rect 5350 4972 5356 5024
rect 5408 4972 5414 5024
rect 5460 5012 5488 5052
rect 5626 5040 5632 5092
rect 5684 5080 5690 5092
rect 6454 5080 6460 5092
rect 5684 5052 6460 5080
rect 5684 5040 5690 5052
rect 6454 5040 6460 5052
rect 6512 5040 6518 5092
rect 5534 5012 5540 5024
rect 5460 4984 5540 5012
rect 5534 4972 5540 4984
rect 5592 4972 5598 5024
rect 6089 5015 6147 5021
rect 6089 4981 6101 5015
rect 6135 5012 6147 5015
rect 6178 5012 6184 5024
rect 6135 4984 6184 5012
rect 6135 4981 6147 4984
rect 6089 4975 6147 4981
rect 6178 4972 6184 4984
rect 6236 4972 6242 5024
rect 6564 5012 6592 5120
rect 6638 5108 6644 5160
rect 6696 5108 6702 5160
rect 6733 5151 6791 5157
rect 6733 5117 6745 5151
rect 6779 5117 6791 5151
rect 6733 5111 6791 5117
rect 6748 5080 6776 5111
rect 6914 5108 6920 5160
rect 6972 5108 6978 5160
rect 7006 5108 7012 5160
rect 7064 5108 7070 5160
rect 7116 5157 7144 5188
rect 7377 5185 7389 5219
rect 7423 5216 7435 5219
rect 8570 5216 8576 5228
rect 7423 5188 8576 5216
rect 7423 5185 7435 5188
rect 7377 5179 7435 5185
rect 8570 5176 8576 5188
rect 8628 5176 8634 5228
rect 9048 5216 9076 5256
rect 10134 5244 10140 5256
rect 10192 5244 10198 5296
rect 11992 5284 12020 5324
rect 12437 5321 12449 5324
rect 12483 5321 12495 5355
rect 12437 5315 12495 5321
rect 12710 5312 12716 5364
rect 12768 5352 12774 5364
rect 12805 5355 12863 5361
rect 12805 5352 12817 5355
rect 12768 5324 12817 5352
rect 12768 5312 12774 5324
rect 12805 5321 12817 5324
rect 12851 5321 12863 5355
rect 12805 5315 12863 5321
rect 12986 5312 12992 5364
rect 13044 5352 13050 5364
rect 17037 5355 17095 5361
rect 13044 5324 16896 5352
rect 13044 5312 13050 5324
rect 11532 5256 12020 5284
rect 8956 5188 9076 5216
rect 7101 5151 7159 5157
rect 7101 5117 7113 5151
rect 7147 5117 7159 5151
rect 7101 5111 7159 5117
rect 7561 5151 7619 5157
rect 7561 5117 7573 5151
rect 7607 5148 7619 5151
rect 7650 5148 7656 5160
rect 7607 5120 7656 5148
rect 7607 5117 7619 5120
rect 7561 5111 7619 5117
rect 7650 5108 7656 5120
rect 7708 5108 7714 5160
rect 7745 5151 7803 5157
rect 7745 5117 7757 5151
rect 7791 5117 7803 5151
rect 7745 5111 7803 5117
rect 7837 5151 7895 5157
rect 7837 5117 7849 5151
rect 7883 5117 7895 5151
rect 7837 5111 7895 5117
rect 7929 5151 7987 5157
rect 7929 5117 7941 5151
rect 7975 5148 7987 5151
rect 8754 5148 8760 5160
rect 7975 5120 8760 5148
rect 7975 5117 7987 5120
rect 7929 5111 7987 5117
rect 7190 5080 7196 5092
rect 6748 5052 7196 5080
rect 7190 5040 7196 5052
rect 7248 5040 7254 5092
rect 6914 5012 6920 5024
rect 6564 4984 6920 5012
rect 6914 4972 6920 4984
rect 6972 4972 6978 5024
rect 7760 5012 7788 5111
rect 7852 5080 7880 5111
rect 8754 5108 8760 5120
rect 8812 5148 8818 5160
rect 8956 5148 8984 5188
rect 9122 5176 9128 5228
rect 9180 5176 9186 5228
rect 9769 5219 9827 5225
rect 9769 5185 9781 5219
rect 9815 5216 9827 5219
rect 10042 5216 10048 5228
rect 9815 5188 10048 5216
rect 9815 5185 9827 5188
rect 9769 5179 9827 5185
rect 10042 5176 10048 5188
rect 10100 5176 10106 5228
rect 10965 5219 11023 5225
rect 10965 5185 10977 5219
rect 11011 5216 11023 5219
rect 11054 5216 11060 5228
rect 11011 5188 11060 5216
rect 11011 5185 11023 5188
rect 10965 5179 11023 5185
rect 11054 5176 11060 5188
rect 11112 5176 11118 5228
rect 11532 5216 11560 5256
rect 12894 5244 12900 5296
rect 12952 5284 12958 5296
rect 16868 5284 16896 5324
rect 17037 5321 17049 5355
rect 17083 5352 17095 5355
rect 19058 5352 19064 5364
rect 17083 5324 19064 5352
rect 17083 5321 17095 5324
rect 17037 5315 17095 5321
rect 19058 5312 19064 5324
rect 19116 5312 19122 5364
rect 19613 5355 19671 5361
rect 19613 5321 19625 5355
rect 19659 5352 19671 5355
rect 19794 5352 19800 5364
rect 19659 5324 19800 5352
rect 19659 5321 19671 5324
rect 19613 5315 19671 5321
rect 19794 5312 19800 5324
rect 19852 5312 19858 5364
rect 20162 5312 20168 5364
rect 20220 5352 20226 5364
rect 20441 5355 20499 5361
rect 20441 5352 20453 5355
rect 20220 5324 20453 5352
rect 20220 5312 20226 5324
rect 20441 5321 20453 5324
rect 20487 5321 20499 5355
rect 20441 5315 20499 5321
rect 20533 5355 20591 5361
rect 20533 5321 20545 5355
rect 20579 5352 20591 5355
rect 20714 5352 20720 5364
rect 20579 5324 20720 5352
rect 20579 5321 20591 5324
rect 20533 5315 20591 5321
rect 20714 5312 20720 5324
rect 20772 5352 20778 5364
rect 21450 5352 21456 5364
rect 20772 5324 21456 5352
rect 20772 5312 20778 5324
rect 21450 5312 21456 5324
rect 21508 5312 21514 5364
rect 21821 5355 21879 5361
rect 21821 5321 21833 5355
rect 21867 5352 21879 5355
rect 22002 5352 22008 5364
rect 21867 5324 22008 5352
rect 21867 5321 21879 5324
rect 21821 5315 21879 5321
rect 22002 5312 22008 5324
rect 22060 5312 22066 5364
rect 20254 5284 20260 5296
rect 12952 5256 16804 5284
rect 16868 5256 20260 5284
rect 12952 5244 12958 5256
rect 12986 5216 12992 5228
rect 11164 5188 11560 5216
rect 8812 5120 8984 5148
rect 9033 5151 9091 5157
rect 8812 5108 8818 5120
rect 9033 5117 9045 5151
rect 9079 5148 9091 5151
rect 9214 5148 9220 5160
rect 9079 5120 9220 5148
rect 9079 5117 9091 5120
rect 9033 5111 9091 5117
rect 9214 5108 9220 5120
rect 9272 5148 9278 5160
rect 10781 5151 10839 5157
rect 10781 5148 10793 5151
rect 9272 5120 10793 5148
rect 9272 5108 9278 5120
rect 10781 5117 10793 5120
rect 10827 5148 10839 5151
rect 11164 5148 11192 5188
rect 10827 5120 11192 5148
rect 10827 5117 10839 5120
rect 10781 5111 10839 5117
rect 11238 5108 11244 5160
rect 11296 5108 11302 5160
rect 11330 5108 11336 5160
rect 11388 5108 11394 5160
rect 11532 5157 11560 5188
rect 12728 5188 12992 5216
rect 11517 5151 11575 5157
rect 11517 5117 11529 5151
rect 11563 5117 11575 5151
rect 11517 5111 11575 5117
rect 11609 5151 11667 5157
rect 11609 5117 11621 5151
rect 11655 5148 11667 5151
rect 11790 5148 11796 5160
rect 11655 5120 11796 5148
rect 11655 5117 11667 5120
rect 11609 5111 11667 5117
rect 11790 5108 11796 5120
rect 11848 5108 11854 5160
rect 12069 5151 12127 5157
rect 12069 5117 12081 5151
rect 12115 5148 12127 5151
rect 12158 5148 12164 5160
rect 12115 5120 12164 5148
rect 12115 5117 12127 5120
rect 12069 5111 12127 5117
rect 12158 5108 12164 5120
rect 12216 5108 12222 5160
rect 12728 5157 12756 5188
rect 12986 5176 12992 5188
rect 13044 5176 13050 5228
rect 14090 5176 14096 5228
rect 14148 5176 14154 5228
rect 14458 5176 14464 5228
rect 14516 5216 14522 5228
rect 15565 5219 15623 5225
rect 14516 5188 14964 5216
rect 14516 5176 14522 5188
rect 12345 5151 12403 5157
rect 12345 5117 12357 5151
rect 12391 5148 12403 5151
rect 12621 5151 12679 5157
rect 12621 5148 12633 5151
rect 12391 5120 12633 5148
rect 12391 5117 12403 5120
rect 12345 5111 12403 5117
rect 12621 5117 12633 5120
rect 12667 5117 12679 5151
rect 12621 5111 12679 5117
rect 12713 5151 12771 5157
rect 12713 5117 12725 5151
rect 12759 5117 12771 5151
rect 12713 5111 12771 5117
rect 12897 5151 12955 5157
rect 12897 5117 12909 5151
rect 12943 5148 12955 5151
rect 13262 5148 13268 5160
rect 12943 5120 13268 5148
rect 12943 5117 12955 5120
rect 12897 5111 12955 5117
rect 8110 5080 8116 5092
rect 7852 5052 8116 5080
rect 8110 5040 8116 5052
rect 8168 5040 8174 5092
rect 8941 5083 8999 5089
rect 8941 5049 8953 5083
rect 8987 5080 8999 5083
rect 9306 5080 9312 5092
rect 8987 5052 9312 5080
rect 8987 5049 8999 5052
rect 8941 5043 8999 5049
rect 9306 5040 9312 5052
rect 9364 5040 9370 5092
rect 9861 5083 9919 5089
rect 9861 5049 9873 5083
rect 9907 5080 9919 5083
rect 10134 5080 10140 5092
rect 9907 5052 10140 5080
rect 9907 5049 9919 5052
rect 9861 5043 9919 5049
rect 10134 5040 10140 5052
rect 10192 5080 10198 5092
rect 10873 5083 10931 5089
rect 10873 5080 10885 5083
rect 10192 5052 10885 5080
rect 10192 5040 10198 5052
rect 10873 5049 10885 5052
rect 10919 5080 10931 5083
rect 12636 5080 12664 5111
rect 13262 5108 13268 5120
rect 13320 5108 13326 5160
rect 13814 5108 13820 5160
rect 13872 5148 13878 5160
rect 13998 5148 14004 5160
rect 13872 5120 14004 5148
rect 13872 5108 13878 5120
rect 13998 5108 14004 5120
rect 14056 5108 14062 5160
rect 14182 5108 14188 5160
rect 14240 5148 14246 5160
rect 14553 5151 14611 5157
rect 14553 5148 14565 5151
rect 14240 5120 14565 5148
rect 14240 5108 14246 5120
rect 14553 5117 14565 5120
rect 14599 5148 14611 5151
rect 14734 5148 14740 5160
rect 14599 5120 14740 5148
rect 14599 5117 14611 5120
rect 14553 5111 14611 5117
rect 14734 5108 14740 5120
rect 14792 5148 14798 5160
rect 14829 5151 14887 5157
rect 14829 5148 14841 5151
rect 14792 5120 14841 5148
rect 14792 5108 14798 5120
rect 14829 5117 14841 5120
rect 14875 5117 14887 5151
rect 14936 5148 14964 5188
rect 15565 5185 15577 5219
rect 15611 5216 15623 5219
rect 16574 5216 16580 5228
rect 15611 5188 16580 5216
rect 15611 5185 15623 5188
rect 15565 5179 15623 5185
rect 16574 5176 16580 5188
rect 16632 5176 16638 5228
rect 16666 5176 16672 5228
rect 16724 5176 16730 5228
rect 16776 5225 16804 5256
rect 20254 5244 20260 5256
rect 20312 5284 20318 5296
rect 20312 5256 21956 5284
rect 20312 5244 20318 5256
rect 16761 5219 16819 5225
rect 16761 5185 16773 5219
rect 16807 5185 16819 5219
rect 16761 5179 16819 5185
rect 15749 5151 15807 5157
rect 15749 5148 15761 5151
rect 14936 5120 15761 5148
rect 14829 5111 14887 5117
rect 15749 5117 15761 5120
rect 15795 5117 15807 5151
rect 15749 5111 15807 5117
rect 16485 5151 16543 5157
rect 16485 5117 16497 5151
rect 16531 5117 16543 5151
rect 16776 5148 16804 5179
rect 17034 5176 17040 5228
rect 17092 5216 17098 5228
rect 17497 5219 17555 5225
rect 17497 5216 17509 5219
rect 17092 5188 17509 5216
rect 17092 5176 17098 5188
rect 17497 5185 17509 5188
rect 17543 5185 17555 5219
rect 17497 5179 17555 5185
rect 19058 5176 19064 5228
rect 19116 5176 19122 5228
rect 19978 5216 19984 5228
rect 19536 5188 19984 5216
rect 17221 5151 17279 5157
rect 17221 5148 17233 5151
rect 16776 5120 17233 5148
rect 16485 5111 16543 5117
rect 17221 5117 17233 5120
rect 17267 5117 17279 5151
rect 17221 5111 17279 5117
rect 10919 5052 12434 5080
rect 12636 5052 14688 5080
rect 10919 5049 10931 5052
rect 10873 5043 10931 5049
rect 7926 5012 7932 5024
rect 7760 4984 7932 5012
rect 7926 4972 7932 4984
rect 7984 4972 7990 5024
rect 9766 4972 9772 5024
rect 9824 5012 9830 5024
rect 9953 5015 10011 5021
rect 9953 5012 9965 5015
rect 9824 4984 9965 5012
rect 9824 4972 9830 4984
rect 9953 4981 9965 4984
rect 9999 5012 10011 5015
rect 12161 5015 12219 5021
rect 12161 5012 12173 5015
rect 9999 4984 12173 5012
rect 9999 4981 10011 4984
rect 9953 4975 10011 4981
rect 12161 4981 12173 4984
rect 12207 5012 12219 5015
rect 12250 5012 12256 5024
rect 12207 4984 12256 5012
rect 12207 4981 12219 4984
rect 12161 4975 12219 4981
rect 12250 4972 12256 4984
rect 12308 4972 12314 5024
rect 12406 5012 12434 5052
rect 14660 5024 14688 5052
rect 16022 5040 16028 5092
rect 16080 5080 16086 5092
rect 16301 5083 16359 5089
rect 16301 5080 16313 5083
rect 16080 5052 16313 5080
rect 16080 5040 16086 5052
rect 16301 5049 16313 5052
rect 16347 5049 16359 5083
rect 16500 5080 16528 5111
rect 17402 5108 17408 5160
rect 17460 5108 17466 5160
rect 17586 5108 17592 5160
rect 17644 5108 17650 5160
rect 17773 5151 17831 5157
rect 17773 5117 17785 5151
rect 17819 5117 17831 5151
rect 17773 5111 17831 5117
rect 17788 5080 17816 5111
rect 18690 5108 18696 5160
rect 18748 5148 18754 5160
rect 18785 5151 18843 5157
rect 18785 5148 18797 5151
rect 18748 5120 18797 5148
rect 18748 5108 18754 5120
rect 18785 5117 18797 5120
rect 18831 5117 18843 5151
rect 18785 5111 18843 5117
rect 18877 5151 18935 5157
rect 18877 5117 18889 5151
rect 18923 5117 18935 5151
rect 18877 5111 18935 5117
rect 17862 5080 17868 5092
rect 16500 5052 17868 5080
rect 16301 5043 16359 5049
rect 17862 5040 17868 5052
rect 17920 5040 17926 5092
rect 12710 5012 12716 5024
rect 12406 4984 12716 5012
rect 12710 4972 12716 4984
rect 12768 4972 12774 5024
rect 12986 4972 12992 5024
rect 13044 5012 13050 5024
rect 13541 5015 13599 5021
rect 13541 5012 13553 5015
rect 13044 4984 13553 5012
rect 13044 4972 13050 4984
rect 13541 4981 13553 4984
rect 13587 4981 13599 5015
rect 13541 4975 13599 4981
rect 13909 5015 13967 5021
rect 13909 4981 13921 5015
rect 13955 5012 13967 5015
rect 14366 5012 14372 5024
rect 13955 4984 14372 5012
rect 13955 4981 13967 4984
rect 13909 4975 13967 4981
rect 14366 4972 14372 4984
rect 14424 4972 14430 5024
rect 14642 4972 14648 5024
rect 14700 5012 14706 5024
rect 15657 5015 15715 5021
rect 15657 5012 15669 5015
rect 14700 4984 15669 5012
rect 14700 4972 14706 4984
rect 15657 4981 15669 4984
rect 15703 4981 15715 5015
rect 15657 4975 15715 4981
rect 16117 5015 16175 5021
rect 16117 4981 16129 5015
rect 16163 5012 16175 5015
rect 16206 5012 16212 5024
rect 16163 4984 16212 5012
rect 16163 4981 16175 4984
rect 16117 4975 16175 4981
rect 16206 4972 16212 4984
rect 16264 4972 16270 5024
rect 18230 4972 18236 5024
rect 18288 5012 18294 5024
rect 18892 5012 18920 5111
rect 18966 5108 18972 5160
rect 19024 5108 19030 5160
rect 19536 5157 19564 5188
rect 19978 5176 19984 5188
rect 20036 5176 20042 5228
rect 21928 5225 21956 5256
rect 21913 5219 21971 5225
rect 21913 5185 21925 5219
rect 21959 5216 21971 5219
rect 22278 5216 22284 5228
rect 21959 5188 22284 5216
rect 21959 5185 21971 5188
rect 21913 5179 21971 5185
rect 22278 5176 22284 5188
rect 22336 5176 22342 5228
rect 19521 5151 19579 5157
rect 19521 5117 19533 5151
rect 19567 5117 19579 5151
rect 19521 5111 19579 5117
rect 19797 5151 19855 5157
rect 19797 5117 19809 5151
rect 19843 5117 19855 5151
rect 19797 5111 19855 5117
rect 19058 5040 19064 5092
rect 19116 5080 19122 5092
rect 19812 5080 19840 5111
rect 19886 5108 19892 5160
rect 19944 5148 19950 5160
rect 20257 5151 20315 5157
rect 20257 5148 20269 5151
rect 19944 5120 20269 5148
rect 19944 5108 19950 5120
rect 20257 5117 20269 5120
rect 20303 5117 20315 5151
rect 20257 5111 20315 5117
rect 20717 5151 20775 5157
rect 20717 5117 20729 5151
rect 20763 5148 20775 5151
rect 21082 5148 21088 5160
rect 20763 5120 21088 5148
rect 20763 5117 20775 5120
rect 20717 5111 20775 5117
rect 21082 5108 21088 5120
rect 21140 5108 21146 5160
rect 21174 5108 21180 5160
rect 21232 5108 21238 5160
rect 21542 5108 21548 5160
rect 21600 5108 21606 5160
rect 20073 5083 20131 5089
rect 20073 5080 20085 5083
rect 19116 5052 19380 5080
rect 19812 5052 20085 5080
rect 19116 5040 19122 5052
rect 18288 4984 18920 5012
rect 18288 4972 18294 4984
rect 19150 4972 19156 5024
rect 19208 5012 19214 5024
rect 19352 5021 19380 5052
rect 20073 5049 20085 5052
rect 20119 5080 20131 5083
rect 20901 5083 20959 5089
rect 20119 5052 20668 5080
rect 20119 5049 20131 5052
rect 20073 5043 20131 5049
rect 20640 5024 20668 5052
rect 20901 5049 20913 5083
rect 20947 5049 20959 5083
rect 20901 5043 20959 5049
rect 19245 5015 19303 5021
rect 19245 5012 19257 5015
rect 19208 4984 19257 5012
rect 19208 4972 19214 4984
rect 19245 4981 19257 4984
rect 19291 4981 19303 5015
rect 19245 4975 19303 4981
rect 19337 5015 19395 5021
rect 19337 4981 19349 5015
rect 19383 4981 19395 5015
rect 19337 4975 19395 4981
rect 19702 4972 19708 5024
rect 19760 5012 19766 5024
rect 19978 5012 19984 5024
rect 19760 4984 19984 5012
rect 19760 4972 19766 4984
rect 19978 4972 19984 4984
rect 20036 4972 20042 5024
rect 20622 4972 20628 5024
rect 20680 5012 20686 5024
rect 20916 5012 20944 5043
rect 21358 5040 21364 5092
rect 21416 5080 21422 5092
rect 21637 5083 21695 5089
rect 21637 5080 21649 5083
rect 21416 5052 21649 5080
rect 21416 5040 21422 5052
rect 21637 5049 21649 5052
rect 21683 5049 21695 5083
rect 21637 5043 21695 5049
rect 21726 5040 21732 5092
rect 21784 5080 21790 5092
rect 22005 5083 22063 5089
rect 22005 5080 22017 5083
rect 21784 5052 22017 5080
rect 21784 5040 21790 5052
rect 22005 5049 22017 5052
rect 22051 5049 22063 5083
rect 22005 5043 22063 5049
rect 20993 5015 21051 5021
rect 20993 5012 21005 5015
rect 20680 4984 21005 5012
rect 20680 4972 20686 4984
rect 20993 4981 21005 4984
rect 21039 4981 21051 5015
rect 20993 4975 21051 4981
rect 552 4922 23368 4944
rect 552 4870 4366 4922
rect 4418 4870 4430 4922
rect 4482 4870 4494 4922
rect 4546 4870 4558 4922
rect 4610 4870 4622 4922
rect 4674 4870 4686 4922
rect 4738 4870 10366 4922
rect 10418 4870 10430 4922
rect 10482 4870 10494 4922
rect 10546 4870 10558 4922
rect 10610 4870 10622 4922
rect 10674 4870 10686 4922
rect 10738 4870 16366 4922
rect 16418 4870 16430 4922
rect 16482 4870 16494 4922
rect 16546 4870 16558 4922
rect 16610 4870 16622 4922
rect 16674 4870 16686 4922
rect 16738 4870 22366 4922
rect 22418 4870 22430 4922
rect 22482 4870 22494 4922
rect 22546 4870 22558 4922
rect 22610 4870 22622 4922
rect 22674 4870 22686 4922
rect 22738 4870 23368 4922
rect 552 4848 23368 4870
rect 1118 4768 1124 4820
rect 1176 4768 1182 4820
rect 2314 4808 2320 4820
rect 2148 4780 2320 4808
rect 1486 4740 1492 4752
rect 1044 4712 1492 4740
rect 658 4632 664 4684
rect 716 4672 722 4684
rect 1044 4681 1072 4712
rect 1486 4700 1492 4712
rect 1544 4700 1550 4752
rect 2148 4740 2176 4780
rect 2314 4768 2320 4780
rect 2372 4768 2378 4820
rect 2409 4811 2467 4817
rect 2409 4777 2421 4811
rect 2455 4808 2467 4811
rect 2682 4808 2688 4820
rect 2455 4780 2688 4808
rect 2455 4777 2467 4780
rect 2409 4771 2467 4777
rect 2682 4768 2688 4780
rect 2740 4768 2746 4820
rect 2774 4768 2780 4820
rect 2832 4808 2838 4820
rect 3234 4808 3240 4820
rect 2832 4780 3240 4808
rect 2832 4768 2838 4780
rect 3234 4768 3240 4780
rect 3292 4768 3298 4820
rect 3421 4811 3479 4817
rect 3421 4777 3433 4811
rect 3467 4808 3479 4811
rect 3510 4808 3516 4820
rect 3467 4780 3516 4808
rect 3467 4777 3479 4780
rect 3421 4771 3479 4777
rect 3510 4768 3516 4780
rect 3568 4768 3574 4820
rect 3786 4768 3792 4820
rect 3844 4808 3850 4820
rect 3881 4811 3939 4817
rect 3881 4808 3893 4811
rect 3844 4780 3893 4808
rect 3844 4768 3850 4780
rect 3881 4777 3893 4780
rect 3927 4777 3939 4811
rect 3881 4771 3939 4777
rect 4341 4811 4399 4817
rect 4341 4777 4353 4811
rect 4387 4808 4399 4811
rect 4798 4808 4804 4820
rect 4387 4780 4804 4808
rect 4387 4777 4399 4780
rect 4341 4771 4399 4777
rect 2056 4712 2176 4740
rect 2056 4684 2084 4712
rect 2222 4700 2228 4752
rect 2280 4740 2286 4752
rect 3145 4743 3203 4749
rect 3145 4740 3157 4743
rect 2280 4712 3157 4740
rect 2280 4700 2286 4712
rect 3145 4709 3157 4712
rect 3191 4709 3203 4743
rect 3896 4740 3924 4771
rect 4798 4768 4804 4780
rect 4856 4768 4862 4820
rect 4985 4811 5043 4817
rect 4985 4777 4997 4811
rect 5031 4808 5043 4811
rect 5258 4808 5264 4820
rect 5031 4780 5264 4808
rect 5031 4777 5043 4780
rect 4985 4771 5043 4777
rect 5258 4768 5264 4780
rect 5316 4768 5322 4820
rect 5626 4768 5632 4820
rect 5684 4768 5690 4820
rect 6733 4811 6791 4817
rect 6733 4777 6745 4811
rect 6779 4808 6791 4811
rect 7006 4808 7012 4820
rect 6779 4780 7012 4808
rect 6779 4777 6791 4780
rect 6733 4771 6791 4777
rect 7006 4768 7012 4780
rect 7064 4768 7070 4820
rect 9214 4768 9220 4820
rect 9272 4768 9278 4820
rect 9309 4811 9367 4817
rect 9309 4777 9321 4811
rect 9355 4808 9367 4811
rect 10134 4808 10140 4820
rect 9355 4780 10140 4808
rect 9355 4777 9367 4780
rect 9309 4771 9367 4777
rect 10134 4768 10140 4780
rect 10192 4768 10198 4820
rect 12250 4808 12256 4820
rect 10244 4780 12256 4808
rect 4522 4740 4528 4752
rect 3896 4712 4528 4740
rect 3145 4703 3203 4709
rect 4522 4700 4528 4712
rect 4580 4700 4586 4752
rect 4617 4743 4675 4749
rect 4617 4709 4629 4743
rect 4663 4740 4675 4743
rect 4890 4740 4896 4752
rect 4663 4712 4896 4740
rect 4663 4709 4675 4712
rect 4617 4703 4675 4709
rect 4890 4700 4896 4712
rect 4948 4700 4954 4752
rect 5718 4740 5724 4752
rect 5000 4712 5724 4740
rect 845 4675 903 4681
rect 845 4672 857 4675
rect 716 4644 857 4672
rect 716 4632 722 4644
rect 845 4641 857 4644
rect 891 4641 903 4675
rect 845 4635 903 4641
rect 1029 4675 1087 4681
rect 1029 4641 1041 4675
rect 1075 4641 1087 4675
rect 1029 4635 1087 4641
rect 860 4536 888 4635
rect 1302 4632 1308 4684
rect 1360 4632 1366 4684
rect 1397 4675 1455 4681
rect 1397 4641 1409 4675
rect 1443 4672 1455 4675
rect 1443 4644 1808 4672
rect 1443 4641 1455 4644
rect 1397 4635 1455 4641
rect 937 4607 995 4613
rect 937 4573 949 4607
rect 983 4604 995 4607
rect 1118 4604 1124 4616
rect 983 4576 1124 4604
rect 983 4573 995 4576
rect 937 4567 995 4573
rect 1118 4564 1124 4576
rect 1176 4564 1182 4616
rect 1780 4548 1808 4644
rect 1854 4632 1860 4684
rect 1912 4632 1918 4684
rect 2038 4632 2044 4684
rect 2096 4632 2102 4684
rect 2133 4675 2191 4681
rect 2133 4641 2145 4675
rect 2179 4641 2191 4675
rect 2133 4635 2191 4641
rect 2148 4604 2176 4635
rect 2314 4632 2320 4684
rect 2372 4672 2378 4684
rect 2593 4675 2651 4681
rect 2593 4672 2605 4675
rect 2372 4644 2605 4672
rect 2372 4632 2378 4644
rect 2593 4641 2605 4644
rect 2639 4641 2651 4675
rect 2593 4635 2651 4641
rect 2869 4675 2927 4681
rect 2869 4641 2881 4675
rect 2915 4672 2927 4675
rect 2958 4672 2964 4684
rect 2915 4644 2964 4672
rect 2915 4641 2927 4644
rect 2869 4635 2927 4641
rect 2958 4632 2964 4644
rect 3016 4632 3022 4684
rect 3329 4675 3387 4681
rect 3329 4641 3341 4675
rect 3375 4641 3387 4675
rect 3329 4635 3387 4641
rect 3605 4675 3663 4681
rect 3605 4641 3617 4675
rect 3651 4672 3663 4675
rect 3694 4672 3700 4684
rect 3651 4644 3700 4672
rect 3651 4641 3663 4644
rect 3605 4635 3663 4641
rect 3344 4604 3372 4635
rect 3694 4632 3700 4644
rect 3752 4632 3758 4684
rect 4062 4632 4068 4684
rect 4120 4632 4126 4684
rect 4154 4632 4160 4684
rect 4212 4632 4218 4684
rect 4801 4675 4859 4681
rect 4801 4641 4813 4675
rect 4847 4672 4859 4675
rect 5000 4672 5028 4712
rect 5718 4700 5724 4712
rect 5776 4700 5782 4752
rect 7190 4700 7196 4752
rect 7248 4740 7254 4752
rect 7529 4743 7587 4749
rect 7529 4740 7541 4743
rect 7248 4712 7541 4740
rect 7248 4700 7254 4712
rect 7529 4709 7541 4712
rect 7575 4709 7587 4743
rect 7529 4703 7587 4709
rect 7650 4700 7656 4752
rect 7708 4740 7714 4752
rect 7745 4743 7803 4749
rect 7745 4740 7757 4743
rect 7708 4712 7757 4740
rect 7708 4700 7714 4712
rect 7745 4709 7757 4712
rect 7791 4709 7803 4743
rect 7745 4703 7803 4709
rect 9766 4700 9772 4752
rect 9824 4740 9830 4752
rect 10045 4743 10103 4749
rect 10045 4740 10057 4743
rect 9824 4712 10057 4740
rect 9824 4700 9830 4712
rect 10045 4709 10057 4712
rect 10091 4709 10103 4743
rect 10045 4703 10103 4709
rect 4847 4644 5028 4672
rect 5261 4675 5319 4681
rect 4847 4641 4859 4644
rect 4801 4635 4859 4641
rect 4908 4616 4936 4644
rect 5261 4641 5273 4675
rect 5307 4672 5319 4675
rect 5813 4675 5871 4681
rect 5813 4672 5825 4675
rect 5307 4644 5825 4672
rect 5307 4641 5319 4644
rect 5261 4635 5319 4641
rect 5813 4641 5825 4644
rect 5859 4641 5871 4675
rect 5813 4635 5871 4641
rect 2148 4576 3372 4604
rect 1673 4539 1731 4545
rect 1673 4536 1685 4539
rect 860 4508 1685 4536
rect 1673 4505 1685 4508
rect 1719 4505 1731 4539
rect 1673 4499 1731 4505
rect 1762 4496 1768 4548
rect 1820 4536 1826 4548
rect 2590 4536 2596 4548
rect 1820 4508 2596 4536
rect 1820 4496 1826 4508
rect 2590 4496 2596 4508
rect 2648 4496 2654 4548
rect 3344 4536 3372 4576
rect 4246 4564 4252 4616
rect 4304 4604 4310 4616
rect 4341 4607 4399 4613
rect 4341 4604 4353 4607
rect 4304 4576 4353 4604
rect 4304 4564 4310 4576
rect 4341 4573 4353 4576
rect 4387 4573 4399 4607
rect 4341 4567 4399 4573
rect 4890 4564 4896 4616
rect 4948 4564 4954 4616
rect 4982 4536 4988 4548
rect 3344 4508 4988 4536
rect 4982 4496 4988 4508
rect 5040 4536 5046 4548
rect 5276 4536 5304 4635
rect 6178 4632 6184 4684
rect 6236 4672 6242 4684
rect 7101 4675 7159 4681
rect 7101 4672 7113 4675
rect 6236 4644 7113 4672
rect 6236 4632 6242 4644
rect 7101 4641 7113 4644
rect 7147 4641 7159 4675
rect 7101 4635 7159 4641
rect 8205 4675 8263 4681
rect 8205 4641 8217 4675
rect 8251 4672 8263 4675
rect 8386 4672 8392 4684
rect 8251 4644 8392 4672
rect 8251 4641 8263 4644
rect 8205 4635 8263 4641
rect 8386 4632 8392 4644
rect 8444 4632 8450 4684
rect 8570 4632 8576 4684
rect 8628 4672 8634 4684
rect 10244 4672 10272 4780
rect 12250 4768 12256 4780
rect 12308 4768 12314 4820
rect 12452 4780 13952 4808
rect 12452 4740 12480 4780
rect 12268 4712 12480 4740
rect 12529 4743 12587 4749
rect 8628 4644 10272 4672
rect 8628 4632 8634 4644
rect 11514 4632 11520 4684
rect 11572 4672 11578 4684
rect 11793 4675 11851 4681
rect 11793 4672 11805 4675
rect 11572 4644 11805 4672
rect 11572 4632 11578 4644
rect 11793 4641 11805 4644
rect 11839 4641 11851 4675
rect 11793 4635 11851 4641
rect 11882 4632 11888 4684
rect 11940 4672 11946 4684
rect 12268 4681 12296 4712
rect 12529 4709 12541 4743
rect 12575 4740 12587 4743
rect 12618 4740 12624 4752
rect 12575 4712 12624 4740
rect 12575 4709 12587 4712
rect 12529 4703 12587 4709
rect 12618 4700 12624 4712
rect 12676 4700 12682 4752
rect 13924 4740 13952 4780
rect 13998 4768 14004 4820
rect 14056 4808 14062 4820
rect 14458 4808 14464 4820
rect 14056 4780 14464 4808
rect 14056 4768 14062 4780
rect 14458 4768 14464 4780
rect 14516 4768 14522 4820
rect 14553 4811 14611 4817
rect 14553 4777 14565 4811
rect 14599 4808 14611 4811
rect 14642 4808 14648 4820
rect 14599 4780 14648 4808
rect 14599 4777 14611 4780
rect 14553 4771 14611 4777
rect 14642 4768 14648 4780
rect 14700 4768 14706 4820
rect 17862 4768 17868 4820
rect 17920 4808 17926 4820
rect 18325 4811 18383 4817
rect 17920 4780 18276 4808
rect 17920 4768 17926 4780
rect 15470 4740 15476 4752
rect 12728 4712 13584 4740
rect 13924 4712 15476 4740
rect 12069 4675 12127 4681
rect 12069 4672 12081 4675
rect 11940 4644 12081 4672
rect 11940 4632 11946 4644
rect 12069 4641 12081 4644
rect 12115 4641 12127 4675
rect 12069 4635 12127 4641
rect 12253 4675 12311 4681
rect 12253 4641 12265 4675
rect 12299 4641 12311 4675
rect 12253 4635 12311 4641
rect 12345 4675 12403 4681
rect 12345 4641 12357 4675
rect 12391 4672 12403 4675
rect 12728 4672 12756 4712
rect 12391 4644 12756 4672
rect 12391 4641 12403 4644
rect 12345 4635 12403 4641
rect 5350 4564 5356 4616
rect 5408 4564 5414 4616
rect 6089 4607 6147 4613
rect 6089 4604 6101 4607
rect 5552 4576 6101 4604
rect 5040 4508 5304 4536
rect 5040 4496 5046 4508
rect 2958 4428 2964 4480
rect 3016 4428 3022 4480
rect 5258 4428 5264 4480
rect 5316 4468 5322 4480
rect 5552 4468 5580 4576
rect 6089 4573 6101 4576
rect 6135 4604 6147 4607
rect 6730 4604 6736 4616
rect 6135 4576 6736 4604
rect 6135 4573 6147 4576
rect 6089 4567 6147 4573
rect 6730 4564 6736 4576
rect 6788 4564 6794 4616
rect 6917 4607 6975 4613
rect 6917 4573 6929 4607
rect 6963 4573 6975 4607
rect 6917 4567 6975 4573
rect 5902 4496 5908 4548
rect 5960 4536 5966 4548
rect 6932 4536 6960 4567
rect 7006 4564 7012 4616
rect 7064 4564 7070 4616
rect 7193 4607 7251 4613
rect 7193 4573 7205 4607
rect 7239 4604 7251 4607
rect 7834 4604 7840 4616
rect 7239 4576 7840 4604
rect 7239 4573 7251 4576
rect 7193 4567 7251 4573
rect 7834 4564 7840 4576
rect 7892 4604 7898 4616
rect 8110 4604 8116 4616
rect 7892 4576 8116 4604
rect 7892 4564 7898 4576
rect 8110 4564 8116 4576
rect 8168 4564 8174 4616
rect 8294 4564 8300 4616
rect 8352 4604 8358 4616
rect 9493 4607 9551 4613
rect 9493 4604 9505 4607
rect 8352 4576 9505 4604
rect 8352 4564 8358 4576
rect 9493 4573 9505 4576
rect 9539 4573 9551 4607
rect 9493 4567 9551 4573
rect 5960 4508 6960 4536
rect 7377 4539 7435 4545
rect 5960 4496 5966 4508
rect 7377 4505 7389 4539
rect 7423 4536 7435 4539
rect 8386 4536 8392 4548
rect 7423 4508 8392 4536
rect 7423 4505 7435 4508
rect 7377 4499 7435 4505
rect 8386 4496 8392 4508
rect 8444 4496 8450 4548
rect 8849 4539 8907 4545
rect 8849 4536 8861 4539
rect 8588 4508 8861 4536
rect 5316 4440 5580 4468
rect 7561 4471 7619 4477
rect 5316 4428 5322 4440
rect 7561 4437 7573 4471
rect 7607 4468 7619 4471
rect 7834 4468 7840 4480
rect 7607 4440 7840 4468
rect 7607 4437 7619 4440
rect 7561 4431 7619 4437
rect 7834 4428 7840 4440
rect 7892 4428 7898 4480
rect 8588 4477 8616 4508
rect 8849 4505 8861 4508
rect 8895 4505 8907 4539
rect 9508 4536 9536 4567
rect 9950 4564 9956 4616
rect 10008 4604 10014 4616
rect 10226 4604 10232 4616
rect 10008 4576 10232 4604
rect 10008 4564 10014 4576
rect 10226 4564 10232 4576
rect 10284 4564 10290 4616
rect 11238 4564 11244 4616
rect 11296 4604 11302 4616
rect 12158 4604 12164 4616
rect 11296 4576 12164 4604
rect 11296 4564 11302 4576
rect 12158 4564 12164 4576
rect 12216 4604 12222 4616
rect 12360 4604 12388 4635
rect 12986 4632 12992 4684
rect 13044 4632 13050 4684
rect 13170 4632 13176 4684
rect 13228 4672 13234 4684
rect 13449 4675 13507 4681
rect 13449 4672 13461 4675
rect 13228 4644 13461 4672
rect 13228 4632 13234 4644
rect 13449 4641 13461 4644
rect 13495 4641 13507 4675
rect 13556 4672 13584 4712
rect 15470 4700 15476 4712
rect 15528 4700 15534 4752
rect 17586 4700 17592 4752
rect 17644 4740 17650 4752
rect 18248 4740 18276 4780
rect 18325 4777 18337 4811
rect 18371 4808 18383 4811
rect 18966 4808 18972 4820
rect 18371 4780 18972 4808
rect 18371 4777 18383 4780
rect 18325 4771 18383 4777
rect 18966 4768 18972 4780
rect 19024 4768 19030 4820
rect 19702 4768 19708 4820
rect 19760 4808 19766 4820
rect 19886 4808 19892 4820
rect 19760 4780 19892 4808
rect 19760 4768 19766 4780
rect 19886 4768 19892 4780
rect 19944 4768 19950 4820
rect 20349 4811 20407 4817
rect 20349 4777 20361 4811
rect 20395 4777 20407 4811
rect 20349 4771 20407 4777
rect 20993 4811 21051 4817
rect 20993 4777 21005 4811
rect 21039 4808 21051 4811
rect 21818 4808 21824 4820
rect 21039 4780 21824 4808
rect 21039 4777 21051 4780
rect 20993 4771 21051 4777
rect 20364 4740 20392 4771
rect 21818 4768 21824 4780
rect 21876 4768 21882 4820
rect 21910 4768 21916 4820
rect 21968 4808 21974 4820
rect 21968 4780 22508 4808
rect 21968 4768 21974 4780
rect 21174 4740 21180 4752
rect 17644 4712 18184 4740
rect 18248 4712 20392 4740
rect 17644 4700 17650 4712
rect 13906 4672 13912 4684
rect 13556 4644 13912 4672
rect 13449 4635 13507 4641
rect 13906 4632 13912 4644
rect 13964 4632 13970 4684
rect 15105 4675 15163 4681
rect 15105 4672 15117 4675
rect 14384 4644 15117 4672
rect 12216 4576 12388 4604
rect 12713 4607 12771 4613
rect 12216 4564 12222 4576
rect 12713 4573 12725 4607
rect 12759 4604 12771 4607
rect 12894 4604 12900 4616
rect 12759 4576 12900 4604
rect 12759 4573 12771 4576
rect 12713 4567 12771 4573
rect 12894 4564 12900 4576
rect 12952 4564 12958 4616
rect 13081 4607 13139 4613
rect 13081 4573 13093 4607
rect 13127 4604 13139 4607
rect 13725 4607 13783 4613
rect 13725 4604 13737 4607
rect 13127 4576 13737 4604
rect 13127 4573 13139 4576
rect 13081 4567 13139 4573
rect 13188 4548 13216 4576
rect 13725 4573 13737 4576
rect 13771 4604 13783 4607
rect 14384 4604 14412 4644
rect 15105 4641 15117 4644
rect 15151 4641 15163 4675
rect 15105 4635 15163 4641
rect 13771 4576 14412 4604
rect 14737 4607 14795 4613
rect 13771 4573 13783 4576
rect 13725 4567 13783 4573
rect 14737 4573 14749 4607
rect 14783 4604 14795 4607
rect 14826 4604 14832 4616
rect 14783 4576 14832 4604
rect 14783 4573 14795 4576
rect 14737 4567 14795 4573
rect 14826 4564 14832 4576
rect 14884 4564 14890 4616
rect 15120 4604 15148 4635
rect 16114 4632 16120 4684
rect 16172 4632 16178 4684
rect 17218 4632 17224 4684
rect 17276 4632 17282 4684
rect 17862 4632 17868 4684
rect 17920 4632 17926 4684
rect 18156 4681 18184 4712
rect 18141 4675 18199 4681
rect 18141 4641 18153 4675
rect 18187 4641 18199 4675
rect 18141 4635 18199 4641
rect 18325 4675 18383 4681
rect 18325 4641 18337 4675
rect 18371 4641 18383 4675
rect 18325 4635 18383 4641
rect 16393 4607 16451 4613
rect 16393 4604 16405 4607
rect 15120 4576 16405 4604
rect 16393 4573 16405 4576
rect 16439 4573 16451 4607
rect 17313 4607 17371 4613
rect 17313 4604 17325 4607
rect 16393 4567 16451 4573
rect 16684 4576 17325 4604
rect 11146 4536 11152 4548
rect 9508 4508 11152 4536
rect 8849 4499 8907 4505
rect 11146 4496 11152 4508
rect 11204 4496 11210 4548
rect 11256 4508 13032 4536
rect 8573 4471 8631 4477
rect 8573 4437 8585 4471
rect 8619 4437 8631 4471
rect 8573 4431 8631 4437
rect 8662 4428 8668 4480
rect 8720 4468 8726 4480
rect 8757 4471 8815 4477
rect 8757 4468 8769 4471
rect 8720 4440 8769 4468
rect 8720 4428 8726 4440
rect 8757 4437 8769 4440
rect 8803 4437 8815 4471
rect 8757 4431 8815 4437
rect 8938 4428 8944 4480
rect 8996 4468 9002 4480
rect 9677 4471 9735 4477
rect 9677 4468 9689 4471
rect 8996 4440 9689 4468
rect 8996 4428 9002 4440
rect 9677 4437 9689 4440
rect 9723 4437 9735 4471
rect 9677 4431 9735 4437
rect 9766 4428 9772 4480
rect 9824 4468 9830 4480
rect 11256 4468 11284 4508
rect 9824 4440 11284 4468
rect 11609 4471 11667 4477
rect 9824 4428 9830 4440
rect 11609 4437 11621 4471
rect 11655 4468 11667 4471
rect 12342 4468 12348 4480
rect 11655 4440 12348 4468
rect 11655 4437 11667 4440
rect 11609 4431 11667 4437
rect 12342 4428 12348 4440
rect 12400 4428 12406 4480
rect 13004 4477 13032 4508
rect 13170 4496 13176 4548
rect 13228 4496 13234 4548
rect 14093 4539 14151 4545
rect 14093 4536 14105 4539
rect 13832 4508 14105 4536
rect 12989 4471 13047 4477
rect 12989 4437 13001 4471
rect 13035 4437 13047 4471
rect 12989 4431 13047 4437
rect 13262 4428 13268 4480
rect 13320 4468 13326 4480
rect 13832 4477 13860 4508
rect 14093 4505 14105 4508
rect 14139 4505 14151 4539
rect 14093 4499 14151 4505
rect 15378 4496 15384 4548
rect 15436 4536 15442 4548
rect 16684 4545 16712 4576
rect 17313 4573 17325 4576
rect 17359 4573 17371 4607
rect 17313 4567 17371 4573
rect 17405 4607 17463 4613
rect 17405 4573 17417 4607
rect 17451 4573 17463 4607
rect 17405 4567 17463 4573
rect 17497 4607 17555 4613
rect 17497 4573 17509 4607
rect 17543 4573 17555 4607
rect 17497 4567 17555 4573
rect 16669 4539 16727 4545
rect 15436 4508 16620 4536
rect 15436 4496 15442 4508
rect 13357 4471 13415 4477
rect 13357 4468 13369 4471
rect 13320 4440 13369 4468
rect 13320 4428 13326 4440
rect 13357 4437 13369 4440
rect 13403 4437 13415 4471
rect 13357 4431 13415 4437
rect 13817 4471 13875 4477
rect 13817 4437 13829 4471
rect 13863 4437 13875 4471
rect 13817 4431 13875 4437
rect 13998 4428 14004 4480
rect 14056 4428 14062 4480
rect 14918 4428 14924 4480
rect 14976 4428 14982 4480
rect 16206 4428 16212 4480
rect 16264 4428 16270 4480
rect 16592 4468 16620 4508
rect 16669 4505 16681 4539
rect 16715 4505 16727 4539
rect 17420 4536 17448 4567
rect 16669 4499 16727 4505
rect 16776 4508 17448 4536
rect 17512 4536 17540 4567
rect 18046 4564 18052 4616
rect 18104 4604 18110 4616
rect 18340 4604 18368 4635
rect 18414 4632 18420 4684
rect 18472 4632 18478 4684
rect 18506 4632 18512 4684
rect 18564 4632 18570 4684
rect 18693 4675 18751 4681
rect 18693 4641 18705 4675
rect 18739 4672 18751 4675
rect 18874 4672 18880 4684
rect 18739 4644 18880 4672
rect 18739 4641 18751 4644
rect 18693 4635 18751 4641
rect 18874 4632 18880 4644
rect 18932 4632 18938 4684
rect 19153 4675 19211 4681
rect 19153 4641 19165 4675
rect 19199 4641 19211 4675
rect 19153 4635 19211 4641
rect 19705 4675 19763 4681
rect 19705 4641 19717 4675
rect 19751 4672 19763 4675
rect 19794 4672 19800 4684
rect 19751 4644 19800 4672
rect 19751 4641 19763 4644
rect 19705 4635 19763 4641
rect 18104 4576 18368 4604
rect 18104 4564 18110 4576
rect 18598 4564 18604 4616
rect 18656 4604 18662 4616
rect 18785 4607 18843 4613
rect 18785 4604 18797 4607
rect 18656 4576 18797 4604
rect 18656 4564 18662 4576
rect 18785 4573 18797 4576
rect 18831 4604 18843 4607
rect 19061 4607 19119 4613
rect 19061 4604 19073 4607
rect 18831 4576 19073 4604
rect 18831 4573 18843 4576
rect 18785 4567 18843 4573
rect 19061 4573 19073 4576
rect 19107 4573 19119 4607
rect 19061 4567 19119 4573
rect 18690 4536 18696 4548
rect 17512 4508 18696 4536
rect 16776 4468 16804 4508
rect 16592 4440 16804 4468
rect 17034 4428 17040 4480
rect 17092 4428 17098 4480
rect 17420 4468 17448 4508
rect 18690 4496 18696 4508
rect 18748 4536 18754 4548
rect 19168 4536 19196 4635
rect 19794 4632 19800 4644
rect 19852 4632 19858 4684
rect 19889 4675 19947 4681
rect 19889 4641 19901 4675
rect 19935 4641 19947 4675
rect 19889 4635 19947 4641
rect 19705 4539 19763 4545
rect 19705 4536 19717 4539
rect 18748 4508 19717 4536
rect 18748 4496 18754 4508
rect 19705 4505 19717 4508
rect 19751 4505 19763 4539
rect 19705 4499 19763 4505
rect 17681 4471 17739 4477
rect 17681 4468 17693 4471
rect 17420 4440 17693 4468
rect 17681 4437 17693 4440
rect 17727 4437 17739 4471
rect 17681 4431 17739 4437
rect 18782 4428 18788 4480
rect 18840 4428 18846 4480
rect 19904 4468 19932 4635
rect 20364 4604 20392 4712
rect 20824 4712 21180 4740
rect 20533 4675 20591 4681
rect 20533 4641 20545 4675
rect 20579 4672 20591 4675
rect 20622 4672 20628 4684
rect 20579 4644 20628 4672
rect 20579 4641 20591 4644
rect 20533 4635 20591 4641
rect 20622 4632 20628 4644
rect 20680 4632 20686 4684
rect 20824 4681 20852 4712
rect 21174 4700 21180 4712
rect 21232 4700 21238 4752
rect 21726 4740 21732 4752
rect 21376 4712 21732 4740
rect 20809 4675 20867 4681
rect 20809 4641 20821 4675
rect 20855 4641 20867 4675
rect 20809 4635 20867 4641
rect 20901 4675 20959 4681
rect 20901 4641 20913 4675
rect 20947 4641 20959 4675
rect 20901 4635 20959 4641
rect 20916 4604 20944 4635
rect 21082 4632 21088 4684
rect 21140 4632 21146 4684
rect 21376 4681 21404 4712
rect 21726 4700 21732 4712
rect 21784 4700 21790 4752
rect 21836 4712 22048 4740
rect 21269 4675 21327 4681
rect 21269 4641 21281 4675
rect 21315 4641 21327 4675
rect 21269 4635 21327 4641
rect 21361 4675 21419 4681
rect 21361 4641 21373 4675
rect 21407 4641 21419 4675
rect 21361 4635 21419 4641
rect 20364 4576 20944 4604
rect 21284 4604 21312 4635
rect 21542 4632 21548 4684
rect 21600 4632 21606 4684
rect 21634 4632 21640 4684
rect 21692 4632 21698 4684
rect 21836 4672 21864 4712
rect 21744 4644 21864 4672
rect 21913 4675 21971 4681
rect 21744 4604 21772 4644
rect 21913 4641 21925 4675
rect 21959 4641 21971 4675
rect 21913 4635 21971 4641
rect 21284 4576 21772 4604
rect 20438 4496 20444 4548
rect 20496 4536 20502 4548
rect 20625 4539 20683 4545
rect 20625 4536 20637 4539
rect 20496 4508 20637 4536
rect 20496 4496 20502 4508
rect 20625 4505 20637 4508
rect 20671 4536 20683 4539
rect 21928 4536 21956 4635
rect 22020 4616 22048 4712
rect 22097 4675 22155 4681
rect 22097 4641 22109 4675
rect 22143 4641 22155 4675
rect 22097 4635 22155 4641
rect 22002 4564 22008 4616
rect 22060 4564 22066 4616
rect 22112 4604 22140 4635
rect 22278 4632 22284 4684
rect 22336 4632 22342 4684
rect 22480 4681 22508 4780
rect 22465 4675 22523 4681
rect 22465 4641 22477 4675
rect 22511 4641 22523 4675
rect 22465 4635 22523 4641
rect 23382 4604 23388 4616
rect 22112 4576 23388 4604
rect 22296 4548 22324 4576
rect 23382 4564 23388 4576
rect 23440 4564 23446 4616
rect 20671 4508 21956 4536
rect 20671 4505 20683 4508
rect 20625 4499 20683 4505
rect 22278 4496 22284 4548
rect 22336 4496 22342 4548
rect 21082 4468 21088 4480
rect 19904 4440 21088 4468
rect 21082 4428 21088 4440
rect 21140 4428 21146 4480
rect 21634 4428 21640 4480
rect 21692 4468 21698 4480
rect 21821 4471 21879 4477
rect 21821 4468 21833 4471
rect 21692 4440 21833 4468
rect 21692 4428 21698 4440
rect 21821 4437 21833 4440
rect 21867 4437 21879 4471
rect 21821 4431 21879 4437
rect 22094 4428 22100 4480
rect 22152 4468 22158 4480
rect 22465 4471 22523 4477
rect 22465 4468 22477 4471
rect 22152 4440 22477 4468
rect 22152 4428 22158 4440
rect 22465 4437 22477 4440
rect 22511 4437 22523 4471
rect 22465 4431 22523 4437
rect 552 4378 23368 4400
rect 552 4326 1366 4378
rect 1418 4326 1430 4378
rect 1482 4326 1494 4378
rect 1546 4326 1558 4378
rect 1610 4326 1622 4378
rect 1674 4326 1686 4378
rect 1738 4326 7366 4378
rect 7418 4326 7430 4378
rect 7482 4326 7494 4378
rect 7546 4326 7558 4378
rect 7610 4326 7622 4378
rect 7674 4326 7686 4378
rect 7738 4326 13366 4378
rect 13418 4326 13430 4378
rect 13482 4326 13494 4378
rect 13546 4326 13558 4378
rect 13610 4326 13622 4378
rect 13674 4326 13686 4378
rect 13738 4326 19366 4378
rect 19418 4326 19430 4378
rect 19482 4326 19494 4378
rect 19546 4326 19558 4378
rect 19610 4326 19622 4378
rect 19674 4326 19686 4378
rect 19738 4326 23368 4378
rect 552 4304 23368 4326
rect 2314 4224 2320 4276
rect 2372 4224 2378 4276
rect 4982 4224 4988 4276
rect 5040 4224 5046 4276
rect 5350 4224 5356 4276
rect 5408 4224 5414 4276
rect 6641 4267 6699 4273
rect 6641 4233 6653 4267
rect 6687 4264 6699 4267
rect 7006 4264 7012 4276
rect 6687 4236 7012 4264
rect 6687 4233 6699 4236
rect 6641 4227 6699 4233
rect 7006 4224 7012 4236
rect 7064 4224 7070 4276
rect 7561 4267 7619 4273
rect 7561 4233 7573 4267
rect 7607 4264 7619 4267
rect 7650 4264 7656 4276
rect 7607 4236 7656 4264
rect 7607 4233 7619 4236
rect 7561 4227 7619 4233
rect 7650 4224 7656 4236
rect 7708 4224 7714 4276
rect 7745 4267 7803 4273
rect 7745 4233 7757 4267
rect 7791 4264 7803 4267
rect 7834 4264 7840 4276
rect 7791 4236 7840 4264
rect 7791 4233 7803 4236
rect 7745 4227 7803 4233
rect 7834 4224 7840 4236
rect 7892 4224 7898 4276
rect 8018 4224 8024 4276
rect 8076 4224 8082 4276
rect 8386 4224 8392 4276
rect 8444 4224 8450 4276
rect 9674 4224 9680 4276
rect 9732 4264 9738 4276
rect 10413 4267 10471 4273
rect 10413 4264 10425 4267
rect 9732 4236 10425 4264
rect 9732 4224 9738 4236
rect 10413 4233 10425 4236
rect 10459 4233 10471 4267
rect 10413 4227 10471 4233
rect 12526 4224 12532 4276
rect 12584 4224 12590 4276
rect 12710 4224 12716 4276
rect 12768 4264 12774 4276
rect 13173 4267 13231 4273
rect 13173 4264 13185 4267
rect 12768 4236 13185 4264
rect 12768 4224 12774 4236
rect 13173 4233 13185 4236
rect 13219 4233 13231 4267
rect 14182 4264 14188 4276
rect 13173 4227 13231 4233
rect 13280 4236 14188 4264
rect 1765 4199 1823 4205
rect 1765 4165 1777 4199
rect 1811 4196 1823 4199
rect 3050 4196 3056 4208
rect 1811 4168 3056 4196
rect 1811 4165 1823 4168
rect 1765 4159 1823 4165
rect 3050 4156 3056 4168
rect 3108 4156 3114 4208
rect 4249 4199 4307 4205
rect 4249 4165 4261 4199
rect 4295 4196 4307 4199
rect 6365 4199 6423 4205
rect 4295 4168 5672 4196
rect 4295 4165 4307 4168
rect 4249 4159 4307 4165
rect 1489 4131 1547 4137
rect 1489 4097 1501 4131
rect 1535 4128 1547 4131
rect 1670 4128 1676 4140
rect 1535 4100 1676 4128
rect 1535 4097 1547 4100
rect 1489 4091 1547 4097
rect 1670 4088 1676 4100
rect 1728 4088 1734 4140
rect 1949 4131 2007 4137
rect 1949 4097 1961 4131
rect 1995 4128 2007 4131
rect 2593 4131 2651 4137
rect 2593 4128 2605 4131
rect 1995 4100 2605 4128
rect 1995 4097 2007 4100
rect 1949 4091 2007 4097
rect 2593 4097 2605 4100
rect 2639 4097 2651 4131
rect 2593 4091 2651 4097
rect 3973 4131 4031 4137
rect 3973 4097 3985 4131
rect 4019 4128 4031 4131
rect 4154 4128 4160 4140
rect 4019 4100 4160 4128
rect 4019 4097 4031 4100
rect 3973 4091 4031 4097
rect 4154 4088 4160 4100
rect 4212 4088 4218 4140
rect 4801 4131 4859 4137
rect 4801 4097 4813 4131
rect 4847 4128 4859 4131
rect 4847 4100 5488 4128
rect 4847 4097 4859 4100
rect 4801 4091 4859 4097
rect 5460 4072 5488 4100
rect 1397 4063 1455 4069
rect 1397 4029 1409 4063
rect 1443 4060 1455 4063
rect 1762 4060 1768 4072
rect 1443 4032 1768 4060
rect 1443 4029 1455 4032
rect 1397 4023 1455 4029
rect 1762 4020 1768 4032
rect 1820 4020 1826 4072
rect 2409 4063 2467 4069
rect 2409 4029 2421 4063
rect 2455 4029 2467 4063
rect 2409 4023 2467 4029
rect 2685 4063 2743 4069
rect 2685 4029 2697 4063
rect 2731 4060 2743 4063
rect 2774 4060 2780 4072
rect 2731 4032 2780 4060
rect 2731 4029 2743 4032
rect 2685 4023 2743 4029
rect 2424 3992 2452 4023
rect 2774 4020 2780 4032
rect 2832 4020 2838 4072
rect 3418 4020 3424 4072
rect 3476 4060 3482 4072
rect 3881 4063 3939 4069
rect 3881 4060 3893 4063
rect 3476 4032 3893 4060
rect 3476 4020 3482 4032
rect 3881 4029 3893 4032
rect 3927 4029 3939 4063
rect 3881 4023 3939 4029
rect 4338 4020 4344 4072
rect 4396 4020 4402 4072
rect 4522 4020 4528 4072
rect 4580 4060 4586 4072
rect 4709 4063 4767 4069
rect 4709 4060 4721 4063
rect 4580 4032 4721 4060
rect 4580 4020 4586 4032
rect 4709 4029 4721 4032
rect 4755 4029 4767 4063
rect 4709 4023 4767 4029
rect 4890 4020 4896 4072
rect 4948 4020 4954 4072
rect 4982 4020 4988 4072
rect 5040 4060 5046 4072
rect 5169 4063 5227 4069
rect 5169 4060 5181 4063
rect 5040 4032 5181 4060
rect 5040 4020 5046 4032
rect 5169 4029 5181 4032
rect 5215 4029 5227 4063
rect 5169 4023 5227 4029
rect 2958 3992 2964 4004
rect 2424 3964 2964 3992
rect 2958 3952 2964 3964
rect 3016 3952 3022 4004
rect 5184 3992 5212 4023
rect 5258 4020 5264 4072
rect 5316 4020 5322 4072
rect 5442 4020 5448 4072
rect 5500 4060 5506 4072
rect 5537 4063 5595 4069
rect 5537 4060 5549 4063
rect 5500 4032 5549 4060
rect 5500 4020 5506 4032
rect 5537 4029 5549 4032
rect 5583 4029 5595 4063
rect 5644 4060 5672 4168
rect 6365 4165 6377 4199
rect 6411 4165 6423 4199
rect 6365 4159 6423 4165
rect 5721 4131 5779 4137
rect 5721 4097 5733 4131
rect 5767 4128 5779 4131
rect 5905 4131 5963 4137
rect 5905 4128 5917 4131
rect 5767 4100 5917 4128
rect 5767 4097 5779 4100
rect 5721 4091 5779 4097
rect 5905 4097 5917 4100
rect 5951 4128 5963 4131
rect 6086 4128 6092 4140
rect 5951 4100 6092 4128
rect 5951 4097 5963 4100
rect 5905 4091 5963 4097
rect 6086 4088 6092 4100
rect 6144 4088 6150 4140
rect 5997 4063 6055 4069
rect 5997 4060 6009 4063
rect 5644 4032 6009 4060
rect 5537 4023 5595 4029
rect 5997 4029 6009 4032
rect 6043 4060 6055 4063
rect 6270 4060 6276 4072
rect 6043 4032 6276 4060
rect 6043 4029 6055 4032
rect 5997 4023 6055 4029
rect 6270 4020 6276 4032
rect 6328 4020 6334 4072
rect 6380 4060 6408 4159
rect 7024 4128 7052 4224
rect 7098 4156 7104 4208
rect 7156 4196 7162 4208
rect 8036 4196 8064 4224
rect 7156 4168 8064 4196
rect 7156 4156 7162 4168
rect 9398 4156 9404 4208
rect 9456 4196 9462 4208
rect 9582 4196 9588 4208
rect 9456 4168 9588 4196
rect 9456 4156 9462 4168
rect 9582 4156 9588 4168
rect 9640 4156 9646 4208
rect 9766 4156 9772 4208
rect 9824 4196 9830 4208
rect 10965 4199 11023 4205
rect 10965 4196 10977 4199
rect 9824 4168 10977 4196
rect 9824 4156 9830 4168
rect 10965 4165 10977 4168
rect 11011 4196 11023 4199
rect 11054 4196 11060 4208
rect 11011 4168 11060 4196
rect 11011 4165 11023 4168
rect 10965 4159 11023 4165
rect 11054 4156 11060 4168
rect 11112 4156 11118 4208
rect 11422 4156 11428 4208
rect 11480 4196 11486 4208
rect 11790 4196 11796 4208
rect 11480 4168 11796 4196
rect 11480 4156 11486 4168
rect 11790 4156 11796 4168
rect 11848 4196 11854 4208
rect 11848 4168 12756 4196
rect 11848 4156 11854 4168
rect 7469 4131 7527 4137
rect 7024 4100 7236 4128
rect 6825 4063 6883 4069
rect 6825 4060 6837 4063
rect 6380 4032 6837 4060
rect 6825 4029 6837 4032
rect 6871 4029 6883 4063
rect 6825 4023 6883 4029
rect 5350 3992 5356 4004
rect 5184 3964 5356 3992
rect 5350 3952 5356 3964
rect 5408 3952 5414 4004
rect 6840 3992 6868 4023
rect 7098 4020 7104 4072
rect 7156 4020 7162 4072
rect 7208 4069 7236 4100
rect 7469 4097 7481 4131
rect 7515 4128 7527 4131
rect 8110 4128 8116 4140
rect 7515 4100 8116 4128
rect 7515 4097 7527 4100
rect 7469 4091 7527 4097
rect 8110 4088 8116 4100
rect 8168 4088 8174 4140
rect 8938 4128 8944 4140
rect 8404 4100 8944 4128
rect 7193 4063 7251 4069
rect 7193 4029 7205 4063
rect 7239 4029 7251 4063
rect 7193 4023 7251 4029
rect 7650 4020 7656 4072
rect 7708 4060 7714 4072
rect 8404 4069 8432 4100
rect 8938 4088 8944 4100
rect 8996 4088 9002 4140
rect 9122 4088 9128 4140
rect 9180 4128 9186 4140
rect 11330 4128 11336 4140
rect 9180 4100 10088 4128
rect 9180 4088 9186 4100
rect 8389 4063 8447 4069
rect 7708 4032 8248 4060
rect 7708 4020 7714 4032
rect 8220 4001 8248 4032
rect 8389 4029 8401 4063
rect 8435 4029 8447 4063
rect 8389 4023 8447 4029
rect 8570 4020 8576 4072
rect 8628 4020 8634 4072
rect 9306 4020 9312 4072
rect 9364 4020 9370 4072
rect 9674 4060 9680 4072
rect 9416 4032 9680 4060
rect 7989 3995 8047 4001
rect 7989 3992 8001 3995
rect 6840 3964 8001 3992
rect 7989 3961 8001 3964
rect 8035 3961 8047 3995
rect 7989 3955 8047 3961
rect 8205 3995 8263 4001
rect 8205 3961 8217 3995
rect 8251 3961 8263 3995
rect 8205 3955 8263 3961
rect 8938 3952 8944 4004
rect 8996 3992 9002 4004
rect 9416 3992 9444 4032
rect 9674 4020 9680 4032
rect 9732 4020 9738 4072
rect 10060 4069 10088 4100
rect 11164 4100 11336 4128
rect 10045 4063 10103 4069
rect 10045 4029 10057 4063
rect 10091 4029 10103 4063
rect 10045 4023 10103 4029
rect 10686 4020 10692 4072
rect 10744 4020 10750 4072
rect 11164 4069 11192 4100
rect 11330 4088 11336 4100
rect 11388 4088 11394 4140
rect 11609 4131 11667 4137
rect 11609 4097 11621 4131
rect 11655 4128 11667 4131
rect 11977 4131 12035 4137
rect 11977 4128 11989 4131
rect 11655 4100 11989 4128
rect 11655 4097 11667 4100
rect 11609 4091 11667 4097
rect 11977 4097 11989 4100
rect 12023 4097 12035 4131
rect 11977 4091 12035 4097
rect 12253 4131 12311 4137
rect 12253 4097 12265 4131
rect 12299 4128 12311 4131
rect 12728 4128 12756 4168
rect 13280 4128 13308 4236
rect 14182 4224 14188 4236
rect 14240 4224 14246 4276
rect 14918 4224 14924 4276
rect 14976 4264 14982 4276
rect 21542 4264 21548 4276
rect 14976 4236 21548 4264
rect 14976 4224 14982 4236
rect 21542 4224 21548 4236
rect 21600 4224 21606 4276
rect 14090 4196 14096 4208
rect 12299 4100 12388 4128
rect 12299 4097 12311 4100
rect 12253 4091 12311 4097
rect 11149 4063 11207 4069
rect 11149 4029 11161 4063
rect 11195 4029 11207 4063
rect 11149 4023 11207 4029
rect 11238 4020 11244 4072
rect 11296 4060 11302 4072
rect 11517 4063 11575 4069
rect 11517 4060 11529 4063
rect 11296 4032 11529 4060
rect 11296 4020 11302 4032
rect 11517 4029 11529 4032
rect 11563 4029 11575 4063
rect 11517 4023 11575 4029
rect 11701 4063 11759 4069
rect 11701 4029 11713 4063
rect 11747 4060 11759 4063
rect 11790 4060 11796 4072
rect 11747 4032 11796 4060
rect 11747 4029 11759 4032
rect 11701 4023 11759 4029
rect 11790 4020 11796 4032
rect 11848 4020 11854 4072
rect 12069 4063 12127 4069
rect 12069 4029 12081 4063
rect 12115 4029 12127 4063
rect 12069 4023 12127 4029
rect 12161 4063 12219 4069
rect 12161 4029 12173 4063
rect 12207 4029 12219 4063
rect 12161 4023 12219 4029
rect 8996 3964 9444 3992
rect 8996 3952 9002 3964
rect 9582 3952 9588 4004
rect 9640 3952 9646 4004
rect 9769 3995 9827 4001
rect 9769 3961 9781 3995
rect 9815 3992 9827 3995
rect 10226 3992 10232 4004
rect 9815 3964 10232 3992
rect 9815 3961 9827 3964
rect 9769 3955 9827 3961
rect 10226 3952 10232 3964
rect 10284 3952 10290 4004
rect 10778 3952 10784 4004
rect 10836 3992 10842 4004
rect 12084 3992 12112 4023
rect 10836 3964 11560 3992
rect 10836 3952 10842 3964
rect 3053 3927 3111 3933
rect 3053 3893 3065 3927
rect 3099 3924 3111 3927
rect 3142 3924 3148 3936
rect 3099 3896 3148 3924
rect 3099 3893 3111 3896
rect 3053 3887 3111 3893
rect 3142 3884 3148 3896
rect 3200 3884 3206 3936
rect 4338 3884 4344 3936
rect 4396 3884 4402 3936
rect 6822 3884 6828 3936
rect 6880 3924 6886 3936
rect 7009 3927 7067 3933
rect 7009 3924 7021 3927
rect 6880 3896 7021 3924
rect 6880 3884 6886 3896
rect 7009 3893 7021 3896
rect 7055 3924 7067 3927
rect 7466 3924 7472 3936
rect 7055 3896 7472 3924
rect 7055 3893 7067 3896
rect 7009 3887 7067 3893
rect 7466 3884 7472 3896
rect 7524 3884 7530 3936
rect 7742 3884 7748 3936
rect 7800 3924 7806 3936
rect 7837 3927 7895 3933
rect 7837 3924 7849 3927
rect 7800 3896 7849 3924
rect 7800 3884 7806 3896
rect 7837 3893 7849 3896
rect 7883 3893 7895 3927
rect 7837 3887 7895 3893
rect 8757 3927 8815 3933
rect 8757 3893 8769 3927
rect 8803 3924 8815 3927
rect 9214 3924 9220 3936
rect 8803 3896 9220 3924
rect 8803 3893 8815 3896
rect 8757 3887 8815 3893
rect 9214 3884 9220 3896
rect 9272 3884 9278 3936
rect 9401 3927 9459 3933
rect 9401 3893 9413 3927
rect 9447 3924 9459 3927
rect 9674 3924 9680 3936
rect 9447 3896 9680 3924
rect 9447 3893 9459 3896
rect 9401 3887 9459 3893
rect 9674 3884 9680 3896
rect 9732 3884 9738 3936
rect 9953 3927 10011 3933
rect 9953 3893 9965 3927
rect 9999 3924 10011 3927
rect 10134 3924 10140 3936
rect 9999 3896 10140 3924
rect 9999 3893 10011 3896
rect 9953 3887 10011 3893
rect 10134 3884 10140 3896
rect 10192 3884 10198 3936
rect 10505 3927 10563 3933
rect 10505 3893 10517 3927
rect 10551 3924 10563 3927
rect 11330 3924 11336 3936
rect 10551 3896 11336 3924
rect 10551 3893 10563 3896
rect 10505 3887 10563 3893
rect 11330 3884 11336 3896
rect 11388 3884 11394 3936
rect 11532 3924 11560 3964
rect 11716 3964 12112 3992
rect 11716 3924 11744 3964
rect 11532 3896 11744 3924
rect 11790 3884 11796 3936
rect 11848 3884 11854 3936
rect 11974 3884 11980 3936
rect 12032 3924 12038 3936
rect 12176 3924 12204 4023
rect 12032 3896 12204 3924
rect 12360 3924 12388 4100
rect 12728 4100 13308 4128
rect 13924 4168 14096 4196
rect 12434 4020 12440 4072
rect 12492 4020 12498 4072
rect 12728 4069 12756 4100
rect 12713 4063 12771 4069
rect 12713 4029 12725 4063
rect 12759 4029 12771 4063
rect 12713 4023 12771 4029
rect 12802 4020 12808 4072
rect 12860 4020 12866 4072
rect 12894 4020 12900 4072
rect 12952 4060 12958 4072
rect 12989 4063 13047 4069
rect 12989 4060 13001 4063
rect 12952 4032 13001 4060
rect 12952 4020 12958 4032
rect 12989 4029 13001 4032
rect 13035 4029 13047 4063
rect 12989 4023 13047 4029
rect 13357 4063 13415 4069
rect 13357 4029 13369 4063
rect 13403 4060 13415 4063
rect 13722 4060 13728 4072
rect 13403 4032 13728 4060
rect 13403 4029 13415 4032
rect 13357 4023 13415 4029
rect 13722 4020 13728 4032
rect 13780 4020 13786 4072
rect 13814 4020 13820 4072
rect 13872 4020 13878 4072
rect 13924 4069 13952 4168
rect 14090 4156 14096 4168
rect 14148 4156 14154 4208
rect 14458 4156 14464 4208
rect 14516 4196 14522 4208
rect 14516 4168 16528 4196
rect 14516 4156 14522 4168
rect 13998 4088 14004 4140
rect 14056 4128 14062 4140
rect 14645 4131 14703 4137
rect 14645 4128 14657 4131
rect 14056 4100 14657 4128
rect 14056 4088 14062 4100
rect 14645 4097 14657 4100
rect 14691 4097 14703 4131
rect 14645 4091 14703 4097
rect 14734 4088 14740 4140
rect 14792 4088 14798 4140
rect 15194 4088 15200 4140
rect 15252 4088 15258 4140
rect 15286 4088 15292 4140
rect 15344 4088 15350 4140
rect 15378 4088 15384 4140
rect 15436 4088 15442 4140
rect 13909 4063 13967 4069
rect 13909 4029 13921 4063
rect 13955 4029 13967 4063
rect 13909 4023 13967 4029
rect 14093 4063 14151 4069
rect 14093 4029 14105 4063
rect 14139 4060 14151 4063
rect 14182 4060 14188 4072
rect 14139 4032 14188 4060
rect 14139 4029 14151 4032
rect 14093 4023 14151 4029
rect 14182 4020 14188 4032
rect 14240 4020 14246 4072
rect 14458 4020 14464 4072
rect 14516 4020 14522 4072
rect 14553 4063 14611 4069
rect 14553 4029 14565 4063
rect 14599 4060 14611 4063
rect 15396 4060 15424 4088
rect 14599 4032 15424 4060
rect 15473 4063 15531 4069
rect 14599 4029 14611 4032
rect 14553 4023 14611 4029
rect 15473 4029 15485 4063
rect 15519 4060 15531 4063
rect 15580 4060 15608 4168
rect 15654 4088 15660 4140
rect 15712 4128 15718 4140
rect 16209 4131 16267 4137
rect 16209 4128 16221 4131
rect 15712 4100 16221 4128
rect 15712 4088 15718 4100
rect 16209 4097 16221 4100
rect 16255 4097 16267 4131
rect 16209 4091 16267 4097
rect 16298 4088 16304 4140
rect 16356 4088 16362 4140
rect 16390 4088 16396 4140
rect 16448 4088 16454 4140
rect 15519 4032 15608 4060
rect 15519 4029 15531 4032
rect 15473 4023 15531 4029
rect 15838 4020 15844 4072
rect 15896 4020 15902 4072
rect 16114 4020 16120 4072
rect 16172 4020 16178 4072
rect 12618 3952 12624 4004
rect 12676 3992 12682 4004
rect 16500 3992 16528 4168
rect 18046 4156 18052 4208
rect 18104 4196 18110 4208
rect 22557 4199 22615 4205
rect 18104 4168 22324 4196
rect 18104 4156 18110 4168
rect 16577 4131 16635 4137
rect 16577 4097 16589 4131
rect 16623 4128 16635 4131
rect 16850 4128 16856 4140
rect 16623 4100 16856 4128
rect 16623 4097 16635 4100
rect 16577 4091 16635 4097
rect 16850 4088 16856 4100
rect 16908 4088 16914 4140
rect 19886 4128 19892 4140
rect 19168 4100 19892 4128
rect 19168 4069 19196 4100
rect 19886 4088 19892 4100
rect 19944 4088 19950 4140
rect 20364 4100 20760 4128
rect 19153 4063 19211 4069
rect 19153 4029 19165 4063
rect 19199 4029 19211 4063
rect 19153 4023 19211 4029
rect 19334 4020 19340 4072
rect 19392 4020 19398 4072
rect 19797 4063 19855 4069
rect 19797 4029 19809 4063
rect 19843 4060 19855 4063
rect 19904 4060 19932 4088
rect 20364 4072 20392 4100
rect 19843 4032 19932 4060
rect 19981 4063 20039 4069
rect 19843 4029 19855 4032
rect 19797 4023 19855 4029
rect 19981 4029 19993 4063
rect 20027 4060 20039 4063
rect 20254 4060 20260 4072
rect 20027 4032 20260 4060
rect 20027 4029 20039 4032
rect 19981 4023 20039 4029
rect 20254 4020 20260 4032
rect 20312 4020 20318 4072
rect 20346 4020 20352 4072
rect 20404 4020 20410 4072
rect 20438 4020 20444 4072
rect 20496 4020 20502 4072
rect 20622 4020 20628 4072
rect 20680 4020 20686 4072
rect 20732 4069 20760 4100
rect 21082 4088 21088 4140
rect 21140 4088 21146 4140
rect 20717 4063 20775 4069
rect 20717 4029 20729 4063
rect 20763 4029 20775 4063
rect 20717 4023 20775 4029
rect 21174 4020 21180 4072
rect 21232 4020 21238 4072
rect 21358 4069 21364 4072
rect 21331 4063 21364 4069
rect 21331 4029 21343 4063
rect 21331 4023 21364 4029
rect 21358 4020 21364 4023
rect 21416 4020 21422 4072
rect 21450 4020 21456 4072
rect 21508 4060 21514 4072
rect 21821 4063 21879 4069
rect 21821 4060 21833 4063
rect 21508 4032 21833 4060
rect 21508 4020 21514 4032
rect 21821 4029 21833 4032
rect 21867 4060 21879 4063
rect 21910 4060 21916 4072
rect 21867 4032 21916 4060
rect 21867 4029 21879 4032
rect 21821 4023 21879 4029
rect 21910 4020 21916 4032
rect 21968 4020 21974 4072
rect 22002 4020 22008 4072
rect 22060 4020 22066 4072
rect 22094 4020 22100 4072
rect 22152 4020 22158 4072
rect 22296 4069 22324 4168
rect 22557 4165 22569 4199
rect 22603 4196 22615 4199
rect 22922 4196 22928 4208
rect 22603 4168 22928 4196
rect 22603 4165 22615 4168
rect 22557 4159 22615 4165
rect 22922 4156 22928 4168
rect 22980 4156 22986 4208
rect 22281 4063 22339 4069
rect 22281 4029 22293 4063
rect 22327 4029 22339 4063
rect 22281 4023 22339 4029
rect 22373 4063 22431 4069
rect 22373 4029 22385 4063
rect 22419 4029 22431 4063
rect 22373 4023 22431 4029
rect 22741 4063 22799 4069
rect 22741 4029 22753 4063
rect 22787 4060 22799 4063
rect 23106 4060 23112 4072
rect 22787 4032 23112 4060
rect 22787 4029 22799 4032
rect 22741 4023 22799 4029
rect 19889 3995 19947 4001
rect 19889 3992 19901 3995
rect 12676 3964 15700 3992
rect 16500 3964 19901 3992
rect 12676 3952 12682 3964
rect 15672 3936 15700 3964
rect 19889 3961 19901 3964
rect 19935 3961 19947 3995
rect 19889 3955 19947 3961
rect 21545 3995 21603 4001
rect 21545 3961 21557 3995
rect 21591 3992 21603 3995
rect 21591 3964 22094 3992
rect 21591 3961 21603 3964
rect 21545 3955 21603 3961
rect 12802 3924 12808 3936
rect 12360 3896 12808 3924
rect 12032 3884 12038 3896
rect 12802 3884 12808 3896
rect 12860 3884 12866 3936
rect 12986 3884 12992 3936
rect 13044 3884 13050 3936
rect 13170 3884 13176 3936
rect 13228 3924 13234 3936
rect 13633 3927 13691 3933
rect 13633 3924 13645 3927
rect 13228 3896 13645 3924
rect 13228 3884 13234 3896
rect 13633 3893 13645 3896
rect 13679 3893 13691 3927
rect 13633 3887 13691 3893
rect 13814 3884 13820 3936
rect 13872 3924 13878 3936
rect 14001 3927 14059 3933
rect 14001 3924 14013 3927
rect 13872 3896 14013 3924
rect 13872 3884 13878 3896
rect 14001 3893 14013 3896
rect 14047 3893 14059 3927
rect 14001 3887 14059 3893
rect 14918 3884 14924 3936
rect 14976 3884 14982 3936
rect 15013 3927 15071 3933
rect 15013 3893 15025 3927
rect 15059 3924 15071 3927
rect 15102 3924 15108 3936
rect 15059 3896 15108 3924
rect 15059 3893 15071 3896
rect 15013 3887 15071 3893
rect 15102 3884 15108 3896
rect 15160 3884 15166 3936
rect 15654 3884 15660 3936
rect 15712 3884 15718 3936
rect 16758 3884 16764 3936
rect 16816 3924 16822 3936
rect 19245 3927 19303 3933
rect 19245 3924 19257 3927
rect 16816 3896 19257 3924
rect 16816 3884 16822 3896
rect 19245 3893 19257 3896
rect 19291 3893 19303 3927
rect 19245 3887 19303 3893
rect 19334 3884 19340 3936
rect 19392 3924 19398 3936
rect 20070 3924 20076 3936
rect 19392 3896 20076 3924
rect 19392 3884 19398 3896
rect 20070 3884 20076 3896
rect 20128 3884 20134 3936
rect 20162 3884 20168 3936
rect 20220 3884 20226 3936
rect 20346 3884 20352 3936
rect 20404 3924 20410 3936
rect 20533 3927 20591 3933
rect 20533 3924 20545 3927
rect 20404 3896 20545 3924
rect 20404 3884 20410 3896
rect 20533 3893 20545 3896
rect 20579 3893 20591 3927
rect 20533 3887 20591 3893
rect 20898 3884 20904 3936
rect 20956 3884 20962 3936
rect 21174 3884 21180 3936
rect 21232 3924 21238 3936
rect 21637 3927 21695 3933
rect 21637 3924 21649 3927
rect 21232 3896 21649 3924
rect 21232 3884 21238 3896
rect 21637 3893 21649 3896
rect 21683 3893 21695 3927
rect 22066 3924 22094 3964
rect 22186 3952 22192 4004
rect 22244 3992 22250 4004
rect 22388 3992 22416 4023
rect 23106 4020 23112 4032
rect 23164 4020 23170 4072
rect 23382 3992 23388 4004
rect 22244 3964 22416 3992
rect 22480 3964 23388 3992
rect 22244 3952 22250 3964
rect 22480 3924 22508 3964
rect 23382 3952 23388 3964
rect 23440 3952 23446 4004
rect 22066 3896 22508 3924
rect 21637 3887 21695 3893
rect 22830 3884 22836 3936
rect 22888 3884 22894 3936
rect 552 3834 23368 3856
rect 552 3782 4366 3834
rect 4418 3782 4430 3834
rect 4482 3782 4494 3834
rect 4546 3782 4558 3834
rect 4610 3782 4622 3834
rect 4674 3782 4686 3834
rect 4738 3782 10366 3834
rect 10418 3782 10430 3834
rect 10482 3782 10494 3834
rect 10546 3782 10558 3834
rect 10610 3782 10622 3834
rect 10674 3782 10686 3834
rect 10738 3782 16366 3834
rect 16418 3782 16430 3834
rect 16482 3782 16494 3834
rect 16546 3782 16558 3834
rect 16610 3782 16622 3834
rect 16674 3782 16686 3834
rect 16738 3782 22366 3834
rect 22418 3782 22430 3834
rect 22482 3782 22494 3834
rect 22546 3782 22558 3834
rect 22610 3782 22622 3834
rect 22674 3782 22686 3834
rect 22738 3782 23368 3834
rect 552 3760 23368 3782
rect 1670 3680 1676 3732
rect 1728 3680 1734 3732
rect 3513 3723 3571 3729
rect 3513 3689 3525 3723
rect 3559 3720 3571 3723
rect 7561 3723 7619 3729
rect 3559 3692 7144 3720
rect 3559 3689 3571 3692
rect 3513 3683 3571 3689
rect 1210 3612 1216 3664
rect 1268 3612 1274 3664
rect 6086 3612 6092 3664
rect 6144 3612 6150 3664
rect 6178 3612 6184 3664
rect 6236 3652 6242 3664
rect 6457 3655 6515 3661
rect 6457 3652 6469 3655
rect 6236 3624 6469 3652
rect 6236 3612 6242 3624
rect 6457 3621 6469 3624
rect 6503 3621 6515 3655
rect 6457 3615 6515 3621
rect 3142 3544 3148 3596
rect 3200 3544 3206 3596
rect 4246 3544 4252 3596
rect 4304 3584 4310 3596
rect 4525 3587 4583 3593
rect 4525 3584 4537 3587
rect 4304 3556 4537 3584
rect 4304 3544 4310 3556
rect 4525 3553 4537 3556
rect 4571 3553 4583 3587
rect 4525 3547 4583 3553
rect 4709 3587 4767 3593
rect 4709 3553 4721 3587
rect 4755 3584 4767 3587
rect 5166 3584 5172 3596
rect 4755 3556 5172 3584
rect 4755 3553 4767 3556
rect 4709 3547 4767 3553
rect 5166 3544 5172 3556
rect 5224 3544 5230 3596
rect 6270 3544 6276 3596
rect 6328 3544 6334 3596
rect 7116 3593 7144 3692
rect 7561 3689 7573 3723
rect 7607 3720 7619 3723
rect 7926 3720 7932 3732
rect 7607 3692 7932 3720
rect 7607 3689 7619 3692
rect 7561 3683 7619 3689
rect 7926 3680 7932 3692
rect 7984 3680 7990 3732
rect 8846 3680 8852 3732
rect 8904 3720 8910 3732
rect 9582 3720 9588 3732
rect 8904 3692 9076 3720
rect 8904 3680 8910 3692
rect 7193 3655 7251 3661
rect 7193 3621 7205 3655
rect 7239 3652 7251 3655
rect 7834 3652 7840 3664
rect 7239 3624 7840 3652
rect 7239 3621 7251 3624
rect 7193 3615 7251 3621
rect 7834 3612 7840 3624
rect 7892 3612 7898 3664
rect 7101 3587 7159 3593
rect 7101 3553 7113 3587
rect 7147 3553 7159 3587
rect 7101 3547 7159 3553
rect 7282 3544 7288 3596
rect 7340 3584 7346 3596
rect 7377 3587 7435 3593
rect 7377 3584 7389 3587
rect 7340 3556 7389 3584
rect 7340 3544 7346 3556
rect 7377 3553 7389 3556
rect 7423 3553 7435 3587
rect 7377 3547 7435 3553
rect 8205 3587 8263 3593
rect 8205 3553 8217 3587
rect 8251 3584 8263 3587
rect 8294 3584 8300 3596
rect 8251 3556 8300 3584
rect 8251 3553 8263 3556
rect 8205 3547 8263 3553
rect 8294 3544 8300 3556
rect 8352 3544 8358 3596
rect 8389 3587 8447 3593
rect 8389 3553 8401 3587
rect 8435 3584 8447 3587
rect 8481 3587 8539 3593
rect 8481 3584 8493 3587
rect 8435 3556 8493 3584
rect 8435 3553 8447 3556
rect 8389 3547 8447 3553
rect 8481 3553 8493 3556
rect 8527 3553 8539 3587
rect 8481 3547 8539 3553
rect 8665 3587 8723 3593
rect 8665 3553 8677 3587
rect 8711 3584 8723 3587
rect 8754 3584 8760 3596
rect 8711 3556 8760 3584
rect 8711 3553 8723 3556
rect 8665 3547 8723 3553
rect 3050 3476 3056 3528
rect 3108 3476 3114 3528
rect 8496 3516 8524 3547
rect 8754 3544 8760 3556
rect 8812 3544 8818 3596
rect 8938 3544 8944 3596
rect 8996 3544 9002 3596
rect 9048 3593 9076 3692
rect 9140 3692 9588 3720
rect 9140 3593 9168 3692
rect 9582 3680 9588 3692
rect 9640 3720 9646 3732
rect 9640 3692 9915 3720
rect 9640 3680 9646 3692
rect 9674 3652 9680 3664
rect 9416 3624 9680 3652
rect 9033 3587 9091 3593
rect 9033 3553 9045 3587
rect 9079 3553 9091 3587
rect 9033 3547 9091 3553
rect 9125 3587 9183 3593
rect 9125 3553 9137 3587
rect 9171 3553 9183 3587
rect 9125 3547 9183 3553
rect 9217 3587 9275 3593
rect 9217 3553 9229 3587
rect 9263 3584 9275 3587
rect 9306 3584 9312 3596
rect 9263 3556 9312 3584
rect 9263 3553 9275 3556
rect 9217 3547 9275 3553
rect 9306 3544 9312 3556
rect 9364 3544 9370 3596
rect 9416 3593 9444 3624
rect 9674 3612 9680 3624
rect 9732 3612 9738 3664
rect 9766 3612 9772 3664
rect 9824 3612 9830 3664
rect 9401 3587 9459 3593
rect 9401 3553 9413 3587
rect 9447 3553 9459 3587
rect 9401 3547 9459 3553
rect 9490 3544 9496 3596
rect 9548 3584 9554 3596
rect 9585 3587 9643 3593
rect 9585 3584 9597 3587
rect 9548 3556 9597 3584
rect 9548 3544 9554 3556
rect 9585 3553 9597 3556
rect 9631 3553 9643 3587
rect 9784 3584 9812 3612
rect 9585 3547 9643 3553
rect 9692 3556 9812 3584
rect 9692 3525 9720 3556
rect 9677 3519 9735 3525
rect 9677 3516 9689 3519
rect 8496 3488 9689 3516
rect 9677 3485 9689 3488
rect 9723 3485 9735 3519
rect 9677 3479 9735 3485
rect 9766 3476 9772 3528
rect 9824 3476 9830 3528
rect 9887 3516 9915 3692
rect 10226 3680 10232 3732
rect 10284 3720 10290 3732
rect 12805 3723 12863 3729
rect 10284 3692 12296 3720
rect 10284 3680 10290 3692
rect 12268 3661 12296 3692
rect 12805 3689 12817 3723
rect 12851 3720 12863 3723
rect 12894 3720 12900 3732
rect 12851 3692 12900 3720
rect 12851 3689 12863 3692
rect 12805 3683 12863 3689
rect 12253 3655 12311 3661
rect 9968 3624 11836 3652
rect 9968 3593 9996 3624
rect 9953 3587 10011 3593
rect 9953 3553 9965 3587
rect 9999 3553 10011 3587
rect 9953 3547 10011 3553
rect 10134 3544 10140 3596
rect 10192 3584 10198 3596
rect 10413 3587 10471 3593
rect 10413 3584 10425 3587
rect 10192 3556 10425 3584
rect 10192 3544 10198 3556
rect 10413 3553 10425 3556
rect 10459 3553 10471 3587
rect 10413 3547 10471 3553
rect 10502 3544 10508 3596
rect 10560 3544 10566 3596
rect 10962 3544 10968 3596
rect 11020 3584 11026 3596
rect 11241 3587 11299 3593
rect 11241 3584 11253 3587
rect 11020 3556 11253 3584
rect 11020 3544 11026 3556
rect 11241 3553 11253 3556
rect 11287 3553 11299 3587
rect 11241 3547 11299 3553
rect 11330 3544 11336 3596
rect 11388 3544 11394 3596
rect 9887 3488 10364 3516
rect 1118 3408 1124 3460
rect 1176 3448 1182 3460
rect 1489 3451 1547 3457
rect 1489 3448 1501 3451
rect 1176 3420 1501 3448
rect 1176 3408 1182 3420
rect 1489 3417 1501 3420
rect 1535 3417 1547 3451
rect 1489 3411 1547 3417
rect 8573 3451 8631 3457
rect 8573 3417 8585 3451
rect 8619 3448 8631 3451
rect 9306 3448 9312 3460
rect 8619 3420 9312 3448
rect 8619 3417 8631 3420
rect 8573 3411 8631 3417
rect 9306 3408 9312 3420
rect 9364 3408 9370 3460
rect 9490 3408 9496 3460
rect 9548 3448 9554 3460
rect 10229 3451 10287 3457
rect 10229 3448 10241 3451
rect 9548 3420 10241 3448
rect 9548 3408 9554 3420
rect 10229 3417 10241 3420
rect 10275 3417 10287 3451
rect 10336 3448 10364 3488
rect 10594 3476 10600 3528
rect 10652 3476 10658 3528
rect 10686 3476 10692 3528
rect 10744 3476 10750 3528
rect 10778 3476 10784 3528
rect 10836 3516 10842 3528
rect 11149 3519 11207 3525
rect 11149 3516 11161 3519
rect 10836 3488 11161 3516
rect 10836 3476 10842 3488
rect 11149 3485 11161 3488
rect 11195 3485 11207 3519
rect 11149 3479 11207 3485
rect 11348 3448 11376 3544
rect 11422 3476 11428 3528
rect 11480 3476 11486 3528
rect 11808 3516 11836 3624
rect 12253 3621 12265 3655
rect 12299 3652 12311 3655
rect 12618 3652 12624 3664
rect 12299 3624 12624 3652
rect 12299 3621 12311 3624
rect 12253 3615 12311 3621
rect 12618 3612 12624 3624
rect 12676 3612 12682 3664
rect 11882 3544 11888 3596
rect 11940 3584 11946 3596
rect 11977 3587 12035 3593
rect 11977 3584 11989 3587
rect 11940 3556 11989 3584
rect 11940 3544 11946 3556
rect 11977 3553 11989 3556
rect 12023 3553 12035 3587
rect 11977 3547 12035 3553
rect 12066 3544 12072 3596
rect 12124 3544 12130 3596
rect 12342 3544 12348 3596
rect 12400 3544 12406 3596
rect 12434 3516 12440 3528
rect 11808 3488 12440 3516
rect 12434 3476 12440 3488
rect 12492 3476 12498 3528
rect 12621 3519 12679 3525
rect 12621 3485 12633 3519
rect 12667 3516 12679 3519
rect 12820 3516 12848 3683
rect 12894 3680 12900 3692
rect 12952 3680 12958 3732
rect 14645 3723 14703 3729
rect 14645 3689 14657 3723
rect 14691 3720 14703 3723
rect 14734 3720 14740 3732
rect 14691 3692 14740 3720
rect 14691 3689 14703 3692
rect 14645 3683 14703 3689
rect 14734 3680 14740 3692
rect 14792 3680 14798 3732
rect 14826 3680 14832 3732
rect 14884 3680 14890 3732
rect 16114 3680 16120 3732
rect 16172 3720 16178 3732
rect 16666 3720 16672 3732
rect 16172 3692 16672 3720
rect 16172 3680 16178 3692
rect 16666 3680 16672 3692
rect 16724 3680 16730 3732
rect 19794 3720 19800 3732
rect 16776 3692 19800 3720
rect 14844 3652 14872 3680
rect 15013 3655 15071 3661
rect 15013 3652 15025 3655
rect 14844 3624 15025 3652
rect 15013 3621 15025 3624
rect 15059 3621 15071 3655
rect 15013 3615 15071 3621
rect 15654 3612 15660 3664
rect 15712 3652 15718 3664
rect 16776 3652 16804 3692
rect 19794 3680 19800 3692
rect 19852 3680 19858 3732
rect 21358 3720 21364 3732
rect 21284 3692 21364 3720
rect 17954 3652 17960 3664
rect 15712 3624 16436 3652
rect 15712 3612 15718 3624
rect 12897 3587 12955 3593
rect 12897 3553 12909 3587
rect 12943 3584 12955 3587
rect 12943 3556 13216 3584
rect 12943 3553 12955 3556
rect 12897 3547 12955 3553
rect 12667 3488 12848 3516
rect 12667 3485 12679 3488
rect 12621 3479 12679 3485
rect 12529 3451 12587 3457
rect 12529 3448 12541 3451
rect 10336 3420 11376 3448
rect 11992 3420 12541 3448
rect 10229 3411 10287 3417
rect 11992 3392 12020 3420
rect 12529 3417 12541 3420
rect 12575 3417 12587 3451
rect 12529 3411 12587 3417
rect 12802 3408 12808 3460
rect 12860 3448 12866 3460
rect 13188 3448 13216 3556
rect 13814 3544 13820 3596
rect 13872 3544 13878 3596
rect 14090 3544 14096 3596
rect 14148 3544 14154 3596
rect 14829 3587 14887 3593
rect 14829 3553 14841 3587
rect 14875 3584 14887 3587
rect 14875 3556 15884 3584
rect 14875 3553 14887 3556
rect 14829 3547 14887 3553
rect 15856 3528 15884 3556
rect 15930 3544 15936 3596
rect 15988 3584 15994 3596
rect 16408 3593 16436 3624
rect 16500 3624 16804 3652
rect 17236 3624 17960 3652
rect 16301 3587 16359 3593
rect 16301 3584 16313 3587
rect 15988 3556 16313 3584
rect 15988 3544 15994 3556
rect 16301 3553 16313 3556
rect 16347 3553 16359 3587
rect 16301 3547 16359 3553
rect 16393 3587 16451 3593
rect 16393 3553 16405 3587
rect 16439 3553 16451 3587
rect 16393 3547 16451 3553
rect 13262 3476 13268 3528
rect 13320 3516 13326 3528
rect 13909 3519 13967 3525
rect 13909 3516 13921 3519
rect 13320 3488 13921 3516
rect 13320 3476 13326 3488
rect 13909 3485 13921 3488
rect 13955 3485 13967 3519
rect 13909 3479 13967 3485
rect 14001 3519 14059 3525
rect 14001 3485 14013 3519
rect 14047 3516 14059 3519
rect 15378 3516 15384 3528
rect 14047 3488 15384 3516
rect 14047 3485 14059 3488
rect 14001 3479 14059 3485
rect 15378 3476 15384 3488
rect 15436 3476 15442 3528
rect 15838 3476 15844 3528
rect 15896 3516 15902 3528
rect 16500 3516 16528 3624
rect 16577 3587 16635 3593
rect 16577 3553 16589 3587
rect 16623 3553 16635 3587
rect 16577 3547 16635 3553
rect 15896 3488 16528 3516
rect 16592 3516 16620 3547
rect 16666 3544 16672 3596
rect 16724 3544 16730 3596
rect 17236 3593 17264 3624
rect 17954 3612 17960 3624
rect 18012 3612 18018 3664
rect 18874 3652 18880 3664
rect 18524 3624 18880 3652
rect 17221 3587 17279 3593
rect 17221 3553 17233 3587
rect 17267 3553 17279 3587
rect 17221 3547 17279 3553
rect 17405 3587 17463 3593
rect 17405 3553 17417 3587
rect 17451 3584 17463 3587
rect 17681 3587 17739 3593
rect 17681 3584 17693 3587
rect 17451 3556 17693 3584
rect 17451 3553 17463 3556
rect 17405 3547 17463 3553
rect 17681 3553 17693 3556
rect 17727 3553 17739 3587
rect 17681 3547 17739 3553
rect 17865 3587 17923 3593
rect 17865 3553 17877 3587
rect 17911 3584 17923 3587
rect 18524 3584 18552 3624
rect 18874 3612 18880 3624
rect 18932 3612 18938 3664
rect 20162 3652 20168 3664
rect 19306 3624 20168 3652
rect 17911 3556 18552 3584
rect 18601 3587 18659 3593
rect 17911 3553 17923 3556
rect 17865 3547 17923 3553
rect 18601 3553 18613 3587
rect 18647 3584 18659 3587
rect 19153 3587 19211 3593
rect 19153 3584 19165 3587
rect 18647 3556 19165 3584
rect 18647 3553 18659 3556
rect 18601 3547 18659 3553
rect 19153 3553 19165 3556
rect 19199 3584 19211 3587
rect 19306 3584 19334 3624
rect 20162 3612 20168 3624
rect 20220 3652 20226 3664
rect 21284 3652 21312 3692
rect 21358 3680 21364 3692
rect 21416 3680 21422 3732
rect 22278 3652 22284 3664
rect 20220 3624 21312 3652
rect 20220 3612 20226 3624
rect 19199 3556 19334 3584
rect 19199 3553 19211 3556
rect 19153 3547 19211 3553
rect 17313 3519 17371 3525
rect 17313 3516 17325 3519
rect 16592 3488 17325 3516
rect 15896 3476 15902 3488
rect 17313 3485 17325 3488
rect 17359 3485 17371 3519
rect 17696 3516 17724 3547
rect 19518 3544 19524 3596
rect 19576 3544 19582 3596
rect 19705 3587 19763 3593
rect 19705 3553 19717 3587
rect 19751 3584 19763 3587
rect 19794 3584 19800 3596
rect 19751 3556 19800 3584
rect 19751 3553 19763 3556
rect 19705 3547 19763 3553
rect 19794 3544 19800 3556
rect 19852 3544 19858 3596
rect 19886 3544 19892 3596
rect 19944 3544 19950 3596
rect 20257 3587 20315 3593
rect 20257 3553 20269 3587
rect 20303 3584 20315 3587
rect 20809 3587 20867 3593
rect 20809 3584 20821 3587
rect 20303 3556 20821 3584
rect 20303 3553 20315 3556
rect 20257 3547 20315 3553
rect 20809 3553 20821 3556
rect 20855 3584 20867 3587
rect 20898 3584 20904 3596
rect 20855 3556 20904 3584
rect 20855 3553 20867 3556
rect 20809 3547 20867 3553
rect 20898 3544 20904 3556
rect 20956 3544 20962 3596
rect 18506 3516 18512 3528
rect 17696 3488 18512 3516
rect 17313 3479 17371 3485
rect 18506 3476 18512 3488
rect 18564 3476 18570 3528
rect 18874 3476 18880 3528
rect 18932 3476 18938 3528
rect 19334 3516 19340 3528
rect 19306 3476 19340 3516
rect 19392 3476 19398 3528
rect 19429 3519 19487 3525
rect 19429 3485 19441 3519
rect 19475 3516 19487 3519
rect 19904 3516 19932 3544
rect 19475 3488 19932 3516
rect 19475 3485 19487 3488
rect 19429 3479 19487 3485
rect 20070 3476 20076 3528
rect 20128 3516 20134 3528
rect 20533 3519 20591 3525
rect 20533 3516 20545 3519
rect 20128 3488 20545 3516
rect 20128 3476 20134 3488
rect 20533 3485 20545 3488
rect 20579 3485 20591 3519
rect 20533 3479 20591 3485
rect 21082 3476 21088 3528
rect 21140 3476 21146 3528
rect 21284 3516 21312 3624
rect 21560 3624 22284 3652
rect 21361 3587 21419 3593
rect 21361 3553 21373 3587
rect 21407 3584 21419 3587
rect 21560 3584 21588 3624
rect 22278 3612 22284 3624
rect 22336 3612 22342 3664
rect 21407 3556 21588 3584
rect 21637 3587 21695 3593
rect 21407 3553 21419 3556
rect 21361 3547 21419 3553
rect 21637 3553 21649 3587
rect 21683 3553 21695 3587
rect 21637 3547 21695 3553
rect 21652 3516 21680 3547
rect 21910 3544 21916 3596
rect 21968 3584 21974 3596
rect 22097 3587 22155 3593
rect 22097 3584 22109 3587
rect 21968 3556 22109 3584
rect 21968 3544 21974 3556
rect 22097 3553 22109 3556
rect 22143 3553 22155 3587
rect 22097 3547 22155 3553
rect 22189 3587 22247 3593
rect 22189 3553 22201 3587
rect 22235 3553 22247 3587
rect 22189 3547 22247 3553
rect 22649 3587 22707 3593
rect 22649 3553 22661 3587
rect 22695 3584 22707 3587
rect 23014 3584 23020 3596
rect 22695 3556 23020 3584
rect 22695 3553 22707 3556
rect 22649 3547 22707 3553
rect 21284 3488 21680 3516
rect 22204 3516 22232 3547
rect 23014 3544 23020 3556
rect 23072 3544 23078 3596
rect 23198 3516 23204 3528
rect 22204 3488 23204 3516
rect 23198 3476 23204 3488
rect 23256 3476 23262 3528
rect 16758 3448 16764 3460
rect 12860 3420 16764 3448
rect 12860 3408 12866 3420
rect 16758 3408 16764 3420
rect 16816 3408 16822 3460
rect 17678 3408 17684 3460
rect 17736 3448 17742 3460
rect 17736 3420 18000 3448
rect 17736 3408 17742 3420
rect 4614 3340 4620 3392
rect 4672 3340 4678 3392
rect 8294 3340 8300 3392
rect 8352 3340 8358 3392
rect 8754 3340 8760 3392
rect 8812 3340 8818 3392
rect 8846 3340 8852 3392
rect 8904 3380 8910 3392
rect 9950 3380 9956 3392
rect 8904 3352 9956 3380
rect 8904 3340 8910 3352
rect 9950 3340 9956 3352
rect 10008 3340 10014 3392
rect 10042 3340 10048 3392
rect 10100 3380 10106 3392
rect 10137 3383 10195 3389
rect 10137 3380 10149 3383
rect 10100 3352 10149 3380
rect 10100 3340 10106 3352
rect 10137 3349 10149 3352
rect 10183 3349 10195 3383
rect 10137 3343 10195 3349
rect 10318 3340 10324 3392
rect 10376 3380 10382 3392
rect 10965 3383 11023 3389
rect 10965 3380 10977 3383
rect 10376 3352 10977 3380
rect 10376 3340 10382 3352
rect 10965 3349 10977 3352
rect 11011 3349 11023 3383
rect 10965 3343 11023 3349
rect 11974 3340 11980 3392
rect 12032 3340 12038 3392
rect 12253 3383 12311 3389
rect 12253 3349 12265 3383
rect 12299 3380 12311 3383
rect 12437 3383 12495 3389
rect 12437 3380 12449 3383
rect 12299 3352 12449 3380
rect 12299 3349 12311 3352
rect 12253 3343 12311 3349
rect 12437 3349 12449 3352
rect 12483 3349 12495 3383
rect 12437 3343 12495 3349
rect 13633 3383 13691 3389
rect 13633 3349 13645 3383
rect 13679 3380 13691 3383
rect 13814 3380 13820 3392
rect 13679 3352 13820 3380
rect 13679 3349 13691 3352
rect 13633 3343 13691 3349
rect 13814 3340 13820 3352
rect 13872 3340 13878 3392
rect 14182 3340 14188 3392
rect 14240 3380 14246 3392
rect 15194 3380 15200 3392
rect 14240 3352 15200 3380
rect 14240 3340 14246 3352
rect 15194 3340 15200 3352
rect 15252 3340 15258 3392
rect 15838 3340 15844 3392
rect 15896 3380 15902 3392
rect 16117 3383 16175 3389
rect 16117 3380 16129 3383
rect 15896 3352 16129 3380
rect 15896 3340 15902 3352
rect 16117 3349 16129 3352
rect 16163 3349 16175 3383
rect 16117 3343 16175 3349
rect 17402 3340 17408 3392
rect 17460 3380 17466 3392
rect 17865 3383 17923 3389
rect 17865 3380 17877 3383
rect 17460 3352 17877 3380
rect 17460 3340 17466 3352
rect 17865 3349 17877 3352
rect 17911 3349 17923 3383
rect 17972 3380 18000 3420
rect 18046 3408 18052 3460
rect 18104 3448 18110 3460
rect 18969 3451 19027 3457
rect 18969 3448 18981 3451
rect 18104 3420 18981 3448
rect 18104 3408 18110 3420
rect 18969 3417 18981 3420
rect 19015 3417 19027 3451
rect 18969 3411 19027 3417
rect 18417 3383 18475 3389
rect 18417 3380 18429 3383
rect 17972 3352 18429 3380
rect 17865 3343 17923 3349
rect 18417 3349 18429 3352
rect 18463 3349 18475 3383
rect 18417 3343 18475 3349
rect 18785 3383 18843 3389
rect 18785 3349 18797 3383
rect 18831 3380 18843 3383
rect 19306 3380 19334 3476
rect 20254 3408 20260 3460
rect 20312 3448 20318 3460
rect 20625 3451 20683 3457
rect 20625 3448 20637 3451
rect 20312 3420 20637 3448
rect 20312 3408 20318 3420
rect 20625 3417 20637 3420
rect 20671 3417 20683 3451
rect 20625 3411 20683 3417
rect 20993 3451 21051 3457
rect 20993 3417 21005 3451
rect 21039 3448 21051 3451
rect 21913 3451 21971 3457
rect 21913 3448 21925 3451
rect 21039 3420 21925 3448
rect 21039 3417 21051 3420
rect 20993 3411 21051 3417
rect 21913 3417 21925 3420
rect 21959 3417 21971 3451
rect 21913 3411 21971 3417
rect 18831 3352 19334 3380
rect 20073 3383 20131 3389
rect 18831 3349 18843 3352
rect 18785 3343 18843 3349
rect 20073 3349 20085 3383
rect 20119 3380 20131 3383
rect 20162 3380 20168 3392
rect 20119 3352 20168 3380
rect 20119 3349 20131 3352
rect 20073 3343 20131 3349
rect 20162 3340 20168 3352
rect 20220 3340 20226 3392
rect 20441 3383 20499 3389
rect 20441 3349 20453 3383
rect 20487 3380 20499 3383
rect 20530 3380 20536 3392
rect 20487 3352 20536 3380
rect 20487 3349 20499 3352
rect 20441 3343 20499 3349
rect 20530 3340 20536 3352
rect 20588 3380 20594 3392
rect 21008 3380 21036 3411
rect 20588 3352 21036 3380
rect 20588 3340 20594 3352
rect 21174 3340 21180 3392
rect 21232 3380 21238 3392
rect 21453 3383 21511 3389
rect 21453 3380 21465 3383
rect 21232 3352 21465 3380
rect 21232 3340 21238 3352
rect 21453 3349 21465 3352
rect 21499 3349 21511 3383
rect 21453 3343 21511 3349
rect 21726 3340 21732 3392
rect 21784 3380 21790 3392
rect 21821 3383 21879 3389
rect 21821 3380 21833 3383
rect 21784 3352 21833 3380
rect 21784 3340 21790 3352
rect 21821 3349 21833 3352
rect 21867 3349 21879 3383
rect 21821 3343 21879 3349
rect 22278 3340 22284 3392
rect 22336 3340 22342 3392
rect 22738 3340 22744 3392
rect 22796 3340 22802 3392
rect 552 3290 23368 3312
rect 552 3238 1366 3290
rect 1418 3238 1430 3290
rect 1482 3238 1494 3290
rect 1546 3238 1558 3290
rect 1610 3238 1622 3290
rect 1674 3238 1686 3290
rect 1738 3238 7366 3290
rect 7418 3238 7430 3290
rect 7482 3238 7494 3290
rect 7546 3238 7558 3290
rect 7610 3238 7622 3290
rect 7674 3238 7686 3290
rect 7738 3238 13366 3290
rect 13418 3238 13430 3290
rect 13482 3238 13494 3290
rect 13546 3238 13558 3290
rect 13610 3238 13622 3290
rect 13674 3238 13686 3290
rect 13738 3238 19366 3290
rect 19418 3238 19430 3290
rect 19482 3238 19494 3290
rect 19546 3238 19558 3290
rect 19610 3238 19622 3290
rect 19674 3238 19686 3290
rect 19738 3238 23368 3290
rect 552 3216 23368 3238
rect 2038 3176 2044 3188
rect 1320 3148 2044 3176
rect 1026 3000 1032 3052
rect 1084 3040 1090 3052
rect 1213 3043 1271 3049
rect 1213 3040 1225 3043
rect 1084 3012 1225 3040
rect 1084 3000 1090 3012
rect 1213 3009 1225 3012
rect 1259 3009 1271 3043
rect 1213 3003 1271 3009
rect 1320 2981 1348 3148
rect 2038 3136 2044 3148
rect 2096 3136 2102 3188
rect 5261 3179 5319 3185
rect 5261 3145 5273 3179
rect 5307 3176 5319 3179
rect 6730 3176 6736 3188
rect 5307 3148 6736 3176
rect 5307 3145 5319 3148
rect 5261 3139 5319 3145
rect 6730 3136 6736 3148
rect 6788 3136 6794 3188
rect 7009 3179 7067 3185
rect 7009 3145 7021 3179
rect 7055 3176 7067 3179
rect 7190 3176 7196 3188
rect 7055 3148 7196 3176
rect 7055 3145 7067 3148
rect 7009 3139 7067 3145
rect 7190 3136 7196 3148
rect 7248 3136 7254 3188
rect 8662 3136 8668 3188
rect 8720 3136 8726 3188
rect 9398 3136 9404 3188
rect 9456 3176 9462 3188
rect 10137 3179 10195 3185
rect 10137 3176 10149 3179
rect 9456 3148 10149 3176
rect 9456 3136 9462 3148
rect 10137 3145 10149 3148
rect 10183 3176 10195 3179
rect 10686 3176 10692 3188
rect 10183 3148 10692 3176
rect 10183 3145 10195 3148
rect 10137 3139 10195 3145
rect 10686 3136 10692 3148
rect 10744 3136 10750 3188
rect 10778 3136 10784 3188
rect 10836 3136 10842 3188
rect 11514 3136 11520 3188
rect 11572 3176 11578 3188
rect 11882 3176 11888 3188
rect 11572 3148 11888 3176
rect 11572 3136 11578 3148
rect 11882 3136 11888 3148
rect 11940 3176 11946 3188
rect 19797 3179 19855 3185
rect 19797 3176 19809 3179
rect 11940 3148 19809 3176
rect 11940 3136 11946 3148
rect 19797 3145 19809 3148
rect 19843 3145 19855 3179
rect 19797 3139 19855 3145
rect 1946 3108 1952 3120
rect 1872 3080 1952 3108
rect 1872 3049 1900 3080
rect 1946 3068 1952 3080
rect 2004 3068 2010 3120
rect 2317 3111 2375 3117
rect 2317 3077 2329 3111
rect 2363 3108 2375 3111
rect 3789 3111 3847 3117
rect 2363 3080 2774 3108
rect 2363 3077 2375 3080
rect 2317 3071 2375 3077
rect 1857 3043 1915 3049
rect 1857 3009 1869 3043
rect 1903 3009 1915 3043
rect 2746 3040 2774 3080
rect 3789 3077 3801 3111
rect 3835 3108 3847 3111
rect 3878 3108 3884 3120
rect 3835 3080 3884 3108
rect 3835 3077 3847 3080
rect 3789 3071 3847 3077
rect 3878 3068 3884 3080
rect 3936 3068 3942 3120
rect 4525 3111 4583 3117
rect 4525 3077 4537 3111
rect 4571 3108 4583 3111
rect 5537 3111 5595 3117
rect 4571 3080 5028 3108
rect 4571 3077 4583 3080
rect 4525 3071 4583 3077
rect 5000 3052 5028 3080
rect 5537 3077 5549 3111
rect 5583 3077 5595 3111
rect 5537 3071 5595 3077
rect 3329 3043 3387 3049
rect 3329 3040 3341 3043
rect 2746 3012 3341 3040
rect 1857 3003 1915 3009
rect 3329 3009 3341 3012
rect 3375 3009 3387 3043
rect 3329 3003 3387 3009
rect 4614 3000 4620 3052
rect 4672 3000 4678 3052
rect 4982 3000 4988 3052
rect 5040 3000 5046 3052
rect 1305 2975 1363 2981
rect 1305 2941 1317 2975
rect 1351 2941 1363 2975
rect 1949 2975 2007 2981
rect 1949 2972 1961 2975
rect 1305 2935 1363 2941
rect 1688 2944 1961 2972
rect 1688 2845 1716 2944
rect 1949 2941 1961 2944
rect 1995 2941 2007 2975
rect 1949 2935 2007 2941
rect 3142 2932 3148 2984
rect 3200 2972 3206 2984
rect 3421 2975 3479 2981
rect 3421 2972 3433 2975
rect 3200 2944 3433 2972
rect 3200 2932 3206 2944
rect 3421 2941 3433 2944
rect 3467 2941 3479 2975
rect 3421 2935 3479 2941
rect 4246 2932 4252 2984
rect 4304 2972 4310 2984
rect 4341 2975 4399 2981
rect 4341 2972 4353 2975
rect 4304 2944 4353 2972
rect 4304 2932 4310 2944
rect 4341 2941 4353 2944
rect 4387 2941 4399 2975
rect 4632 2972 4660 3000
rect 4893 2975 4951 2981
rect 4893 2972 4905 2975
rect 4632 2944 4905 2972
rect 4341 2935 4399 2941
rect 4893 2941 4905 2944
rect 4939 2941 4951 2975
rect 4893 2935 4951 2941
rect 5350 2932 5356 2984
rect 5408 2932 5414 2984
rect 5552 2972 5580 3071
rect 5994 3068 6000 3120
rect 6052 3068 6058 3120
rect 8680 3108 8708 3136
rect 8680 3080 8800 3108
rect 6012 3040 6040 3068
rect 6181 3043 6239 3049
rect 6181 3040 6193 3043
rect 6012 3012 6193 3040
rect 6181 3009 6193 3012
rect 6227 3040 6239 3043
rect 6822 3040 6828 3052
rect 6227 3012 6828 3040
rect 6227 3009 6239 3012
rect 6181 3003 6239 3009
rect 6822 3000 6828 3012
rect 6880 3000 6886 3052
rect 8294 3000 8300 3052
rect 8352 3040 8358 3052
rect 8772 3049 8800 3080
rect 9214 3068 9220 3120
rect 9272 3108 9278 3120
rect 9582 3108 9588 3120
rect 9272 3080 9444 3108
rect 9272 3068 9278 3080
rect 8665 3043 8723 3049
rect 8665 3040 8677 3043
rect 8352 3012 8677 3040
rect 8352 3000 8358 3012
rect 8665 3009 8677 3012
rect 8711 3009 8723 3043
rect 8665 3003 8723 3009
rect 8757 3043 8815 3049
rect 8757 3009 8769 3043
rect 8803 3009 8815 3043
rect 8757 3003 8815 3009
rect 8849 3043 8907 3049
rect 8849 3009 8861 3043
rect 8895 3040 8907 3043
rect 8895 3012 9260 3040
rect 8895 3009 8907 3012
rect 8849 3003 8907 3009
rect 5718 2972 5724 2984
rect 5552 2944 5724 2972
rect 5718 2932 5724 2944
rect 5776 2972 5782 2984
rect 5997 2975 6055 2981
rect 5997 2972 6009 2975
rect 5776 2944 6009 2972
rect 5776 2932 5782 2944
rect 5997 2941 6009 2944
rect 6043 2941 6055 2975
rect 5997 2935 6055 2941
rect 7193 2975 7251 2981
rect 7193 2941 7205 2975
rect 7239 2972 7251 2975
rect 7282 2972 7288 2984
rect 7239 2944 7288 2972
rect 7239 2941 7251 2944
rect 7193 2935 7251 2941
rect 7282 2932 7288 2944
rect 7340 2932 7346 2984
rect 7466 2932 7472 2984
rect 7524 2932 7530 2984
rect 8941 2975 8999 2981
rect 8941 2941 8953 2975
rect 8987 2941 8999 2975
rect 9232 2972 9260 3012
rect 9306 3000 9312 3052
rect 9364 3000 9370 3052
rect 9416 3049 9444 3080
rect 9508 3080 9588 3108
rect 9508 3049 9536 3080
rect 9582 3068 9588 3080
rect 9640 3068 9646 3120
rect 12526 3068 12532 3120
rect 12584 3108 12590 3120
rect 12805 3111 12863 3117
rect 12805 3108 12817 3111
rect 12584 3080 12817 3108
rect 12584 3068 12590 3080
rect 12805 3077 12817 3080
rect 12851 3077 12863 3111
rect 12805 3071 12863 3077
rect 13446 3068 13452 3120
rect 13504 3108 13510 3120
rect 13541 3111 13599 3117
rect 13541 3108 13553 3111
rect 13504 3080 13553 3108
rect 13504 3068 13510 3080
rect 13541 3077 13553 3080
rect 13587 3077 13599 3111
rect 13541 3071 13599 3077
rect 15194 3068 15200 3120
rect 15252 3108 15258 3120
rect 17126 3108 17132 3120
rect 15252 3080 17132 3108
rect 15252 3068 15258 3080
rect 17126 3068 17132 3080
rect 17184 3068 17190 3120
rect 17310 3068 17316 3120
rect 17368 3068 17374 3120
rect 17402 3068 17408 3120
rect 17460 3068 17466 3120
rect 17770 3068 17776 3120
rect 17828 3068 17834 3120
rect 19812 3108 19840 3139
rect 19886 3136 19892 3188
rect 19944 3176 19950 3188
rect 20438 3176 20444 3188
rect 19944 3148 20444 3176
rect 19944 3136 19950 3148
rect 20438 3136 20444 3148
rect 20496 3136 20502 3188
rect 20530 3136 20536 3188
rect 20588 3176 20594 3188
rect 21085 3179 21143 3185
rect 21085 3176 21097 3179
rect 20588 3148 21097 3176
rect 20588 3136 20594 3148
rect 21085 3145 21097 3148
rect 21131 3145 21143 3179
rect 21085 3139 21143 3145
rect 19812 3080 21312 3108
rect 9401 3043 9459 3049
rect 9401 3009 9413 3043
rect 9447 3009 9459 3043
rect 9401 3003 9459 3009
rect 9493 3043 9551 3049
rect 9493 3009 9505 3043
rect 9539 3009 9551 3043
rect 10226 3040 10232 3052
rect 9493 3003 9551 3009
rect 9968 3012 10232 3040
rect 9508 2972 9536 3003
rect 9232 2944 9536 2972
rect 8941 2935 8999 2941
rect 8956 2904 8984 2935
rect 9582 2932 9588 2984
rect 9640 2932 9646 2984
rect 9968 2981 9996 3012
rect 10226 3000 10232 3012
rect 10284 3000 10290 3052
rect 10620 3012 11376 3040
rect 9953 2975 10011 2981
rect 9953 2941 9965 2975
rect 9999 2941 10011 2975
rect 9953 2935 10011 2941
rect 10134 2932 10140 2984
rect 10192 2932 10198 2984
rect 10620 2981 10648 3012
rect 11348 2984 11376 3012
rect 11790 3000 11796 3052
rect 11848 3040 11854 3052
rect 12250 3040 12256 3052
rect 11848 3012 12256 3040
rect 11848 3000 11854 3012
rect 12250 3000 12256 3012
rect 12308 3000 12314 3052
rect 19794 3040 19800 3052
rect 13740 3012 18000 3040
rect 13740 2984 13768 3012
rect 10597 2975 10655 2981
rect 10597 2941 10609 2975
rect 10643 2941 10655 2975
rect 10597 2935 10655 2941
rect 10689 2975 10747 2981
rect 10689 2941 10701 2975
rect 10735 2972 10747 2975
rect 10778 2972 10784 2984
rect 10735 2944 10784 2972
rect 10735 2941 10747 2944
rect 10689 2935 10747 2941
rect 10778 2932 10784 2944
rect 10836 2932 10842 2984
rect 10873 2975 10931 2981
rect 10873 2941 10885 2975
rect 10919 2972 10931 2975
rect 11054 2972 11060 2984
rect 10919 2944 11060 2972
rect 10919 2941 10931 2944
rect 10873 2935 10931 2941
rect 11054 2932 11060 2944
rect 11112 2932 11118 2984
rect 11149 2975 11207 2981
rect 11149 2941 11161 2975
rect 11195 2972 11207 2975
rect 11238 2972 11244 2984
rect 11195 2944 11244 2972
rect 11195 2941 11207 2944
rect 11149 2935 11207 2941
rect 11238 2932 11244 2944
rect 11296 2932 11302 2984
rect 11330 2932 11336 2984
rect 11388 2932 11394 2984
rect 11514 2932 11520 2984
rect 11572 2932 11578 2984
rect 11606 2932 11612 2984
rect 11664 2932 11670 2984
rect 12069 2975 12127 2981
rect 12069 2941 12081 2975
rect 12115 2941 12127 2975
rect 12069 2935 12127 2941
rect 12529 2975 12587 2981
rect 12529 2941 12541 2975
rect 12575 2972 12587 2975
rect 12894 2972 12900 2984
rect 12575 2944 12900 2972
rect 12575 2941 12587 2944
rect 12529 2935 12587 2941
rect 9600 2904 9628 2932
rect 8956 2876 9628 2904
rect 12084 2904 12112 2935
rect 12894 2932 12900 2944
rect 12952 2932 12958 2984
rect 13722 2932 13728 2984
rect 13780 2932 13786 2984
rect 13817 2975 13875 2981
rect 13817 2941 13829 2975
rect 13863 2972 13875 2975
rect 14001 2975 14059 2981
rect 14001 2972 14013 2975
rect 13863 2944 14013 2972
rect 13863 2941 13875 2944
rect 13817 2935 13875 2941
rect 14001 2941 14013 2944
rect 14047 2941 14059 2975
rect 14001 2935 14059 2941
rect 14090 2932 14096 2984
rect 14148 2932 14154 2984
rect 14458 2932 14464 2984
rect 14516 2972 14522 2984
rect 15105 2975 15163 2981
rect 15105 2972 15117 2975
rect 14516 2944 15117 2972
rect 14516 2932 14522 2944
rect 15105 2941 15117 2944
rect 15151 2941 15163 2975
rect 15105 2935 15163 2941
rect 16485 2975 16543 2981
rect 16485 2941 16497 2975
rect 16531 2972 16543 2975
rect 16666 2972 16672 2984
rect 16531 2944 16672 2972
rect 16531 2941 16543 2944
rect 16485 2935 16543 2941
rect 16666 2932 16672 2944
rect 16724 2972 16730 2984
rect 17221 2975 17279 2981
rect 17221 2972 17233 2975
rect 16724 2944 17233 2972
rect 16724 2932 16730 2944
rect 17221 2941 17233 2944
rect 17267 2972 17279 2975
rect 17402 2972 17408 2984
rect 17267 2944 17408 2972
rect 17267 2941 17279 2944
rect 17221 2935 17279 2941
rect 17402 2932 17408 2944
rect 17460 2932 17466 2984
rect 17497 2975 17555 2981
rect 17497 2941 17509 2975
rect 17543 2941 17555 2975
rect 17497 2935 17555 2941
rect 12342 2904 12348 2916
rect 12084 2876 12348 2904
rect 12342 2864 12348 2876
rect 12400 2904 12406 2916
rect 12805 2907 12863 2913
rect 12400 2876 12756 2904
rect 12400 2864 12406 2876
rect 1673 2839 1731 2845
rect 1673 2805 1685 2839
rect 1719 2805 1731 2839
rect 1673 2799 1731 2805
rect 4157 2839 4215 2845
rect 4157 2805 4169 2839
rect 4203 2836 4215 2839
rect 4246 2836 4252 2848
rect 4203 2808 4252 2836
rect 4203 2805 4215 2808
rect 4157 2799 4215 2805
rect 4246 2796 4252 2808
rect 4304 2796 4310 2848
rect 5810 2796 5816 2848
rect 5868 2796 5874 2848
rect 7282 2796 7288 2848
rect 7340 2836 7346 2848
rect 7377 2839 7435 2845
rect 7377 2836 7389 2839
rect 7340 2808 7389 2836
rect 7340 2796 7346 2808
rect 7377 2805 7389 2808
rect 7423 2805 7435 2839
rect 7377 2799 7435 2805
rect 8478 2796 8484 2848
rect 8536 2796 8542 2848
rect 9122 2796 9128 2848
rect 9180 2796 9186 2848
rect 10505 2839 10563 2845
rect 10505 2805 10517 2839
rect 10551 2836 10563 2839
rect 11514 2836 11520 2848
rect 10551 2808 11520 2836
rect 10551 2805 10563 2808
rect 10505 2799 10563 2805
rect 11514 2796 11520 2808
rect 11572 2796 11578 2848
rect 11885 2839 11943 2845
rect 11885 2805 11897 2839
rect 11931 2836 11943 2839
rect 12066 2836 12072 2848
rect 11931 2808 12072 2836
rect 11931 2805 11943 2808
rect 11885 2799 11943 2805
rect 12066 2796 12072 2808
rect 12124 2796 12130 2848
rect 12618 2796 12624 2848
rect 12676 2796 12682 2848
rect 12728 2836 12756 2876
rect 12805 2873 12817 2907
rect 12851 2904 12863 2907
rect 13538 2904 13544 2916
rect 12851 2876 13544 2904
rect 12851 2873 12863 2876
rect 12805 2867 12863 2873
rect 13538 2864 13544 2876
rect 13596 2864 13602 2916
rect 17524 2904 17552 2935
rect 17586 2932 17592 2984
rect 17644 2972 17650 2984
rect 17972 2981 18000 3012
rect 19168 3012 19800 3040
rect 17957 2975 18015 2981
rect 17644 2944 17908 2972
rect 17644 2932 17650 2944
rect 13648 2876 17552 2904
rect 17773 2907 17831 2913
rect 13648 2836 13676 2876
rect 17773 2873 17785 2907
rect 17819 2873 17831 2907
rect 17880 2904 17908 2944
rect 17957 2941 17969 2975
rect 18003 2941 18015 2975
rect 17957 2935 18015 2941
rect 18049 2975 18107 2981
rect 18049 2941 18061 2975
rect 18095 2972 18107 2975
rect 18598 2972 18604 2984
rect 18095 2944 18604 2972
rect 18095 2941 18107 2944
rect 18049 2935 18107 2941
rect 18598 2932 18604 2944
rect 18656 2932 18662 2984
rect 19168 2981 19196 3012
rect 19794 3000 19800 3012
rect 19852 3000 19858 3052
rect 19904 3012 20483 3040
rect 19153 2975 19211 2981
rect 19153 2941 19165 2975
rect 19199 2941 19211 2975
rect 19153 2935 19211 2941
rect 19337 2975 19395 2981
rect 19337 2941 19349 2975
rect 19383 2972 19395 2975
rect 19904 2972 19932 3012
rect 19383 2944 19932 2972
rect 19383 2941 19395 2944
rect 19337 2935 19395 2941
rect 19978 2932 19984 2984
rect 20036 2932 20042 2984
rect 20349 2975 20407 2981
rect 20349 2941 20361 2975
rect 20395 2941 20407 2975
rect 20455 2972 20483 3012
rect 20622 3000 20628 3052
rect 20680 3000 20686 3052
rect 20990 3000 20996 3052
rect 21048 3040 21054 3052
rect 21177 3043 21235 3049
rect 21177 3040 21189 3043
rect 21048 3012 21189 3040
rect 21048 3000 21054 3012
rect 21177 3009 21189 3012
rect 21223 3009 21235 3043
rect 21284 3040 21312 3080
rect 21910 3068 21916 3120
rect 21968 3108 21974 3120
rect 22189 3111 22247 3117
rect 22189 3108 22201 3111
rect 21968 3080 22201 3108
rect 21968 3068 21974 3080
rect 22189 3077 22201 3080
rect 22235 3077 22247 3111
rect 22189 3071 22247 3077
rect 22465 3111 22523 3117
rect 22465 3077 22477 3111
rect 22511 3108 22523 3111
rect 23566 3108 23572 3120
rect 22511 3080 23572 3108
rect 22511 3077 22523 3080
rect 22465 3071 22523 3077
rect 23566 3068 23572 3080
rect 23624 3068 23630 3120
rect 22002 3040 22008 3052
rect 21284 3012 21404 3040
rect 21177 3003 21235 3009
rect 20640 2972 20668 3000
rect 20898 2972 20904 2984
rect 20455 2944 20668 2972
rect 20732 2944 20904 2972
rect 20349 2935 20407 2941
rect 19245 2907 19303 2913
rect 19245 2904 19257 2907
rect 17880 2876 19257 2904
rect 17773 2867 17831 2873
rect 19245 2873 19257 2876
rect 19291 2873 19303 2907
rect 20364 2904 20392 2935
rect 20732 2904 20760 2944
rect 20898 2932 20904 2944
rect 20956 2932 20962 2984
rect 21266 2932 21272 2984
rect 21324 2932 21330 2984
rect 21376 2981 21404 3012
rect 21560 3012 22008 3040
rect 21560 2981 21588 3012
rect 22002 3000 22008 3012
rect 22060 3040 22066 3052
rect 22830 3040 22836 3052
rect 22060 3012 22140 3040
rect 22060 3000 22066 3012
rect 21361 2975 21419 2981
rect 21361 2941 21373 2975
rect 21407 2941 21419 2975
rect 21361 2935 21419 2941
rect 21545 2975 21603 2981
rect 21545 2941 21557 2975
rect 21591 2941 21603 2975
rect 21545 2935 21603 2941
rect 21818 2932 21824 2984
rect 21876 2932 21882 2984
rect 22112 2981 22140 3012
rect 22664 3012 22836 3040
rect 22664 2981 22692 3012
rect 22830 3000 22836 3012
rect 22888 3000 22894 3052
rect 22097 2975 22155 2981
rect 22097 2941 22109 2975
rect 22143 2941 22155 2975
rect 22097 2935 22155 2941
rect 22649 2975 22707 2981
rect 22649 2941 22661 2975
rect 22695 2941 22707 2975
rect 22649 2935 22707 2941
rect 22738 2932 22744 2984
rect 22796 2932 22802 2984
rect 20364 2876 20760 2904
rect 19245 2867 19303 2873
rect 12728 2808 13676 2836
rect 15010 2796 15016 2848
rect 15068 2796 15074 2848
rect 16206 2796 16212 2848
rect 16264 2836 16270 2848
rect 16393 2839 16451 2845
rect 16393 2836 16405 2839
rect 16264 2808 16405 2836
rect 16264 2796 16270 2808
rect 16393 2805 16405 2808
rect 16439 2805 16451 2839
rect 16393 2799 16451 2805
rect 16758 2796 16764 2848
rect 16816 2836 16822 2848
rect 17037 2839 17095 2845
rect 17037 2836 17049 2839
rect 16816 2808 17049 2836
rect 16816 2796 16822 2808
rect 17037 2805 17049 2808
rect 17083 2805 17095 2839
rect 17037 2799 17095 2805
rect 17126 2796 17132 2848
rect 17184 2836 17190 2848
rect 17788 2836 17816 2867
rect 20806 2864 20812 2916
rect 20864 2904 20870 2916
rect 21836 2904 21864 2932
rect 23290 2904 23296 2916
rect 20864 2876 21864 2904
rect 22020 2876 23296 2904
rect 20864 2864 20870 2876
rect 19886 2836 19892 2848
rect 17184 2808 19892 2836
rect 17184 2796 17190 2808
rect 19886 2796 19892 2808
rect 19944 2796 19950 2848
rect 19978 2796 19984 2848
rect 20036 2836 20042 2848
rect 20165 2839 20223 2845
rect 20165 2836 20177 2839
rect 20036 2808 20177 2836
rect 20036 2796 20042 2808
rect 20165 2805 20177 2808
rect 20211 2805 20223 2839
rect 20165 2799 20223 2805
rect 20717 2839 20775 2845
rect 20717 2805 20729 2839
rect 20763 2836 20775 2839
rect 20898 2836 20904 2848
rect 20763 2808 20904 2836
rect 20763 2805 20775 2808
rect 20717 2799 20775 2805
rect 20898 2796 20904 2808
rect 20956 2796 20962 2848
rect 21450 2796 21456 2848
rect 21508 2836 21514 2848
rect 21729 2839 21787 2845
rect 21729 2836 21741 2839
rect 21508 2808 21741 2836
rect 21508 2796 21514 2808
rect 21729 2805 21741 2808
rect 21775 2805 21787 2839
rect 21729 2799 21787 2805
rect 21818 2796 21824 2848
rect 21876 2836 21882 2848
rect 22020 2845 22048 2876
rect 23290 2864 23296 2876
rect 23348 2864 23354 2916
rect 22005 2839 22063 2845
rect 22005 2836 22017 2839
rect 21876 2808 22017 2836
rect 21876 2796 21882 2808
rect 22005 2805 22017 2808
rect 22051 2805 22063 2839
rect 22005 2799 22063 2805
rect 22830 2796 22836 2848
rect 22888 2836 22894 2848
rect 22925 2839 22983 2845
rect 22925 2836 22937 2839
rect 22888 2808 22937 2836
rect 22888 2796 22894 2808
rect 22925 2805 22937 2808
rect 22971 2805 22983 2839
rect 22925 2799 22983 2805
rect 552 2746 23368 2768
rect 552 2694 4366 2746
rect 4418 2694 4430 2746
rect 4482 2694 4494 2746
rect 4546 2694 4558 2746
rect 4610 2694 4622 2746
rect 4674 2694 4686 2746
rect 4738 2694 10366 2746
rect 10418 2694 10430 2746
rect 10482 2694 10494 2746
rect 10546 2694 10558 2746
rect 10610 2694 10622 2746
rect 10674 2694 10686 2746
rect 10738 2694 16366 2746
rect 16418 2694 16430 2746
rect 16482 2694 16494 2746
rect 16546 2694 16558 2746
rect 16610 2694 16622 2746
rect 16674 2694 16686 2746
rect 16738 2694 22366 2746
rect 22418 2694 22430 2746
rect 22482 2694 22494 2746
rect 22546 2694 22558 2746
rect 22610 2694 22622 2746
rect 22674 2694 22686 2746
rect 22738 2694 23368 2746
rect 552 2672 23368 2694
rect 2961 2635 3019 2641
rect 2961 2601 2973 2635
rect 3007 2632 3019 2635
rect 4801 2635 4859 2641
rect 3007 2604 4476 2632
rect 3007 2601 3019 2604
rect 2961 2595 3019 2601
rect 3326 2564 3332 2576
rect 2884 2536 3332 2564
rect 2884 2505 2912 2536
rect 3326 2524 3332 2536
rect 3384 2564 3390 2576
rect 3384 2536 3740 2564
rect 3384 2524 3390 2536
rect 2869 2499 2927 2505
rect 2869 2465 2881 2499
rect 2915 2465 2927 2499
rect 2869 2459 2927 2465
rect 3145 2499 3203 2505
rect 3145 2465 3157 2499
rect 3191 2496 3203 2499
rect 3191 2468 3280 2496
rect 3191 2465 3203 2468
rect 3145 2459 3203 2465
rect 3142 2320 3148 2372
rect 3200 2320 3206 2372
rect 3252 2301 3280 2468
rect 3418 2456 3424 2508
rect 3476 2456 3482 2508
rect 3712 2505 3740 2536
rect 4448 2505 4476 2604
rect 4801 2601 4813 2635
rect 4847 2632 4859 2635
rect 5074 2632 5080 2644
rect 4847 2604 5080 2632
rect 4847 2601 4859 2604
rect 4801 2595 4859 2601
rect 5074 2592 5080 2604
rect 5132 2592 5138 2644
rect 5534 2592 5540 2644
rect 5592 2592 5598 2644
rect 5718 2592 5724 2644
rect 5776 2632 5782 2644
rect 5776 2604 6316 2632
rect 5776 2592 5782 2604
rect 5552 2564 5580 2592
rect 6288 2564 6316 2604
rect 6546 2592 6552 2644
rect 6604 2592 6610 2644
rect 7466 2592 7472 2644
rect 7524 2632 7530 2644
rect 7561 2635 7619 2641
rect 7561 2632 7573 2635
rect 7524 2604 7573 2632
rect 7524 2592 7530 2604
rect 7561 2601 7573 2604
rect 7607 2601 7619 2635
rect 7561 2595 7619 2601
rect 8021 2635 8079 2641
rect 8021 2601 8033 2635
rect 8067 2632 8079 2635
rect 8389 2635 8447 2641
rect 8389 2632 8401 2635
rect 8067 2604 8401 2632
rect 8067 2601 8079 2604
rect 8021 2595 8079 2601
rect 8389 2601 8401 2604
rect 8435 2632 8447 2635
rect 8849 2635 8907 2641
rect 8849 2632 8861 2635
rect 8435 2604 8861 2632
rect 8435 2601 8447 2604
rect 8389 2595 8447 2601
rect 8849 2601 8861 2604
rect 8895 2632 8907 2635
rect 10778 2632 10784 2644
rect 8895 2604 10784 2632
rect 8895 2601 8907 2604
rect 8849 2595 8907 2601
rect 10778 2592 10784 2604
rect 10836 2592 10842 2644
rect 11149 2635 11207 2641
rect 11149 2601 11161 2635
rect 11195 2632 11207 2635
rect 11330 2632 11336 2644
rect 11195 2604 11336 2632
rect 11195 2601 11207 2604
rect 11149 2595 11207 2601
rect 11330 2592 11336 2604
rect 11388 2592 11394 2644
rect 11514 2592 11520 2644
rect 11572 2632 11578 2644
rect 11698 2632 11704 2644
rect 11572 2604 11704 2632
rect 11572 2592 11578 2604
rect 11698 2592 11704 2604
rect 11756 2592 11762 2644
rect 11790 2592 11796 2644
rect 11848 2592 11854 2644
rect 11882 2592 11888 2644
rect 11940 2592 11946 2644
rect 12253 2635 12311 2641
rect 12253 2632 12265 2635
rect 11992 2604 12265 2632
rect 6641 2567 6699 2573
rect 6641 2564 6653 2567
rect 5552 2536 6132 2564
rect 6288 2536 6653 2564
rect 3697 2499 3755 2505
rect 3697 2465 3709 2499
rect 3743 2465 3755 2499
rect 3697 2459 3755 2465
rect 4433 2499 4491 2505
rect 4433 2465 4445 2499
rect 4479 2496 4491 2499
rect 5169 2499 5227 2505
rect 5169 2496 5181 2499
rect 4479 2468 5181 2496
rect 4479 2465 4491 2468
rect 4433 2459 4491 2465
rect 5169 2465 5181 2468
rect 5215 2465 5227 2499
rect 5169 2459 5227 2465
rect 5353 2499 5411 2505
rect 5353 2465 5365 2499
rect 5399 2465 5411 2499
rect 5353 2459 5411 2465
rect 5629 2499 5687 2505
rect 5629 2465 5641 2499
rect 5675 2496 5687 2499
rect 5994 2496 6000 2508
rect 5675 2468 6000 2496
rect 5675 2465 5687 2468
rect 5629 2459 5687 2465
rect 3605 2431 3663 2437
rect 3605 2397 3617 2431
rect 3651 2428 3663 2431
rect 3878 2428 3884 2440
rect 3651 2400 3884 2428
rect 3651 2397 3663 2400
rect 3605 2391 3663 2397
rect 3878 2388 3884 2400
rect 3936 2388 3942 2440
rect 4157 2431 4215 2437
rect 4157 2397 4169 2431
rect 4203 2428 4215 2431
rect 4341 2431 4399 2437
rect 4341 2428 4353 2431
rect 4203 2400 4353 2428
rect 4203 2397 4215 2400
rect 4157 2391 4215 2397
rect 4341 2397 4353 2400
rect 4387 2397 4399 2431
rect 5368 2428 5396 2459
rect 5994 2456 6000 2468
rect 6052 2456 6058 2508
rect 6104 2494 6132 2536
rect 6641 2533 6653 2536
rect 6687 2533 6699 2567
rect 6641 2527 6699 2533
rect 6822 2524 6828 2576
rect 6880 2524 6886 2576
rect 9122 2564 9128 2576
rect 8128 2536 9128 2564
rect 6181 2499 6239 2505
rect 6181 2494 6193 2499
rect 6104 2466 6193 2494
rect 6181 2465 6193 2466
rect 6227 2465 6239 2499
rect 6181 2459 6239 2465
rect 6730 2456 6736 2508
rect 6788 2496 6794 2508
rect 7193 2499 7251 2505
rect 7193 2496 7205 2499
rect 6788 2468 7205 2496
rect 6788 2456 6794 2468
rect 7193 2465 7205 2468
rect 7239 2465 7251 2499
rect 7193 2459 7251 2465
rect 7377 2499 7435 2505
rect 7377 2465 7389 2499
rect 7423 2496 7435 2499
rect 7742 2496 7748 2508
rect 7423 2468 7748 2496
rect 7423 2465 7435 2468
rect 7377 2459 7435 2465
rect 7742 2456 7748 2468
rect 7800 2456 7806 2508
rect 8128 2505 8156 2536
rect 9122 2524 9128 2536
rect 9180 2524 9186 2576
rect 9401 2567 9459 2573
rect 9401 2533 9413 2567
rect 9447 2564 9459 2567
rect 9582 2564 9588 2576
rect 9447 2536 9588 2564
rect 9447 2533 9459 2536
rect 9401 2527 9459 2533
rect 9582 2524 9588 2536
rect 9640 2524 9646 2576
rect 9674 2524 9680 2576
rect 9732 2564 9738 2576
rect 10597 2567 10655 2573
rect 9732 2536 10364 2564
rect 9732 2524 9738 2536
rect 7837 2499 7895 2505
rect 7837 2465 7849 2499
rect 7883 2465 7895 2499
rect 7837 2459 7895 2465
rect 8113 2499 8171 2505
rect 8113 2465 8125 2499
rect 8159 2465 8171 2499
rect 8113 2459 8171 2465
rect 8205 2499 8263 2505
rect 8205 2465 8217 2499
rect 8251 2465 8263 2499
rect 8205 2459 8263 2465
rect 5810 2428 5816 2440
rect 5368 2400 5816 2428
rect 4341 2391 4399 2397
rect 5810 2388 5816 2400
rect 5868 2388 5874 2440
rect 6089 2431 6147 2437
rect 6089 2397 6101 2431
rect 6135 2397 6147 2431
rect 6089 2391 6147 2397
rect 6104 2360 6132 2391
rect 7006 2388 7012 2440
rect 7064 2388 7070 2440
rect 7098 2388 7104 2440
rect 7156 2388 7162 2440
rect 7852 2428 7880 2459
rect 8220 2428 8248 2459
rect 8478 2456 8484 2508
rect 8536 2456 8542 2508
rect 8754 2456 8760 2508
rect 8812 2456 8818 2508
rect 9033 2499 9091 2505
rect 9033 2465 9045 2499
rect 9079 2496 9091 2499
rect 9217 2499 9275 2505
rect 9217 2496 9229 2499
rect 9079 2468 9229 2496
rect 9079 2465 9091 2468
rect 9033 2459 9091 2465
rect 9217 2465 9229 2468
rect 9263 2465 9275 2499
rect 9217 2459 9275 2465
rect 8938 2428 8944 2440
rect 7852 2400 8944 2428
rect 8938 2388 8944 2400
rect 8996 2388 9002 2440
rect 9232 2428 9260 2459
rect 9490 2456 9496 2508
rect 9548 2456 9554 2508
rect 9769 2499 9827 2505
rect 9769 2465 9781 2499
rect 9815 2496 9827 2499
rect 9815 2468 9996 2496
rect 9815 2465 9827 2468
rect 9769 2459 9827 2465
rect 9968 2428 9996 2468
rect 10042 2456 10048 2508
rect 10100 2456 10106 2508
rect 10336 2505 10364 2536
rect 10597 2533 10609 2567
rect 10643 2564 10655 2567
rect 11808 2564 11836 2592
rect 10643 2536 11100 2564
rect 10643 2533 10655 2536
rect 10597 2527 10655 2533
rect 10229 2499 10287 2505
rect 10229 2465 10241 2499
rect 10275 2465 10287 2499
rect 10229 2459 10287 2465
rect 10321 2499 10379 2505
rect 10321 2465 10333 2499
rect 10367 2465 10379 2499
rect 10321 2459 10379 2465
rect 9232 2400 9996 2428
rect 6178 2360 6184 2372
rect 6104 2332 6184 2360
rect 6178 2320 6184 2332
rect 6236 2320 6242 2372
rect 8294 2360 8300 2372
rect 7760 2332 8300 2360
rect 3237 2295 3295 2301
rect 3237 2261 3249 2295
rect 3283 2292 3295 2295
rect 3789 2295 3847 2301
rect 3789 2292 3801 2295
rect 3283 2264 3801 2292
rect 3283 2261 3295 2264
rect 3237 2255 3295 2261
rect 3789 2261 3801 2264
rect 3835 2261 3847 2295
rect 3789 2255 3847 2261
rect 3970 2252 3976 2304
rect 4028 2292 4034 2304
rect 7760 2292 7788 2332
rect 8294 2320 8300 2332
rect 8352 2320 8358 2372
rect 9217 2363 9275 2369
rect 9217 2329 9229 2363
rect 9263 2360 9275 2363
rect 9766 2360 9772 2372
rect 9263 2332 9772 2360
rect 9263 2329 9275 2332
rect 9217 2323 9275 2329
rect 9766 2320 9772 2332
rect 9824 2320 9830 2372
rect 4028 2264 7788 2292
rect 4028 2252 4034 2264
rect 7834 2252 7840 2304
rect 7892 2252 7898 2304
rect 8110 2252 8116 2304
rect 8168 2292 8174 2304
rect 8205 2295 8263 2301
rect 8205 2292 8217 2295
rect 8168 2264 8217 2292
rect 8168 2252 8174 2264
rect 8205 2261 8217 2264
rect 8251 2292 8263 2295
rect 8754 2292 8760 2304
rect 8251 2264 8760 2292
rect 8251 2261 8263 2264
rect 8205 2255 8263 2261
rect 8754 2252 8760 2264
rect 8812 2252 8818 2304
rect 9033 2295 9091 2301
rect 9033 2261 9045 2295
rect 9079 2292 9091 2295
rect 9122 2292 9128 2304
rect 9079 2264 9128 2292
rect 9079 2261 9091 2264
rect 9033 2255 9091 2261
rect 9122 2252 9128 2264
rect 9180 2252 9186 2304
rect 9398 2252 9404 2304
rect 9456 2292 9462 2304
rect 9585 2295 9643 2301
rect 9585 2292 9597 2295
rect 9456 2264 9597 2292
rect 9456 2252 9462 2264
rect 9585 2261 9597 2264
rect 9631 2261 9643 2295
rect 9968 2292 9996 2400
rect 10244 2360 10272 2459
rect 10410 2456 10416 2508
rect 10468 2456 10474 2508
rect 10962 2456 10968 2508
rect 11020 2456 11026 2508
rect 11072 2428 11100 2536
rect 11624 2536 11836 2564
rect 11624 2505 11652 2536
rect 11333 2499 11391 2505
rect 11333 2465 11345 2499
rect 11379 2465 11391 2499
rect 11333 2459 11391 2465
rect 11609 2499 11667 2505
rect 11609 2465 11621 2499
rect 11655 2465 11667 2499
rect 11609 2459 11667 2465
rect 11238 2428 11244 2440
rect 11072 2400 11244 2428
rect 11238 2388 11244 2400
rect 11296 2388 11302 2440
rect 11348 2428 11376 2459
rect 11698 2456 11704 2508
rect 11756 2456 11762 2508
rect 11793 2499 11851 2505
rect 11793 2465 11805 2499
rect 11839 2496 11851 2499
rect 11900 2496 11928 2592
rect 11992 2573 12020 2604
rect 12253 2601 12265 2604
rect 12299 2632 12311 2635
rect 12342 2632 12348 2644
rect 12299 2604 12348 2632
rect 12299 2601 12311 2604
rect 12253 2595 12311 2601
rect 12342 2592 12348 2604
rect 12400 2592 12406 2644
rect 13265 2635 13323 2641
rect 13265 2601 13277 2635
rect 13311 2632 13323 2635
rect 13538 2632 13544 2644
rect 13311 2604 13544 2632
rect 13311 2601 13323 2604
rect 13265 2595 13323 2601
rect 13538 2592 13544 2604
rect 13596 2632 13602 2644
rect 13596 2604 15148 2632
rect 13596 2592 13602 2604
rect 11977 2567 12035 2573
rect 11977 2533 11989 2567
rect 12023 2533 12035 2567
rect 11977 2527 12035 2533
rect 12434 2524 12440 2576
rect 12492 2524 12498 2576
rect 14737 2567 14795 2573
rect 14737 2533 14749 2567
rect 14783 2564 14795 2567
rect 15120 2564 15148 2604
rect 16574 2592 16580 2644
rect 16632 2632 16638 2644
rect 19061 2635 19119 2641
rect 19061 2632 19073 2635
rect 16632 2604 19073 2632
rect 16632 2592 16638 2604
rect 19061 2601 19073 2604
rect 19107 2632 19119 2635
rect 19107 2604 22324 2632
rect 19107 2601 19119 2604
rect 19061 2595 19119 2601
rect 15289 2567 15347 2573
rect 15289 2564 15301 2567
rect 14783 2536 15056 2564
rect 15120 2536 15301 2564
rect 14783 2533 14795 2536
rect 14737 2527 14795 2533
rect 15028 2508 15056 2536
rect 15289 2533 15301 2536
rect 15335 2564 15347 2567
rect 16117 2567 16175 2573
rect 16117 2564 16129 2567
rect 15335 2536 16129 2564
rect 15335 2533 15347 2536
rect 15289 2527 15347 2533
rect 16117 2533 16129 2536
rect 16163 2533 16175 2567
rect 16117 2527 16175 2533
rect 16206 2524 16212 2576
rect 16264 2564 16270 2576
rect 16850 2564 16856 2576
rect 16264 2536 16436 2564
rect 16264 2524 16270 2536
rect 11839 2468 11928 2496
rect 12069 2499 12127 2505
rect 11839 2465 11851 2468
rect 11793 2459 11851 2465
rect 12069 2465 12081 2499
rect 12115 2494 12127 2499
rect 12158 2494 12164 2508
rect 12115 2466 12164 2494
rect 12115 2465 12127 2466
rect 12069 2459 12127 2465
rect 12158 2456 12164 2466
rect 12216 2456 12222 2508
rect 12250 2456 12256 2508
rect 12308 2496 12314 2508
rect 12345 2499 12403 2505
rect 12345 2496 12357 2499
rect 12308 2468 12357 2496
rect 12308 2456 12314 2468
rect 12345 2465 12357 2468
rect 12391 2465 12403 2499
rect 12345 2459 12403 2465
rect 12526 2456 12532 2508
rect 12584 2496 12590 2508
rect 12621 2499 12679 2505
rect 12621 2496 12633 2499
rect 12584 2468 12633 2496
rect 12584 2456 12590 2468
rect 12621 2465 12633 2468
rect 12667 2465 12679 2499
rect 12621 2459 12679 2465
rect 12894 2456 12900 2508
rect 12952 2456 12958 2508
rect 12989 2499 13047 2505
rect 12989 2465 13001 2499
rect 13035 2496 13047 2499
rect 13078 2496 13084 2508
rect 13035 2468 13084 2496
rect 13035 2465 13047 2468
rect 12989 2459 13047 2465
rect 13078 2456 13084 2468
rect 13136 2456 13142 2508
rect 13449 2499 13507 2505
rect 13449 2496 13461 2499
rect 13188 2468 13461 2496
rect 11348 2400 12112 2428
rect 11348 2360 11376 2400
rect 10244 2332 11376 2360
rect 11422 2320 11428 2372
rect 11480 2360 11486 2372
rect 11977 2363 12035 2369
rect 11977 2360 11989 2363
rect 11480 2332 11989 2360
rect 11480 2320 11486 2332
rect 11977 2329 11989 2332
rect 12023 2329 12035 2363
rect 11977 2323 12035 2329
rect 10597 2295 10655 2301
rect 10597 2292 10609 2295
rect 9968 2264 10609 2292
rect 9585 2255 9643 2261
rect 10597 2261 10609 2264
rect 10643 2261 10655 2295
rect 10597 2255 10655 2261
rect 11333 2295 11391 2301
rect 11333 2261 11345 2295
rect 11379 2292 11391 2295
rect 11514 2292 11520 2304
rect 11379 2264 11520 2292
rect 11379 2261 11391 2264
rect 11333 2255 11391 2261
rect 11514 2252 11520 2264
rect 11572 2252 11578 2304
rect 12084 2292 12112 2400
rect 12544 2332 12848 2360
rect 12544 2292 12572 2332
rect 12084 2264 12572 2292
rect 12618 2252 12624 2304
rect 12676 2252 12682 2304
rect 12820 2301 12848 2332
rect 12894 2320 12900 2372
rect 12952 2360 12958 2372
rect 13188 2369 13216 2468
rect 13449 2465 13461 2468
rect 13495 2465 13507 2499
rect 13449 2459 13507 2465
rect 13464 2428 13492 2459
rect 13538 2456 13544 2508
rect 13596 2456 13602 2508
rect 13722 2456 13728 2508
rect 13780 2456 13786 2508
rect 13814 2456 13820 2508
rect 13872 2456 13878 2508
rect 13909 2499 13967 2505
rect 13909 2465 13921 2499
rect 13955 2465 13967 2499
rect 13909 2459 13967 2465
rect 13924 2428 13952 2459
rect 14550 2456 14556 2508
rect 14608 2496 14614 2508
rect 14645 2499 14703 2505
rect 14645 2496 14657 2499
rect 14608 2468 14657 2496
rect 14608 2456 14614 2468
rect 14645 2465 14657 2468
rect 14691 2465 14703 2499
rect 14921 2499 14979 2505
rect 14921 2496 14933 2499
rect 14645 2459 14703 2465
rect 14752 2468 14933 2496
rect 13464 2400 13952 2428
rect 13173 2363 13231 2369
rect 13173 2360 13185 2363
rect 12952 2332 13185 2360
rect 12952 2320 12958 2332
rect 13173 2329 13185 2332
rect 13219 2329 13231 2363
rect 14752 2360 14780 2468
rect 14921 2465 14933 2468
rect 14967 2465 14979 2499
rect 14921 2459 14979 2465
rect 15010 2456 15016 2508
rect 15068 2456 15074 2508
rect 15105 2499 15163 2505
rect 15105 2465 15117 2499
rect 15151 2496 15163 2499
rect 15194 2496 15200 2508
rect 15151 2468 15200 2496
rect 15151 2465 15163 2468
rect 15105 2459 15163 2465
rect 15194 2456 15200 2468
rect 15252 2456 15258 2508
rect 15378 2456 15384 2508
rect 15436 2456 15442 2508
rect 15565 2499 15623 2505
rect 15565 2465 15577 2499
rect 15611 2465 15623 2499
rect 15565 2459 15623 2465
rect 15580 2428 15608 2459
rect 16298 2456 16304 2508
rect 16356 2456 16362 2508
rect 16408 2505 16436 2536
rect 16500 2536 16856 2564
rect 16500 2505 16528 2536
rect 16850 2524 16856 2536
rect 16908 2524 16914 2576
rect 17313 2567 17371 2573
rect 17313 2533 17325 2567
rect 17359 2564 17371 2567
rect 17770 2564 17776 2576
rect 17359 2536 17776 2564
rect 17359 2533 17371 2536
rect 17313 2527 17371 2533
rect 17770 2524 17776 2536
rect 17828 2564 17834 2576
rect 18509 2567 18567 2573
rect 18509 2564 18521 2567
rect 17828 2536 18521 2564
rect 17828 2524 17834 2536
rect 18509 2533 18521 2536
rect 18555 2564 18567 2567
rect 18877 2567 18935 2573
rect 18877 2564 18889 2567
rect 18555 2536 18889 2564
rect 18555 2533 18567 2536
rect 18509 2527 18567 2533
rect 18877 2533 18889 2536
rect 18923 2533 18935 2567
rect 21450 2564 21456 2576
rect 18877 2527 18935 2533
rect 18984 2536 20944 2564
rect 16393 2499 16451 2505
rect 16393 2465 16405 2499
rect 16439 2465 16451 2499
rect 16393 2459 16451 2465
rect 16485 2499 16543 2505
rect 16485 2465 16497 2499
rect 16531 2465 16543 2499
rect 16485 2459 16543 2465
rect 16761 2499 16819 2505
rect 16761 2465 16773 2499
rect 16807 2465 16819 2499
rect 16761 2459 16819 2465
rect 14936 2400 15608 2428
rect 14936 2369 14964 2400
rect 16206 2388 16212 2440
rect 16264 2428 16270 2440
rect 16776 2428 16804 2459
rect 17034 2456 17040 2508
rect 17092 2456 17098 2508
rect 17129 2499 17187 2505
rect 17129 2465 17141 2499
rect 17175 2465 17187 2499
rect 17129 2459 17187 2465
rect 16264 2400 16804 2428
rect 16264 2388 16270 2400
rect 16850 2388 16856 2440
rect 16908 2428 16914 2440
rect 17144 2428 17172 2459
rect 17678 2456 17684 2508
rect 17736 2496 17742 2508
rect 18693 2499 18751 2505
rect 18693 2496 18705 2499
rect 17736 2468 18705 2496
rect 17736 2456 17742 2468
rect 18693 2465 18705 2468
rect 18739 2465 18751 2499
rect 18693 2459 18751 2465
rect 16908 2400 17172 2428
rect 18708 2428 18736 2459
rect 18782 2456 18788 2508
rect 18840 2456 18846 2508
rect 18984 2428 19012 2536
rect 19150 2456 19156 2508
rect 19208 2456 19214 2508
rect 20257 2499 20315 2505
rect 19260 2468 20208 2496
rect 18708 2400 19012 2428
rect 16908 2388 16914 2400
rect 13173 2323 13231 2329
rect 13280 2332 14780 2360
rect 14921 2363 14979 2369
rect 12805 2295 12863 2301
rect 12805 2261 12817 2295
rect 12851 2292 12863 2295
rect 13280 2292 13308 2332
rect 14921 2329 14933 2363
rect 14967 2329 14979 2363
rect 14921 2323 14979 2329
rect 15289 2363 15347 2369
rect 15289 2329 15301 2363
rect 15335 2360 15347 2363
rect 15378 2360 15384 2372
rect 15335 2332 15384 2360
rect 15335 2329 15347 2332
rect 15289 2323 15347 2329
rect 15378 2320 15384 2332
rect 15436 2320 15442 2372
rect 15565 2363 15623 2369
rect 15565 2329 15577 2363
rect 15611 2360 15623 2363
rect 17862 2360 17868 2372
rect 15611 2332 17868 2360
rect 15611 2329 15623 2332
rect 15565 2323 15623 2329
rect 17862 2320 17868 2332
rect 17920 2320 17926 2372
rect 19260 2360 19288 2468
rect 17972 2332 19288 2360
rect 12851 2264 13308 2292
rect 13541 2295 13599 2301
rect 12851 2261 12863 2264
rect 12805 2255 12863 2261
rect 13541 2261 13553 2295
rect 13587 2292 13599 2295
rect 13998 2292 14004 2304
rect 13587 2264 14004 2292
rect 13587 2261 13599 2264
rect 13541 2255 13599 2261
rect 13998 2252 14004 2264
rect 14056 2252 14062 2304
rect 14090 2252 14096 2304
rect 14148 2252 14154 2304
rect 16117 2295 16175 2301
rect 16117 2261 16129 2295
rect 16163 2292 16175 2295
rect 16206 2292 16212 2304
rect 16163 2264 16212 2292
rect 16163 2261 16175 2264
rect 16117 2255 16175 2261
rect 16206 2252 16212 2264
rect 16264 2252 16270 2304
rect 16761 2295 16819 2301
rect 16761 2261 16773 2295
rect 16807 2292 16819 2295
rect 17034 2292 17040 2304
rect 16807 2264 17040 2292
rect 16807 2261 16819 2264
rect 16761 2255 16819 2261
rect 17034 2252 17040 2264
rect 17092 2252 17098 2304
rect 17126 2252 17132 2304
rect 17184 2292 17190 2304
rect 17313 2295 17371 2301
rect 17313 2292 17325 2295
rect 17184 2264 17325 2292
rect 17184 2252 17190 2264
rect 17313 2261 17325 2264
rect 17359 2261 17371 2295
rect 17313 2255 17371 2261
rect 17402 2252 17408 2304
rect 17460 2292 17466 2304
rect 17972 2292 18000 2332
rect 19794 2320 19800 2372
rect 19852 2360 19858 2372
rect 20073 2363 20131 2369
rect 20073 2360 20085 2363
rect 19852 2332 20085 2360
rect 19852 2320 19858 2332
rect 20073 2329 20085 2332
rect 20119 2329 20131 2363
rect 20180 2360 20208 2468
rect 20257 2465 20269 2499
rect 20303 2465 20315 2499
rect 20257 2459 20315 2465
rect 20625 2499 20683 2505
rect 20625 2465 20637 2499
rect 20671 2496 20683 2499
rect 20714 2496 20720 2508
rect 20671 2468 20720 2496
rect 20671 2465 20683 2468
rect 20625 2459 20683 2465
rect 20272 2428 20300 2459
rect 20714 2456 20720 2468
rect 20772 2456 20778 2508
rect 20806 2428 20812 2440
rect 20272 2400 20812 2428
rect 20806 2388 20812 2400
rect 20864 2388 20870 2440
rect 20916 2428 20944 2536
rect 21284 2536 21456 2564
rect 21284 2505 21312 2536
rect 21450 2524 21456 2536
rect 21508 2524 21514 2576
rect 21545 2567 21603 2573
rect 21545 2533 21557 2567
rect 21591 2564 21603 2567
rect 21913 2567 21971 2573
rect 21913 2564 21925 2567
rect 21591 2536 21925 2564
rect 21591 2533 21603 2536
rect 21545 2527 21603 2533
rect 21269 2499 21327 2505
rect 21269 2465 21281 2499
rect 21315 2465 21327 2499
rect 21269 2459 21327 2465
rect 21361 2499 21419 2505
rect 21361 2465 21373 2499
rect 21407 2465 21419 2499
rect 21361 2459 21419 2465
rect 21376 2428 21404 2459
rect 21634 2456 21640 2508
rect 21692 2456 21698 2508
rect 21729 2499 21787 2505
rect 21729 2465 21741 2499
rect 21775 2465 21787 2499
rect 21729 2459 21787 2465
rect 20916 2400 21404 2428
rect 20254 2360 20260 2372
rect 20180 2332 20260 2360
rect 20073 2323 20131 2329
rect 20254 2320 20260 2332
rect 20312 2320 20318 2372
rect 21744 2360 21772 2459
rect 20364 2332 21772 2360
rect 21836 2360 21864 2536
rect 21913 2533 21925 2536
rect 21959 2533 21971 2567
rect 22296 2564 22324 2604
rect 22370 2592 22376 2644
rect 22428 2632 22434 2644
rect 23106 2632 23112 2644
rect 22428 2604 23112 2632
rect 22428 2592 22434 2604
rect 23106 2592 23112 2604
rect 23164 2592 23170 2644
rect 22741 2567 22799 2573
rect 22741 2564 22753 2567
rect 22296 2536 22753 2564
rect 21913 2527 21971 2533
rect 22741 2533 22753 2536
rect 22787 2533 22799 2567
rect 22741 2527 22799 2533
rect 22186 2456 22192 2508
rect 22244 2456 22250 2508
rect 22281 2499 22339 2505
rect 22281 2465 22293 2499
rect 22327 2465 22339 2499
rect 22281 2459 22339 2465
rect 21910 2388 21916 2440
rect 21968 2428 21974 2440
rect 22296 2428 22324 2459
rect 22462 2456 22468 2508
rect 22520 2456 22526 2508
rect 22557 2499 22615 2505
rect 22557 2465 22569 2499
rect 22603 2465 22615 2499
rect 22557 2459 22615 2465
rect 22833 2499 22891 2505
rect 22833 2465 22845 2499
rect 22879 2496 22891 2499
rect 22922 2496 22928 2508
rect 22879 2468 22928 2496
rect 22879 2465 22891 2468
rect 22833 2459 22891 2465
rect 22572 2428 22600 2459
rect 22922 2456 22928 2468
rect 22980 2456 22986 2508
rect 21968 2400 22324 2428
rect 22480 2400 22600 2428
rect 21968 2388 21974 2400
rect 22480 2369 22508 2400
rect 22465 2363 22523 2369
rect 22465 2360 22477 2363
rect 21836 2332 22477 2360
rect 17460 2264 18000 2292
rect 18509 2295 18567 2301
rect 17460 2252 17466 2264
rect 18509 2261 18521 2295
rect 18555 2292 18567 2295
rect 18598 2292 18604 2304
rect 18555 2264 18604 2292
rect 18555 2261 18567 2264
rect 18509 2255 18567 2261
rect 18598 2252 18604 2264
rect 18656 2252 18662 2304
rect 18874 2252 18880 2304
rect 18932 2252 18938 2304
rect 18966 2252 18972 2304
rect 19024 2292 19030 2304
rect 20364 2292 20392 2332
rect 22465 2329 22477 2332
rect 22511 2329 22523 2363
rect 22465 2323 22523 2329
rect 19024 2264 20392 2292
rect 19024 2252 19030 2264
rect 20438 2252 20444 2304
rect 20496 2252 20502 2304
rect 20806 2252 20812 2304
rect 20864 2292 20870 2304
rect 20901 2295 20959 2301
rect 20901 2292 20913 2295
rect 20864 2264 20913 2292
rect 20864 2252 20870 2264
rect 20901 2261 20913 2264
rect 20947 2261 20959 2295
rect 20901 2255 20959 2261
rect 21358 2252 21364 2304
rect 21416 2292 21422 2304
rect 21545 2295 21603 2301
rect 21545 2292 21557 2295
rect 21416 2264 21557 2292
rect 21416 2252 21422 2264
rect 21545 2261 21557 2264
rect 21591 2261 21603 2295
rect 21545 2255 21603 2261
rect 21910 2252 21916 2304
rect 21968 2252 21974 2304
rect 22094 2252 22100 2304
rect 22152 2292 22158 2304
rect 22370 2292 22376 2304
rect 22152 2264 22376 2292
rect 22152 2252 22158 2264
rect 22370 2252 22376 2264
rect 22428 2252 22434 2304
rect 22554 2252 22560 2304
rect 22612 2252 22618 2304
rect 552 2202 23368 2224
rect 552 2150 1366 2202
rect 1418 2150 1430 2202
rect 1482 2150 1494 2202
rect 1546 2150 1558 2202
rect 1610 2150 1622 2202
rect 1674 2150 1686 2202
rect 1738 2150 7366 2202
rect 7418 2150 7430 2202
rect 7482 2150 7494 2202
rect 7546 2150 7558 2202
rect 7610 2150 7622 2202
rect 7674 2150 7686 2202
rect 7738 2150 13366 2202
rect 13418 2150 13430 2202
rect 13482 2150 13494 2202
rect 13546 2150 13558 2202
rect 13610 2150 13622 2202
rect 13674 2150 13686 2202
rect 13738 2150 19366 2202
rect 19418 2150 19430 2202
rect 19482 2150 19494 2202
rect 19546 2150 19558 2202
rect 19610 2150 19622 2202
rect 19674 2150 19686 2202
rect 19738 2150 23368 2202
rect 552 2128 23368 2150
rect 3326 2048 3332 2100
rect 3384 2088 3390 2100
rect 3421 2091 3479 2097
rect 3421 2088 3433 2091
rect 3384 2060 3433 2088
rect 3384 2048 3390 2060
rect 3421 2057 3433 2060
rect 3467 2057 3479 2091
rect 3421 2051 3479 2057
rect 3804 2060 4016 2088
rect 1854 1980 1860 2032
rect 1912 2020 1918 2032
rect 3804 2020 3832 2060
rect 1912 1992 3832 2020
rect 1912 1980 1918 1992
rect 3878 1980 3884 2032
rect 3936 1980 3942 2032
rect 3988 2020 4016 2060
rect 5810 2048 5816 2100
rect 5868 2088 5874 2100
rect 6273 2091 6331 2097
rect 6273 2088 6285 2091
rect 5868 2060 6285 2088
rect 5868 2048 5874 2060
rect 6273 2057 6285 2060
rect 6319 2057 6331 2091
rect 6273 2051 6331 2057
rect 7282 2048 7288 2100
rect 7340 2088 7346 2100
rect 7377 2091 7435 2097
rect 7377 2088 7389 2091
rect 7340 2060 7389 2088
rect 7340 2048 7346 2060
rect 7377 2057 7389 2060
rect 7423 2057 7435 2091
rect 7377 2051 7435 2057
rect 8754 2048 8760 2100
rect 8812 2048 8818 2100
rect 8938 2048 8944 2100
rect 8996 2088 9002 2100
rect 8996 2060 10272 2088
rect 8996 2048 9002 2060
rect 6638 2020 6644 2032
rect 3988 1992 6644 2020
rect 6638 1980 6644 1992
rect 6696 1980 6702 2032
rect 10042 2020 10048 2032
rect 8220 1992 10048 2020
rect 2409 1955 2467 1961
rect 2409 1921 2421 1955
rect 2455 1952 2467 1955
rect 2498 1952 2504 1964
rect 2455 1924 2504 1952
rect 2455 1921 2467 1924
rect 2409 1915 2467 1921
rect 2498 1912 2504 1924
rect 2556 1912 2562 1964
rect 3896 1952 3924 1980
rect 5537 1955 5595 1961
rect 5537 1952 5549 1955
rect 3896 1924 5549 1952
rect 1029 1887 1087 1893
rect 1029 1853 1041 1887
rect 1075 1853 1087 1887
rect 1029 1847 1087 1853
rect 1044 1816 1072 1847
rect 1946 1844 1952 1896
rect 2004 1884 2010 1896
rect 2317 1887 2375 1893
rect 2317 1884 2329 1887
rect 2004 1856 2329 1884
rect 2004 1844 2010 1856
rect 2317 1853 2329 1856
rect 2363 1853 2375 1887
rect 2317 1847 2375 1853
rect 3050 1844 3056 1896
rect 3108 1844 3114 1896
rect 3418 1844 3424 1896
rect 3476 1884 3482 1896
rect 3789 1887 3847 1893
rect 3789 1884 3801 1887
rect 3476 1856 3801 1884
rect 3476 1844 3482 1856
rect 3789 1853 3801 1856
rect 3835 1853 3847 1887
rect 3789 1847 3847 1853
rect 1044 1788 3280 1816
rect 845 1751 903 1757
rect 845 1748 857 1751
rect 492 1720 857 1748
rect 492 1408 520 1720
rect 845 1717 857 1720
rect 891 1717 903 1751
rect 845 1711 903 1717
rect 2682 1708 2688 1760
rect 2740 1708 2746 1760
rect 2774 1708 2780 1760
rect 2832 1748 2838 1760
rect 2961 1751 3019 1757
rect 2961 1748 2973 1751
rect 2832 1720 2973 1748
rect 2832 1708 2838 1720
rect 2961 1717 2973 1720
rect 3007 1717 3019 1751
rect 3252 1748 3280 1788
rect 3326 1776 3332 1828
rect 3384 1816 3390 1828
rect 3605 1819 3663 1825
rect 3605 1816 3617 1819
rect 3384 1788 3617 1816
rect 3384 1776 3390 1788
rect 3605 1785 3617 1788
rect 3651 1816 3663 1819
rect 3896 1816 3924 1924
rect 5537 1921 5549 1924
rect 5583 1921 5595 1955
rect 5537 1915 5595 1921
rect 6089 1955 6147 1961
rect 6089 1921 6101 1955
rect 6135 1952 6147 1955
rect 6178 1952 6184 1964
rect 6135 1924 6184 1952
rect 6135 1921 6147 1924
rect 6089 1915 6147 1921
rect 6178 1912 6184 1924
rect 6236 1912 6242 1964
rect 6730 1912 6736 1964
rect 6788 1952 6794 1964
rect 6788 1924 7512 1952
rect 6788 1912 6794 1924
rect 4065 1887 4123 1893
rect 4065 1853 4077 1887
rect 4111 1853 4123 1887
rect 4065 1847 4123 1853
rect 4525 1887 4583 1893
rect 4525 1853 4537 1887
rect 4571 1884 4583 1887
rect 4982 1884 4988 1896
rect 4571 1856 4988 1884
rect 4571 1853 4583 1856
rect 4525 1847 4583 1853
rect 3651 1788 3924 1816
rect 4080 1816 4108 1847
rect 4982 1844 4988 1856
rect 5040 1844 5046 1896
rect 5258 1844 5264 1896
rect 5316 1844 5322 1896
rect 5718 1844 5724 1896
rect 5776 1844 5782 1896
rect 5994 1844 6000 1896
rect 6052 1884 6058 1896
rect 6549 1887 6607 1893
rect 6549 1884 6561 1887
rect 6052 1856 6561 1884
rect 6052 1844 6058 1856
rect 6549 1853 6561 1856
rect 6595 1884 6607 1887
rect 7006 1884 7012 1896
rect 6595 1856 7012 1884
rect 6595 1853 6607 1856
rect 6549 1847 6607 1853
rect 7006 1844 7012 1856
rect 7064 1844 7070 1896
rect 7098 1844 7104 1896
rect 7156 1884 7162 1896
rect 7484 1893 7512 1924
rect 8220 1893 8248 1992
rect 10042 1980 10048 1992
rect 10100 1980 10106 2032
rect 10137 2023 10195 2029
rect 10137 1989 10149 2023
rect 10183 1989 10195 2023
rect 10244 2020 10272 2060
rect 10410 2048 10416 2100
rect 10468 2088 10474 2100
rect 11606 2088 11612 2100
rect 10468 2060 11612 2088
rect 10468 2048 10474 2060
rect 11606 2048 11612 2060
rect 11664 2048 11670 2100
rect 11882 2048 11888 2100
rect 11940 2048 11946 2100
rect 13262 2088 13268 2100
rect 12406 2060 13268 2088
rect 12406 2020 12434 2060
rect 13262 2048 13268 2060
rect 13320 2048 13326 2100
rect 14090 2048 14096 2100
rect 14148 2088 14154 2100
rect 16574 2088 16580 2100
rect 14148 2060 16580 2088
rect 14148 2048 14154 2060
rect 16574 2048 16580 2060
rect 16632 2048 16638 2100
rect 17034 2048 17040 2100
rect 17092 2088 17098 2100
rect 19705 2091 19763 2097
rect 19705 2088 19717 2091
rect 17092 2060 19717 2088
rect 17092 2048 17098 2060
rect 19705 2057 19717 2060
rect 19751 2057 19763 2091
rect 19705 2051 19763 2057
rect 20070 2048 20076 2100
rect 20128 2048 20134 2100
rect 20901 2091 20959 2097
rect 20901 2057 20913 2091
rect 20947 2088 20959 2091
rect 22186 2088 22192 2100
rect 20947 2060 22192 2088
rect 20947 2057 20959 2060
rect 20901 2051 20959 2057
rect 22186 2048 22192 2060
rect 22244 2048 22250 2100
rect 22370 2048 22376 2100
rect 22428 2048 22434 2100
rect 22465 2091 22523 2097
rect 22465 2057 22477 2091
rect 22511 2088 22523 2091
rect 22554 2088 22560 2100
rect 22511 2060 22560 2088
rect 22511 2057 22523 2060
rect 22465 2051 22523 2057
rect 22554 2048 22560 2060
rect 22612 2048 22618 2100
rect 10244 1992 12434 2020
rect 10137 1983 10195 1989
rect 8573 1955 8631 1961
rect 8573 1952 8585 1955
rect 8404 1924 8585 1952
rect 7285 1887 7343 1893
rect 7285 1884 7297 1887
rect 7156 1856 7297 1884
rect 7156 1844 7162 1856
rect 7285 1853 7297 1856
rect 7331 1853 7343 1887
rect 7285 1847 7343 1853
rect 7469 1887 7527 1893
rect 7469 1853 7481 1887
rect 7515 1853 7527 1887
rect 7469 1847 7527 1853
rect 8205 1887 8263 1893
rect 8205 1853 8217 1887
rect 8251 1853 8263 1887
rect 8205 1847 8263 1853
rect 5442 1816 5448 1828
rect 4080 1788 5448 1816
rect 3651 1785 3663 1788
rect 3605 1779 3663 1785
rect 5442 1776 5448 1788
rect 5500 1776 5506 1828
rect 3970 1748 3976 1760
rect 3252 1720 3976 1748
rect 2961 1711 3019 1717
rect 3970 1708 3976 1720
rect 4028 1708 4034 1760
rect 4154 1708 4160 1760
rect 4212 1748 4218 1760
rect 4433 1751 4491 1757
rect 4433 1748 4445 1751
rect 4212 1720 4445 1748
rect 4212 1708 4218 1720
rect 4433 1717 4445 1720
rect 4479 1717 4491 1751
rect 4433 1711 4491 1717
rect 4890 1708 4896 1760
rect 4948 1748 4954 1760
rect 5169 1751 5227 1757
rect 5169 1748 5181 1751
rect 4948 1720 5181 1748
rect 4948 1708 4954 1720
rect 5169 1717 5181 1720
rect 5215 1717 5227 1751
rect 5169 1711 5227 1717
rect 5902 1708 5908 1760
rect 5960 1708 5966 1760
rect 7926 1708 7932 1760
rect 7984 1748 7990 1760
rect 8021 1751 8079 1757
rect 8021 1748 8033 1751
rect 7984 1720 8033 1748
rect 7984 1708 7990 1720
rect 8021 1717 8033 1720
rect 8067 1748 8079 1751
rect 8404 1748 8432 1924
rect 8573 1921 8585 1924
rect 8619 1921 8631 1955
rect 8941 1955 8999 1961
rect 8941 1952 8953 1955
rect 8573 1915 8631 1921
rect 8772 1924 8953 1952
rect 8478 1844 8484 1896
rect 8536 1884 8542 1896
rect 8772 1884 8800 1924
rect 8941 1921 8953 1924
rect 8987 1921 8999 1955
rect 10152 1952 10180 1983
rect 13998 1980 14004 2032
rect 14056 2020 14062 2032
rect 17865 2023 17923 2029
rect 17865 2020 17877 2023
rect 14056 1992 17877 2020
rect 14056 1980 14062 1992
rect 17865 1989 17877 1992
rect 17911 1989 17923 2023
rect 19978 2020 19984 2032
rect 17865 1983 17923 1989
rect 17972 1992 19984 2020
rect 10152 1924 11284 1952
rect 8941 1915 8999 1921
rect 11256 1896 11284 1924
rect 12434 1912 12440 1964
rect 12492 1952 12498 1964
rect 14274 1952 14280 1964
rect 12492 1924 14280 1952
rect 12492 1912 12498 1924
rect 14274 1912 14280 1924
rect 14332 1912 14338 1964
rect 14366 1912 14372 1964
rect 14424 1952 14430 1964
rect 15841 1955 15899 1961
rect 14424 1924 15792 1952
rect 14424 1912 14430 1924
rect 8536 1856 8800 1884
rect 8849 1887 8907 1893
rect 8536 1844 8542 1856
rect 8849 1853 8861 1887
rect 8895 1884 8907 1887
rect 8895 1856 9076 1884
rect 8895 1853 8907 1856
rect 8849 1847 8907 1853
rect 9048 1828 9076 1856
rect 9122 1844 9128 1896
rect 9180 1844 9186 1896
rect 9217 1887 9275 1893
rect 9217 1853 9229 1887
rect 9263 1853 9275 1887
rect 9217 1847 9275 1853
rect 8662 1776 8668 1828
rect 8720 1816 8726 1828
rect 8941 1819 8999 1825
rect 8941 1816 8953 1819
rect 8720 1788 8953 1816
rect 8720 1776 8726 1788
rect 8941 1785 8953 1788
rect 8987 1785 8999 1819
rect 8941 1779 8999 1785
rect 9030 1776 9036 1828
rect 9088 1816 9094 1828
rect 9232 1816 9260 1847
rect 9306 1844 9312 1896
rect 9364 1844 9370 1896
rect 9858 1844 9864 1896
rect 9916 1844 9922 1896
rect 9950 1844 9956 1896
rect 10008 1844 10014 1896
rect 10226 1844 10232 1896
rect 10284 1844 10290 1896
rect 10318 1844 10324 1896
rect 10376 1884 10382 1896
rect 10689 1887 10747 1893
rect 10689 1884 10701 1887
rect 10376 1856 10701 1884
rect 10376 1844 10382 1856
rect 10689 1853 10701 1856
rect 10735 1853 10747 1887
rect 10689 1847 10747 1853
rect 10870 1844 10876 1896
rect 10928 1893 10934 1896
rect 10928 1887 10950 1893
rect 10938 1853 10950 1887
rect 10928 1847 10950 1853
rect 10928 1844 10934 1847
rect 11238 1844 11244 1896
rect 11296 1844 11302 1896
rect 11333 1887 11391 1893
rect 11333 1853 11345 1887
rect 11379 1884 11391 1887
rect 11422 1884 11428 1896
rect 11379 1856 11428 1884
rect 11379 1853 11391 1856
rect 11333 1847 11391 1853
rect 9088 1788 9260 1816
rect 10975 1819 11033 1825
rect 9088 1776 9094 1788
rect 10975 1785 10987 1819
rect 11021 1816 11033 1819
rect 11348 1816 11376 1847
rect 11422 1844 11428 1856
rect 11480 1844 11486 1896
rect 11514 1844 11520 1896
rect 11572 1844 11578 1896
rect 11606 1844 11612 1896
rect 11664 1844 11670 1896
rect 11701 1887 11759 1893
rect 11701 1853 11713 1887
rect 11747 1884 11759 1887
rect 11882 1884 11888 1896
rect 11747 1856 11888 1884
rect 11747 1853 11759 1856
rect 11701 1847 11759 1853
rect 11882 1844 11888 1856
rect 11940 1844 11946 1896
rect 12069 1887 12127 1893
rect 12069 1853 12081 1887
rect 12115 1884 12127 1887
rect 12342 1884 12348 1896
rect 12115 1856 12348 1884
rect 12115 1853 12127 1856
rect 12069 1847 12127 1853
rect 12342 1844 12348 1856
rect 12400 1844 12406 1896
rect 12621 1887 12679 1893
rect 12621 1853 12633 1887
rect 12667 1884 12679 1887
rect 12710 1884 12716 1896
rect 12667 1856 12716 1884
rect 12667 1853 12679 1856
rect 12621 1847 12679 1853
rect 12710 1844 12716 1856
rect 12768 1844 12774 1896
rect 12894 1844 12900 1896
rect 12952 1844 12958 1896
rect 14001 1887 14059 1893
rect 14001 1853 14013 1887
rect 14047 1884 14059 1887
rect 14458 1884 14464 1896
rect 14047 1856 14464 1884
rect 14047 1853 14059 1856
rect 14001 1847 14059 1853
rect 14458 1844 14464 1856
rect 14516 1844 14522 1896
rect 15562 1844 15568 1896
rect 15620 1844 15626 1896
rect 15654 1844 15660 1896
rect 15712 1844 15718 1896
rect 15764 1884 15792 1924
rect 15841 1921 15853 1955
rect 15887 1952 15899 1955
rect 16114 1952 16120 1964
rect 15887 1924 16120 1952
rect 15887 1921 15899 1924
rect 15841 1915 15899 1921
rect 16114 1912 16120 1924
rect 16172 1952 16178 1964
rect 17972 1952 18000 1992
rect 16172 1924 18000 1952
rect 16172 1912 16178 1924
rect 18046 1912 18052 1964
rect 18104 1912 18110 1964
rect 19904 1961 19932 1992
rect 19978 1980 19984 1992
rect 20036 1980 20042 2032
rect 20349 2023 20407 2029
rect 20349 1989 20361 2023
rect 20395 1989 20407 2023
rect 22002 2020 22008 2032
rect 20349 1983 20407 1989
rect 21100 1992 22008 2020
rect 19889 1955 19947 1961
rect 18616 1924 19656 1952
rect 17402 1884 17408 1896
rect 15764 1856 17408 1884
rect 17402 1844 17408 1856
rect 17460 1844 17466 1896
rect 17770 1844 17776 1896
rect 17828 1884 17834 1896
rect 18616 1884 18644 1924
rect 17828 1856 18644 1884
rect 17828 1844 17834 1856
rect 18690 1844 18696 1896
rect 18748 1844 18754 1896
rect 19628 1893 19656 1924
rect 19889 1921 19901 1955
rect 19935 1921 19947 1955
rect 19889 1915 19947 1921
rect 20254 1912 20260 1964
rect 20312 1912 20318 1964
rect 19521 1887 19579 1893
rect 19521 1853 19533 1887
rect 19567 1853 19579 1887
rect 19521 1847 19579 1853
rect 19613 1887 19671 1893
rect 19613 1853 19625 1887
rect 19659 1884 19671 1887
rect 19981 1887 20039 1893
rect 19981 1884 19993 1887
rect 19659 1856 19993 1884
rect 19659 1853 19671 1856
rect 19613 1847 19671 1853
rect 19981 1853 19993 1856
rect 20027 1884 20039 1887
rect 20364 1884 20392 1983
rect 20027 1856 20392 1884
rect 20533 1887 20591 1893
rect 20027 1853 20039 1856
rect 19981 1847 20039 1853
rect 20533 1853 20545 1887
rect 20579 1884 20591 1887
rect 20806 1884 20812 1896
rect 20579 1856 20812 1884
rect 20579 1853 20591 1856
rect 20533 1847 20591 1853
rect 11021 1788 11376 1816
rect 11021 1785 11033 1788
rect 10975 1779 11033 1785
rect 11256 1760 11284 1788
rect 13262 1776 13268 1828
rect 13320 1816 13326 1828
rect 13722 1816 13728 1828
rect 13320 1788 13728 1816
rect 13320 1776 13326 1788
rect 13722 1776 13728 1788
rect 13780 1816 13786 1828
rect 15841 1819 15899 1825
rect 15841 1816 15853 1819
rect 13780 1788 15853 1816
rect 13780 1776 13786 1788
rect 15841 1785 15853 1788
rect 15887 1785 15899 1819
rect 15841 1779 15899 1785
rect 15930 1776 15936 1828
rect 15988 1816 15994 1828
rect 18049 1819 18107 1825
rect 15988 1788 16988 1816
rect 15988 1776 15994 1788
rect 8067 1720 8432 1748
rect 8573 1751 8631 1757
rect 8067 1717 8079 1720
rect 8021 1711 8079 1717
rect 8573 1717 8585 1751
rect 8619 1748 8631 1751
rect 8846 1748 8852 1760
rect 8619 1720 8852 1748
rect 8619 1717 8631 1720
rect 8573 1711 8631 1717
rect 8846 1708 8852 1720
rect 8904 1708 8910 1760
rect 9214 1708 9220 1760
rect 9272 1748 9278 1760
rect 9493 1751 9551 1757
rect 9493 1748 9505 1751
rect 9272 1720 9505 1748
rect 9272 1708 9278 1720
rect 9493 1717 9505 1720
rect 9539 1717 9551 1751
rect 9493 1711 9551 1717
rect 9582 1708 9588 1760
rect 9640 1748 9646 1760
rect 9677 1751 9735 1757
rect 9677 1748 9689 1751
rect 9640 1720 9689 1748
rect 9640 1708 9646 1720
rect 9677 1717 9689 1720
rect 9723 1717 9735 1751
rect 9677 1711 9735 1717
rect 10778 1708 10784 1760
rect 10836 1748 10842 1760
rect 11057 1751 11115 1757
rect 11057 1748 11069 1751
rect 10836 1720 11069 1748
rect 10836 1708 10842 1720
rect 11057 1717 11069 1720
rect 11103 1717 11115 1751
rect 11057 1711 11115 1717
rect 11238 1708 11244 1760
rect 11296 1708 11302 1760
rect 11422 1708 11428 1760
rect 11480 1708 11486 1760
rect 12529 1751 12587 1757
rect 12529 1717 12541 1751
rect 12575 1748 12587 1751
rect 12618 1748 12624 1760
rect 12575 1720 12624 1748
rect 12575 1717 12587 1720
rect 12529 1711 12587 1717
rect 12618 1708 12624 1720
rect 12676 1708 12682 1760
rect 13078 1708 13084 1760
rect 13136 1708 13142 1760
rect 13170 1708 13176 1760
rect 13228 1748 13234 1760
rect 13630 1748 13636 1760
rect 13228 1720 13636 1748
rect 13228 1708 13234 1720
rect 13630 1708 13636 1720
rect 13688 1708 13694 1760
rect 13909 1751 13967 1757
rect 13909 1717 13921 1751
rect 13955 1748 13967 1751
rect 14642 1748 14648 1760
rect 13955 1720 14648 1748
rect 13955 1717 13967 1720
rect 13909 1711 13967 1717
rect 14642 1708 14648 1720
rect 14700 1708 14706 1760
rect 15746 1708 15752 1760
rect 15804 1748 15810 1760
rect 16850 1748 16856 1760
rect 15804 1720 16856 1748
rect 15804 1708 15810 1720
rect 16850 1708 16856 1720
rect 16908 1708 16914 1760
rect 16960 1748 16988 1788
rect 18049 1785 18061 1819
rect 18095 1816 18107 1819
rect 18322 1816 18328 1828
rect 18095 1788 18328 1816
rect 18095 1785 18107 1788
rect 18049 1779 18107 1785
rect 18322 1776 18328 1788
rect 18380 1776 18386 1828
rect 18966 1816 18972 1828
rect 18800 1788 18972 1816
rect 18800 1748 18828 1788
rect 18966 1776 18972 1788
rect 19024 1776 19030 1828
rect 19536 1816 19564 1847
rect 20548 1816 20576 1847
rect 20806 1844 20812 1856
rect 20864 1844 20870 1896
rect 21100 1893 21128 1992
rect 22002 1980 22008 1992
rect 22060 1980 22066 2032
rect 22094 1980 22100 2032
rect 22152 2020 22158 2032
rect 22833 2023 22891 2029
rect 22833 2020 22845 2023
rect 22152 1992 22845 2020
rect 22152 1980 22158 1992
rect 22833 1989 22845 1992
rect 22879 1989 22891 2023
rect 22833 1983 22891 1989
rect 22281 1955 22339 1961
rect 22281 1952 22293 1955
rect 21744 1924 22293 1952
rect 21744 1896 21772 1924
rect 22281 1921 22293 1924
rect 22327 1921 22339 1955
rect 22281 1915 22339 1921
rect 22370 1912 22376 1964
rect 22428 1952 22434 1964
rect 22428 1924 22692 1952
rect 22428 1912 22434 1924
rect 21085 1887 21143 1893
rect 21085 1853 21097 1887
rect 21131 1853 21143 1887
rect 21085 1847 21143 1853
rect 21358 1844 21364 1896
rect 21416 1844 21422 1896
rect 21542 1844 21548 1896
rect 21600 1844 21606 1896
rect 21726 1844 21732 1896
rect 21784 1844 21790 1896
rect 22189 1887 22247 1893
rect 22189 1853 22201 1887
rect 22235 1884 22247 1887
rect 22235 1856 22508 1884
rect 22235 1853 22247 1856
rect 22189 1847 22247 1853
rect 19536 1788 20576 1816
rect 21634 1776 21640 1828
rect 21692 1776 21698 1828
rect 16960 1720 18828 1748
rect 18877 1751 18935 1757
rect 18877 1717 18889 1751
rect 18923 1748 18935 1751
rect 19242 1748 19248 1760
rect 18923 1720 19248 1748
rect 18923 1717 18935 1720
rect 18877 1711 18935 1717
rect 19242 1708 19248 1720
rect 19300 1708 19306 1760
rect 19334 1708 19340 1760
rect 19392 1708 19398 1760
rect 19886 1708 19892 1760
rect 19944 1708 19950 1760
rect 19978 1708 19984 1760
rect 20036 1748 20042 1760
rect 20257 1751 20315 1757
rect 20257 1748 20269 1751
rect 20036 1720 20269 1748
rect 20036 1708 20042 1720
rect 20257 1717 20269 1720
rect 20303 1748 20315 1751
rect 21818 1748 21824 1760
rect 20303 1720 21824 1748
rect 20303 1717 20315 1720
rect 20257 1711 20315 1717
rect 21818 1708 21824 1720
rect 21876 1708 21882 1760
rect 22005 1751 22063 1757
rect 22005 1717 22017 1751
rect 22051 1748 22063 1751
rect 22186 1748 22192 1760
rect 22051 1720 22192 1748
rect 22051 1717 22063 1720
rect 22005 1711 22063 1717
rect 22186 1708 22192 1720
rect 22244 1708 22250 1760
rect 22480 1748 22508 1856
rect 22554 1844 22560 1896
rect 22612 1844 22618 1896
rect 22664 1893 22692 1924
rect 22649 1887 22707 1893
rect 22649 1853 22661 1887
rect 22695 1853 22707 1887
rect 22649 1847 22707 1853
rect 22738 1844 22744 1896
rect 22796 1884 22802 1896
rect 23198 1884 23204 1896
rect 22796 1856 23204 1884
rect 22796 1844 22802 1856
rect 23198 1844 23204 1856
rect 23256 1844 23262 1896
rect 22572 1816 22600 1844
rect 22922 1816 22928 1828
rect 22572 1788 22928 1816
rect 22922 1776 22928 1788
rect 22980 1776 22986 1828
rect 23014 1748 23020 1760
rect 22480 1720 23020 1748
rect 23014 1708 23020 1720
rect 23072 1708 23078 1760
rect 552 1658 23368 1680
rect 552 1606 4366 1658
rect 4418 1606 4430 1658
rect 4482 1606 4494 1658
rect 4546 1606 4558 1658
rect 4610 1606 4622 1658
rect 4674 1606 4686 1658
rect 4738 1606 10366 1658
rect 10418 1606 10430 1658
rect 10482 1606 10494 1658
rect 10546 1606 10558 1658
rect 10610 1606 10622 1658
rect 10674 1606 10686 1658
rect 10738 1606 16366 1658
rect 16418 1606 16430 1658
rect 16482 1606 16494 1658
rect 16546 1606 16558 1658
rect 16610 1606 16622 1658
rect 16674 1606 16686 1658
rect 16738 1606 22366 1658
rect 22418 1606 22430 1658
rect 22482 1606 22494 1658
rect 22546 1606 22558 1658
rect 22610 1606 22622 1658
rect 22674 1606 22686 1658
rect 22738 1606 23368 1658
rect 552 1584 23368 1606
rect 750 1504 756 1556
rect 808 1544 814 1556
rect 1029 1547 1087 1553
rect 1029 1544 1041 1547
rect 808 1516 1041 1544
rect 808 1504 814 1516
rect 1029 1513 1041 1516
rect 1075 1513 1087 1547
rect 1029 1507 1087 1513
rect 1305 1547 1363 1553
rect 1305 1513 1317 1547
rect 1351 1513 1363 1547
rect 1305 1507 1363 1513
rect 566 1436 572 1488
rect 624 1476 630 1488
rect 1320 1476 1348 1507
rect 2222 1504 2228 1556
rect 2280 1544 2286 1556
rect 2501 1547 2559 1553
rect 2501 1544 2513 1547
rect 2280 1516 2513 1544
rect 2280 1504 2286 1516
rect 2501 1513 2513 1516
rect 2547 1513 2559 1547
rect 2501 1507 2559 1513
rect 2608 1516 5856 1544
rect 2608 1476 2636 1516
rect 624 1448 1348 1476
rect 1504 1448 2636 1476
rect 624 1436 630 1448
rect 1504 1417 1532 1448
rect 2682 1436 2688 1488
rect 2740 1476 2746 1488
rect 2740 1448 4660 1476
rect 2740 1436 2746 1448
rect 845 1411 903 1417
rect 845 1408 857 1411
rect 492 1380 857 1408
rect 845 1377 857 1380
rect 891 1377 903 1411
rect 845 1371 903 1377
rect 1489 1411 1547 1417
rect 1489 1377 1501 1411
rect 1535 1377 1547 1411
rect 1489 1371 1547 1377
rect 1854 1368 1860 1420
rect 1912 1368 1918 1420
rect 1946 1368 1952 1420
rect 2004 1408 2010 1420
rect 2041 1411 2099 1417
rect 2041 1408 2053 1411
rect 2004 1380 2053 1408
rect 2004 1368 2010 1380
rect 2041 1377 2053 1380
rect 2087 1377 2099 1411
rect 2041 1371 2099 1377
rect 2133 1411 2191 1417
rect 2133 1377 2145 1411
rect 2179 1408 2191 1411
rect 2317 1411 2375 1417
rect 2317 1408 2329 1411
rect 2179 1380 2329 1408
rect 2179 1377 2191 1380
rect 2133 1371 2191 1377
rect 2317 1377 2329 1380
rect 2363 1377 2375 1411
rect 2317 1371 2375 1377
rect 2774 1368 2780 1420
rect 2832 1368 2838 1420
rect 3326 1368 3332 1420
rect 3384 1368 3390 1420
rect 3973 1411 4031 1417
rect 3973 1377 3985 1411
rect 4019 1408 4031 1411
rect 4246 1408 4252 1420
rect 4019 1380 4252 1408
rect 4019 1377 4031 1380
rect 3973 1371 4031 1377
rect 4246 1368 4252 1380
rect 4304 1368 4310 1420
rect 4632 1417 4660 1448
rect 5442 1436 5448 1488
rect 5500 1436 5506 1488
rect 5828 1476 5856 1516
rect 6638 1504 6644 1556
rect 6696 1544 6702 1556
rect 7193 1547 7251 1553
rect 7193 1544 7205 1547
rect 6696 1516 7205 1544
rect 6696 1504 6702 1516
rect 7193 1513 7205 1516
rect 7239 1513 7251 1547
rect 7193 1507 7251 1513
rect 7300 1516 8064 1544
rect 7300 1476 7328 1516
rect 8036 1476 8064 1516
rect 8294 1504 8300 1556
rect 8352 1504 8358 1556
rect 9217 1547 9275 1553
rect 9217 1513 9229 1547
rect 9263 1544 9275 1547
rect 9306 1544 9312 1556
rect 9263 1516 9312 1544
rect 9263 1513 9275 1516
rect 9217 1507 9275 1513
rect 9306 1504 9312 1516
rect 9364 1504 9370 1556
rect 12526 1504 12532 1556
rect 12584 1504 12590 1556
rect 13078 1504 13084 1556
rect 13136 1544 13142 1556
rect 15282 1547 15340 1553
rect 15282 1544 15294 1547
rect 13136 1516 14228 1544
rect 13136 1504 13142 1516
rect 8570 1476 8576 1488
rect 5828 1448 7328 1476
rect 7392 1448 7972 1476
rect 8036 1448 8576 1476
rect 4617 1411 4675 1417
rect 4617 1377 4629 1411
rect 4663 1377 4675 1411
rect 4617 1371 4675 1377
rect 5261 1411 5319 1417
rect 5261 1377 5273 1411
rect 5307 1408 5319 1411
rect 5718 1408 5724 1420
rect 5307 1380 5724 1408
rect 5307 1377 5319 1380
rect 5261 1371 5319 1377
rect 5718 1368 5724 1380
rect 5776 1368 5782 1420
rect 5994 1368 6000 1420
rect 6052 1368 6058 1420
rect 6730 1368 6736 1420
rect 6788 1368 6794 1420
rect 7392 1417 7420 1448
rect 7944 1420 7972 1448
rect 8570 1436 8576 1448
rect 8628 1436 8634 1488
rect 9122 1476 9128 1488
rect 8680 1448 9128 1476
rect 7377 1411 7435 1417
rect 7377 1377 7389 1411
rect 7423 1377 7435 1411
rect 7377 1371 7435 1377
rect 7561 1411 7619 1417
rect 7561 1377 7573 1411
rect 7607 1408 7619 1411
rect 7834 1408 7840 1420
rect 7607 1380 7840 1408
rect 7607 1377 7619 1380
rect 7561 1371 7619 1377
rect 7834 1368 7840 1380
rect 7892 1368 7898 1420
rect 7926 1368 7932 1420
rect 7984 1368 7990 1420
rect 8110 1368 8116 1420
rect 8168 1368 8174 1420
rect 8478 1368 8484 1420
rect 8536 1368 8542 1420
rect 8680 1417 8708 1448
rect 9122 1436 9128 1448
rect 9180 1436 9186 1488
rect 12263 1479 12321 1485
rect 9600 1448 10456 1476
rect 8665 1411 8723 1417
rect 8665 1377 8677 1411
rect 8711 1377 8723 1411
rect 8665 1371 8723 1377
rect 8938 1368 8944 1420
rect 8996 1368 9002 1420
rect 9033 1411 9091 1417
rect 9033 1377 9045 1411
rect 9079 1408 9091 1411
rect 9398 1408 9404 1420
rect 9079 1380 9404 1408
rect 9079 1377 9091 1380
rect 9033 1371 9091 1377
rect 9398 1368 9404 1380
rect 9456 1368 9462 1420
rect 9600 1417 9628 1448
rect 9585 1411 9643 1417
rect 9585 1377 9597 1411
rect 9631 1377 9643 1411
rect 9585 1371 9643 1377
rect 3421 1343 3479 1349
rect 3421 1309 3433 1343
rect 3467 1340 3479 1343
rect 3602 1340 3608 1352
rect 3467 1312 3608 1340
rect 3467 1309 3479 1312
rect 3421 1303 3479 1309
rect 3602 1300 3608 1312
rect 3660 1300 3666 1352
rect 3697 1343 3755 1349
rect 3697 1309 3709 1343
rect 3743 1340 3755 1343
rect 3881 1343 3939 1349
rect 3881 1340 3893 1343
rect 3743 1312 3893 1340
rect 3743 1309 3755 1312
rect 3697 1303 3755 1309
rect 3881 1309 3893 1312
rect 3927 1309 3939 1343
rect 4525 1343 4583 1349
rect 4525 1340 4537 1343
rect 3881 1303 3939 1309
rect 4356 1312 4537 1340
rect 4356 1281 4384 1312
rect 4525 1309 4537 1312
rect 4571 1309 4583 1343
rect 5905 1343 5963 1349
rect 5905 1340 5917 1343
rect 4525 1303 4583 1309
rect 5000 1312 5917 1340
rect 5000 1281 5028 1312
rect 5905 1309 5917 1312
rect 5951 1309 5963 1343
rect 5905 1303 5963 1309
rect 6822 1300 6828 1352
rect 6880 1300 6886 1352
rect 7098 1300 7104 1352
rect 7156 1300 7162 1352
rect 7653 1343 7711 1349
rect 7653 1309 7665 1343
rect 7699 1340 7711 1343
rect 8205 1343 8263 1349
rect 8205 1340 8217 1343
rect 7699 1312 8217 1340
rect 7699 1309 7711 1312
rect 7653 1303 7711 1309
rect 8205 1309 8217 1312
rect 8251 1340 8263 1343
rect 8757 1343 8815 1349
rect 8757 1340 8769 1343
rect 8251 1312 8769 1340
rect 8251 1309 8263 1312
rect 8205 1303 8263 1309
rect 8757 1309 8769 1312
rect 8803 1309 8815 1343
rect 8757 1303 8815 1309
rect 4341 1275 4399 1281
rect 4341 1241 4353 1275
rect 4387 1241 4399 1275
rect 4341 1235 4399 1241
rect 4985 1275 5043 1281
rect 4985 1241 4997 1275
rect 5031 1241 5043 1275
rect 4985 1235 5043 1241
rect 6362 1232 6368 1284
rect 6420 1232 6426 1284
rect 7745 1275 7803 1281
rect 7745 1241 7757 1275
rect 7791 1272 7803 1275
rect 8018 1272 8024 1284
rect 7791 1244 8024 1272
rect 7791 1241 7803 1244
rect 7745 1235 7803 1241
rect 8018 1232 8024 1244
rect 8076 1232 8082 1284
rect 8772 1272 8800 1303
rect 9122 1300 9128 1352
rect 9180 1340 9186 1352
rect 9217 1343 9275 1349
rect 9217 1340 9229 1343
rect 9180 1312 9229 1340
rect 9180 1300 9186 1312
rect 9217 1309 9229 1312
rect 9263 1309 9275 1343
rect 9217 1303 9275 1309
rect 9309 1343 9367 1349
rect 9309 1309 9321 1343
rect 9355 1340 9367 1343
rect 9490 1340 9496 1352
rect 9355 1312 9496 1340
rect 9355 1309 9367 1312
rect 9309 1303 9367 1309
rect 9324 1272 9352 1303
rect 9490 1300 9496 1312
rect 9548 1300 9554 1352
rect 8772 1244 9352 1272
rect 1673 1207 1731 1213
rect 1673 1173 1685 1207
rect 1719 1204 1731 1207
rect 1762 1204 1768 1216
rect 1719 1176 1768 1204
rect 1719 1173 1731 1176
rect 1673 1167 1731 1173
rect 1762 1164 1768 1176
rect 1820 1164 1826 1216
rect 2958 1164 2964 1216
rect 3016 1164 3022 1216
rect 5629 1207 5687 1213
rect 5629 1173 5641 1207
rect 5675 1204 5687 1207
rect 6178 1204 6184 1216
rect 5675 1176 6184 1204
rect 5675 1173 5687 1176
rect 5629 1167 5687 1173
rect 6178 1164 6184 1176
rect 6236 1164 6242 1216
rect 8478 1164 8484 1216
rect 8536 1204 8542 1216
rect 9600 1204 9628 1371
rect 9766 1368 9772 1420
rect 9824 1408 9830 1420
rect 10428 1417 10456 1448
rect 11532 1448 11836 1476
rect 9861 1411 9919 1417
rect 9861 1408 9873 1411
rect 9824 1380 9873 1408
rect 9824 1368 9830 1380
rect 9861 1377 9873 1380
rect 9907 1408 9919 1411
rect 10413 1411 10471 1417
rect 9907 1380 10364 1408
rect 9907 1377 9919 1380
rect 9861 1371 9919 1377
rect 9950 1300 9956 1352
rect 10008 1300 10014 1352
rect 10042 1300 10048 1352
rect 10100 1340 10106 1352
rect 10137 1343 10195 1349
rect 10137 1340 10149 1343
rect 10100 1312 10149 1340
rect 10100 1300 10106 1312
rect 10137 1309 10149 1312
rect 10183 1309 10195 1343
rect 10336 1340 10364 1380
rect 10413 1377 10425 1411
rect 10459 1377 10471 1411
rect 10413 1371 10471 1377
rect 11330 1368 11336 1420
rect 11388 1368 11394 1420
rect 11532 1417 11560 1448
rect 11517 1411 11575 1417
rect 11517 1377 11529 1411
rect 11563 1377 11575 1411
rect 11517 1371 11575 1377
rect 11698 1368 11704 1420
rect 11756 1368 11762 1420
rect 11808 1340 11836 1448
rect 12263 1445 12275 1479
rect 12309 1476 12321 1479
rect 12544 1476 12572 1504
rect 13265 1479 13323 1485
rect 13265 1476 13277 1479
rect 12309 1448 13277 1476
rect 12309 1445 12321 1448
rect 12263 1439 12321 1445
rect 13265 1445 13277 1448
rect 13311 1445 13323 1479
rect 13265 1439 13323 1445
rect 13357 1479 13415 1485
rect 13357 1445 13369 1479
rect 13403 1445 13415 1479
rect 13357 1439 13415 1445
rect 11974 1368 11980 1420
rect 12032 1368 12038 1420
rect 12066 1368 12072 1420
rect 12124 1368 12130 1420
rect 12180 1411 12238 1417
rect 12180 1377 12192 1411
rect 12226 1408 12238 1411
rect 12529 1411 12587 1417
rect 12529 1408 12541 1411
rect 12226 1380 12541 1408
rect 12226 1377 12238 1380
rect 12180 1371 12238 1377
rect 12529 1377 12541 1380
rect 12575 1377 12587 1411
rect 12529 1371 12587 1377
rect 12713 1411 12771 1417
rect 12713 1377 12725 1411
rect 12759 1408 12771 1411
rect 12802 1408 12808 1420
rect 12759 1380 12808 1408
rect 12759 1377 12771 1380
rect 12713 1371 12771 1377
rect 12728 1340 12756 1371
rect 12802 1368 12808 1380
rect 12860 1368 12866 1420
rect 12897 1411 12955 1417
rect 12897 1377 12909 1411
rect 12943 1377 12955 1411
rect 12897 1371 12955 1377
rect 10336 1312 11652 1340
rect 11808 1312 12756 1340
rect 12912 1340 12940 1371
rect 12986 1368 12992 1420
rect 13044 1368 13050 1420
rect 13078 1368 13084 1420
rect 13136 1408 13142 1420
rect 13372 1408 13400 1439
rect 13136 1380 13400 1408
rect 13136 1368 13142 1380
rect 13630 1368 13636 1420
rect 13688 1368 13694 1420
rect 13722 1368 13728 1420
rect 13780 1408 13786 1420
rect 13909 1411 13967 1417
rect 13909 1408 13921 1411
rect 13780 1380 13921 1408
rect 13780 1368 13786 1380
rect 13909 1377 13921 1380
rect 13955 1377 13967 1411
rect 13909 1371 13967 1377
rect 13354 1340 13360 1352
rect 12912 1312 13360 1340
rect 10137 1303 10195 1309
rect 9674 1232 9680 1284
rect 9732 1272 9738 1284
rect 9769 1275 9827 1281
rect 9769 1272 9781 1275
rect 9732 1244 9781 1272
rect 9732 1232 9738 1244
rect 9769 1241 9781 1244
rect 9815 1272 9827 1275
rect 9858 1272 9864 1284
rect 9815 1244 9864 1272
rect 9815 1241 9827 1244
rect 9769 1235 9827 1241
rect 9858 1232 9864 1244
rect 9916 1232 9922 1284
rect 9968 1272 9996 1300
rect 10229 1275 10287 1281
rect 10229 1272 10241 1275
rect 9968 1244 10241 1272
rect 10229 1241 10241 1244
rect 10275 1272 10287 1275
rect 10778 1272 10784 1284
rect 10275 1244 10784 1272
rect 10275 1241 10287 1244
rect 10229 1235 10287 1241
rect 10778 1232 10784 1244
rect 10836 1232 10842 1284
rect 10870 1232 10876 1284
rect 10928 1272 10934 1284
rect 11333 1275 11391 1281
rect 11333 1272 11345 1275
rect 10928 1244 11345 1272
rect 10928 1232 10934 1244
rect 11333 1241 11345 1244
rect 11379 1241 11391 1275
rect 11333 1235 11391 1241
rect 8536 1176 9628 1204
rect 9953 1207 10011 1213
rect 8536 1164 8542 1176
rect 9953 1173 9965 1207
rect 9999 1204 10011 1207
rect 10134 1204 10140 1216
rect 9999 1176 10140 1204
rect 9999 1173 10011 1176
rect 9953 1167 10011 1173
rect 10134 1164 10140 1176
rect 10192 1164 10198 1216
rect 10597 1207 10655 1213
rect 10597 1173 10609 1207
rect 10643 1204 10655 1207
rect 11514 1204 11520 1216
rect 10643 1176 11520 1204
rect 10643 1173 10655 1176
rect 10597 1167 10655 1173
rect 11514 1164 11520 1176
rect 11572 1164 11578 1216
rect 11624 1204 11652 1312
rect 13354 1300 13360 1312
rect 13412 1300 13418 1352
rect 14200 1340 14228 1516
rect 14292 1516 15294 1544
rect 14292 1417 14320 1516
rect 15282 1513 15294 1516
rect 15328 1513 15340 1547
rect 15282 1507 15340 1513
rect 15654 1504 15660 1556
rect 15712 1553 15718 1556
rect 15712 1544 15721 1553
rect 15712 1516 15757 1544
rect 15712 1507 15721 1516
rect 15712 1504 15718 1507
rect 16206 1504 16212 1556
rect 16264 1504 16270 1556
rect 18506 1544 18512 1556
rect 17144 1516 18512 1544
rect 14366 1436 14372 1488
rect 14424 1476 14430 1488
rect 14645 1479 14703 1485
rect 14645 1476 14657 1479
rect 14424 1448 14657 1476
rect 14424 1436 14430 1448
rect 14645 1445 14657 1448
rect 14691 1445 14703 1479
rect 14918 1476 14924 1488
rect 14645 1439 14703 1445
rect 14752 1448 14924 1476
rect 14277 1411 14335 1417
rect 14277 1377 14289 1411
rect 14323 1377 14335 1411
rect 14277 1371 14335 1377
rect 14461 1411 14519 1417
rect 14461 1377 14473 1411
rect 14507 1408 14519 1411
rect 14550 1408 14556 1420
rect 14507 1380 14556 1408
rect 14507 1377 14519 1380
rect 14461 1371 14519 1377
rect 14550 1368 14556 1380
rect 14608 1368 14614 1420
rect 14752 1417 14780 1448
rect 14918 1436 14924 1448
rect 14976 1436 14982 1488
rect 15013 1479 15071 1485
rect 15013 1445 15025 1479
rect 15059 1476 15071 1479
rect 15378 1476 15384 1488
rect 15059 1448 15384 1476
rect 15059 1445 15071 1448
rect 15013 1439 15071 1445
rect 15378 1436 15384 1448
rect 15436 1436 15442 1488
rect 15565 1479 15623 1485
rect 15565 1445 15577 1479
rect 15611 1476 15623 1479
rect 16224 1476 16252 1504
rect 17144 1476 17172 1516
rect 18506 1504 18512 1516
rect 18564 1504 18570 1556
rect 18690 1504 18696 1556
rect 18748 1544 18754 1556
rect 19153 1547 19211 1553
rect 19153 1544 19165 1547
rect 18748 1516 19165 1544
rect 18748 1504 18754 1516
rect 19153 1513 19165 1516
rect 19199 1513 19211 1547
rect 19153 1507 19211 1513
rect 19886 1504 19892 1556
rect 19944 1544 19950 1556
rect 22278 1544 22284 1556
rect 19944 1516 22284 1544
rect 19944 1504 19950 1516
rect 22278 1504 22284 1516
rect 22336 1504 22342 1556
rect 22370 1504 22376 1556
rect 22428 1544 22434 1556
rect 23290 1544 23296 1556
rect 22428 1516 23296 1544
rect 22428 1504 22434 1516
rect 23290 1504 23296 1516
rect 23348 1504 23354 1556
rect 15611 1448 16252 1476
rect 17052 1448 17172 1476
rect 17880 1448 20484 1476
rect 15611 1445 15623 1448
rect 15565 1439 15623 1445
rect 14737 1411 14795 1417
rect 14737 1377 14749 1411
rect 14783 1377 14795 1411
rect 14737 1371 14795 1377
rect 14829 1411 14887 1417
rect 14829 1377 14841 1411
rect 14875 1377 14887 1411
rect 14829 1371 14887 1377
rect 14844 1340 14872 1371
rect 15102 1368 15108 1420
rect 15160 1368 15166 1420
rect 15194 1368 15200 1420
rect 15252 1368 15258 1420
rect 15746 1408 15752 1420
rect 15297 1380 15752 1408
rect 15297 1340 15325 1380
rect 15746 1368 15752 1380
rect 15804 1368 15810 1420
rect 15838 1368 15844 1420
rect 15896 1368 15902 1420
rect 16114 1368 16120 1420
rect 16172 1408 16178 1420
rect 16209 1411 16267 1417
rect 16209 1408 16221 1411
rect 16172 1380 16221 1408
rect 16172 1368 16178 1380
rect 16209 1377 16221 1380
rect 16255 1377 16267 1411
rect 16209 1371 16267 1377
rect 16574 1368 16580 1420
rect 16632 1368 16638 1420
rect 17052 1417 17080 1448
rect 17037 1411 17095 1417
rect 17037 1408 17049 1411
rect 16684 1380 17049 1408
rect 14200 1312 15325 1340
rect 15562 1300 15568 1352
rect 15620 1340 15626 1352
rect 16684 1340 16712 1380
rect 17037 1377 17049 1380
rect 17083 1377 17095 1411
rect 17037 1371 17095 1377
rect 17126 1368 17132 1420
rect 17184 1368 17190 1420
rect 17880 1417 17908 1448
rect 17865 1411 17923 1417
rect 17865 1377 17877 1411
rect 17911 1377 17923 1411
rect 17865 1371 17923 1377
rect 18598 1368 18604 1420
rect 18656 1368 18662 1420
rect 18800 1417 18828 1448
rect 18785 1411 18843 1417
rect 18785 1377 18797 1411
rect 18831 1377 18843 1411
rect 18785 1371 18843 1377
rect 18966 1368 18972 1420
rect 19024 1368 19030 1420
rect 19058 1368 19064 1420
rect 19116 1368 19122 1420
rect 19702 1368 19708 1420
rect 19760 1368 19766 1420
rect 19794 1368 19800 1420
rect 19852 1368 19858 1420
rect 19996 1417 20024 1448
rect 19981 1411 20039 1417
rect 19981 1377 19993 1411
rect 20027 1377 20039 1411
rect 19981 1371 20039 1377
rect 20346 1368 20352 1420
rect 20404 1368 20410 1420
rect 20456 1408 20484 1448
rect 20714 1436 20720 1488
rect 20772 1476 20778 1488
rect 20901 1479 20959 1485
rect 20901 1476 20913 1479
rect 20772 1448 20913 1476
rect 20772 1436 20778 1448
rect 20901 1445 20913 1448
rect 20947 1445 20959 1479
rect 20901 1439 20959 1445
rect 21726 1436 21732 1488
rect 21784 1476 21790 1488
rect 22557 1479 22615 1485
rect 21784 1448 22508 1476
rect 21784 1436 21790 1448
rect 20456 1380 20760 1408
rect 15620 1312 16712 1340
rect 16761 1343 16819 1349
rect 15620 1300 15626 1312
rect 16761 1309 16773 1343
rect 16807 1340 16819 1343
rect 16850 1340 16856 1352
rect 16807 1312 16856 1340
rect 16807 1309 16819 1312
rect 16761 1303 16819 1309
rect 16850 1300 16856 1312
rect 16908 1300 16914 1352
rect 17313 1343 17371 1349
rect 17313 1309 17325 1343
rect 17359 1309 17371 1343
rect 17313 1303 17371 1309
rect 12342 1232 12348 1284
rect 12400 1272 12406 1284
rect 12529 1275 12587 1281
rect 12529 1272 12541 1275
rect 12400 1244 12541 1272
rect 12400 1232 12406 1244
rect 12529 1241 12541 1244
rect 12575 1241 12587 1275
rect 13541 1275 13599 1281
rect 13541 1272 13553 1275
rect 12529 1235 12587 1241
rect 13464 1244 13553 1272
rect 13078 1204 13084 1216
rect 11624 1176 13084 1204
rect 13078 1164 13084 1176
rect 13136 1164 13142 1216
rect 13265 1207 13323 1213
rect 13265 1173 13277 1207
rect 13311 1204 13323 1207
rect 13464 1204 13492 1244
rect 13541 1241 13553 1244
rect 13587 1241 13599 1275
rect 13541 1235 13599 1241
rect 14274 1232 14280 1284
rect 14332 1232 14338 1284
rect 14458 1232 14464 1284
rect 14516 1272 14522 1284
rect 17221 1275 17279 1281
rect 17221 1272 17233 1275
rect 14516 1244 17233 1272
rect 14516 1232 14522 1244
rect 17221 1241 17233 1244
rect 17267 1241 17279 1275
rect 17328 1272 17356 1303
rect 17586 1300 17592 1352
rect 17644 1300 17650 1352
rect 18984 1340 19012 1368
rect 19429 1343 19487 1349
rect 19429 1340 19441 1343
rect 17696 1312 19012 1340
rect 19306 1312 19441 1340
rect 17696 1272 17724 1312
rect 17328 1244 17724 1272
rect 17221 1235 17279 1241
rect 18598 1232 18604 1284
rect 18656 1232 18662 1284
rect 18690 1232 18696 1284
rect 18748 1272 18754 1284
rect 19306 1272 19334 1312
rect 19429 1309 19441 1312
rect 19475 1340 19487 1343
rect 19812 1340 19840 1368
rect 19475 1312 19840 1340
rect 19475 1309 19487 1312
rect 19429 1303 19487 1309
rect 20070 1300 20076 1352
rect 20128 1340 20134 1352
rect 20257 1343 20315 1349
rect 20257 1340 20269 1343
rect 20128 1312 20269 1340
rect 20128 1300 20134 1312
rect 20257 1309 20269 1312
rect 20303 1309 20315 1343
rect 20257 1303 20315 1309
rect 20438 1300 20444 1352
rect 20496 1300 20502 1352
rect 20622 1300 20628 1352
rect 20680 1300 20686 1352
rect 20732 1340 20760 1380
rect 20806 1368 20812 1420
rect 20864 1408 20870 1420
rect 21269 1411 21327 1417
rect 21269 1408 21281 1411
rect 20864 1380 21281 1408
rect 20864 1368 20870 1380
rect 21269 1377 21281 1380
rect 21315 1377 21327 1411
rect 21542 1408 21548 1420
rect 21269 1371 21327 1377
rect 21376 1380 21548 1408
rect 21376 1340 21404 1380
rect 21542 1368 21548 1380
rect 21600 1368 21606 1420
rect 22189 1411 22247 1417
rect 22189 1377 22201 1411
rect 22235 1408 22247 1411
rect 22370 1408 22376 1420
rect 22235 1380 22376 1408
rect 22235 1377 22247 1380
rect 22189 1371 22247 1377
rect 22370 1368 22376 1380
rect 22428 1368 22434 1420
rect 20732 1312 21404 1340
rect 21910 1300 21916 1352
rect 21968 1340 21974 1352
rect 22480 1349 22508 1448
rect 22557 1445 22569 1479
rect 22603 1476 22615 1479
rect 23014 1476 23020 1488
rect 22603 1448 23020 1476
rect 22603 1445 22615 1448
rect 22557 1439 22615 1445
rect 23014 1436 23020 1448
rect 23072 1436 23078 1488
rect 22833 1411 22891 1417
rect 22833 1377 22845 1411
rect 22879 1408 22891 1411
rect 22922 1408 22928 1420
rect 22879 1380 22928 1408
rect 22879 1377 22891 1380
rect 22833 1371 22891 1377
rect 22922 1368 22928 1380
rect 22980 1368 22986 1420
rect 22572 1349 22784 1351
rect 22281 1343 22339 1349
rect 22281 1340 22293 1343
rect 21968 1312 22293 1340
rect 21968 1300 21974 1312
rect 22281 1309 22293 1312
rect 22327 1309 22339 1343
rect 22281 1303 22339 1309
rect 22465 1343 22523 1349
rect 22465 1309 22477 1343
rect 22511 1309 22523 1343
rect 22465 1303 22523 1309
rect 22557 1343 22784 1349
rect 22557 1309 22569 1343
rect 22603 1340 22784 1343
rect 23382 1340 23388 1352
rect 22603 1323 23388 1340
rect 22603 1309 22615 1323
rect 22756 1312 23388 1323
rect 22557 1303 22615 1309
rect 23382 1300 23388 1312
rect 23440 1300 23446 1352
rect 18748 1244 19334 1272
rect 18748 1232 18754 1244
rect 19886 1232 19892 1284
rect 19944 1232 19950 1284
rect 20456 1272 20484 1300
rect 22373 1275 22431 1281
rect 22373 1272 22385 1275
rect 20456 1244 22385 1272
rect 22373 1241 22385 1244
rect 22419 1241 22431 1275
rect 22373 1235 22431 1241
rect 22741 1275 22799 1281
rect 22741 1241 22753 1275
rect 22787 1241 22799 1275
rect 22741 1235 22799 1241
rect 13311 1176 13492 1204
rect 13311 1173 13323 1176
rect 13265 1167 13323 1173
rect 13814 1164 13820 1216
rect 13872 1164 13878 1216
rect 15010 1164 15016 1216
rect 15068 1164 15074 1216
rect 15102 1164 15108 1216
rect 15160 1204 15166 1216
rect 16301 1207 16359 1213
rect 16301 1204 16313 1207
rect 15160 1176 16313 1204
rect 15160 1164 15166 1176
rect 16301 1173 16313 1176
rect 16347 1173 16359 1207
rect 16301 1167 16359 1173
rect 17678 1164 17684 1216
rect 17736 1164 17742 1216
rect 17770 1164 17776 1216
rect 17828 1164 17834 1216
rect 18322 1164 18328 1216
rect 18380 1204 18386 1216
rect 19058 1204 19064 1216
rect 18380 1176 19064 1204
rect 18380 1164 18386 1176
rect 19058 1164 19064 1176
rect 19116 1164 19122 1216
rect 19521 1207 19579 1213
rect 19521 1173 19533 1207
rect 19567 1204 19579 1207
rect 20070 1204 20076 1216
rect 19567 1176 20076 1204
rect 19567 1173 19579 1176
rect 19521 1167 19579 1173
rect 20070 1164 20076 1176
rect 20128 1164 20134 1216
rect 20165 1207 20223 1213
rect 20165 1173 20177 1207
rect 20211 1204 20223 1207
rect 20346 1204 20352 1216
rect 20211 1176 20352 1204
rect 20211 1173 20223 1176
rect 20165 1167 20223 1173
rect 20346 1164 20352 1176
rect 20404 1164 20410 1216
rect 20438 1164 20444 1216
rect 20496 1164 20502 1216
rect 20530 1164 20536 1216
rect 20588 1164 20594 1216
rect 20806 1164 20812 1216
rect 20864 1164 20870 1216
rect 20898 1164 20904 1216
rect 20956 1204 20962 1216
rect 22756 1204 22784 1235
rect 20956 1176 22784 1204
rect 20956 1164 20962 1176
rect 552 1114 23368 1136
rect 552 1062 1366 1114
rect 1418 1062 1430 1114
rect 1482 1062 1494 1114
rect 1546 1062 1558 1114
rect 1610 1062 1622 1114
rect 1674 1062 1686 1114
rect 1738 1062 7366 1114
rect 7418 1062 7430 1114
rect 7482 1062 7494 1114
rect 7546 1062 7558 1114
rect 7610 1062 7622 1114
rect 7674 1062 7686 1114
rect 7738 1062 13366 1114
rect 13418 1062 13430 1114
rect 13482 1062 13494 1114
rect 13546 1062 13558 1114
rect 13610 1062 13622 1114
rect 13674 1062 13686 1114
rect 13738 1062 19366 1114
rect 19418 1062 19430 1114
rect 19482 1062 19494 1114
rect 19546 1062 19558 1114
rect 19610 1062 19622 1114
rect 19674 1062 19686 1114
rect 19738 1062 23368 1114
rect 552 1040 23368 1062
rect 2501 1003 2559 1009
rect 2501 969 2513 1003
rect 2547 1000 2559 1003
rect 3326 1000 3332 1012
rect 2547 972 3332 1000
rect 2547 969 2559 972
rect 2501 963 2559 969
rect 3326 960 3332 972
rect 3384 960 3390 1012
rect 5905 1003 5963 1009
rect 5905 969 5917 1003
rect 5951 1000 5963 1003
rect 5994 1000 6000 1012
rect 5951 972 6000 1000
rect 5951 969 5963 972
rect 5905 963 5963 969
rect 5994 960 6000 972
rect 6052 960 6058 1012
rect 6086 960 6092 1012
rect 6144 1000 6150 1012
rect 6457 1003 6515 1009
rect 6457 1000 6469 1003
rect 6144 972 6469 1000
rect 6144 960 6150 972
rect 6457 969 6469 972
rect 6503 969 6515 1003
rect 6457 963 6515 969
rect 6822 960 6828 1012
rect 6880 960 6886 1012
rect 7834 960 7840 1012
rect 7892 1000 7898 1012
rect 7929 1003 7987 1009
rect 7929 1000 7941 1003
rect 7892 972 7941 1000
rect 7892 960 7898 972
rect 7929 969 7941 972
rect 7975 969 7987 1003
rect 7929 963 7987 969
rect 8389 1003 8447 1009
rect 8389 969 8401 1003
rect 8435 1000 8447 1003
rect 8478 1000 8484 1012
rect 8435 972 8484 1000
rect 8435 969 8447 972
rect 8389 963 8447 969
rect 8478 960 8484 972
rect 8536 960 8542 1012
rect 9217 1003 9275 1009
rect 9217 969 9229 1003
rect 9263 1000 9275 1003
rect 9950 1000 9956 1012
rect 9263 972 9956 1000
rect 9263 969 9275 972
rect 9217 963 9275 969
rect 9950 960 9956 972
rect 10008 960 10014 1012
rect 11330 960 11336 1012
rect 11388 960 11394 1012
rect 11514 960 11520 1012
rect 11572 1000 11578 1012
rect 14182 1000 14188 1012
rect 11572 972 14188 1000
rect 11572 960 11578 972
rect 14182 960 14188 972
rect 14240 960 14246 1012
rect 14461 1003 14519 1009
rect 14461 969 14473 1003
rect 14507 1000 14519 1003
rect 15010 1000 15016 1012
rect 14507 972 15016 1000
rect 14507 969 14519 972
rect 14461 963 14519 969
rect 15010 960 15016 972
rect 15068 960 15074 1012
rect 16574 960 16580 1012
rect 16632 1000 16638 1012
rect 16669 1003 16727 1009
rect 16669 1000 16681 1003
rect 16632 972 16681 1000
rect 16632 960 16638 972
rect 16669 969 16681 972
rect 16715 969 16727 1003
rect 20254 1000 20260 1012
rect 16669 963 16727 969
rect 16776 972 20260 1000
rect 2133 935 2191 941
rect 2133 901 2145 935
rect 2179 932 2191 935
rect 2590 932 2596 944
rect 2179 904 2596 932
rect 2179 901 2191 904
rect 2133 895 2191 901
rect 2590 892 2596 904
rect 2648 892 2654 944
rect 3050 932 3056 944
rect 2746 904 3056 932
rect 2746 864 2774 904
rect 3050 892 3056 904
rect 3108 892 3114 944
rect 3605 935 3663 941
rect 3605 901 3617 935
rect 3651 932 3663 935
rect 4062 932 4068 944
rect 3651 904 4068 932
rect 3651 901 3663 904
rect 3605 895 3663 901
rect 4062 892 4068 904
rect 4120 892 4126 944
rect 4709 935 4767 941
rect 4709 901 4721 935
rect 4755 932 4767 935
rect 5166 932 5172 944
rect 4755 904 5172 932
rect 4755 901 4767 904
rect 4709 895 4767 901
rect 5166 892 5172 904
rect 5224 892 5230 944
rect 7098 932 7104 944
rect 5276 904 7104 932
rect 2332 836 2774 864
rect 1210 756 1216 808
rect 1268 756 1274 808
rect 1581 799 1639 805
rect 1581 765 1593 799
rect 1627 796 1639 799
rect 1762 796 1768 808
rect 1627 768 1768 796
rect 1627 765 1639 768
rect 1581 759 1639 765
rect 1762 756 1768 768
rect 1820 756 1826 808
rect 1946 756 1952 808
rect 2004 756 2010 808
rect 2332 805 2360 836
rect 2317 799 2375 805
rect 2317 765 2329 799
rect 2363 765 2375 799
rect 2317 759 2375 765
rect 2685 799 2743 805
rect 2685 765 2697 799
rect 2731 765 2743 799
rect 2685 759 2743 765
rect 3053 799 3111 805
rect 3053 765 3065 799
rect 3099 796 3111 799
rect 3329 799 3387 805
rect 3329 796 3341 799
rect 3099 768 3341 796
rect 3099 765 3111 768
rect 3053 759 3111 765
rect 3329 765 3341 768
rect 3375 765 3387 799
rect 3329 759 3387 765
rect 2700 728 2728 759
rect 3418 756 3424 808
rect 3476 756 3482 808
rect 3789 799 3847 805
rect 3789 765 3801 799
rect 3835 765 3847 799
rect 3789 759 3847 765
rect 3436 728 3464 756
rect 2700 700 3464 728
rect 3804 728 3832 759
rect 4154 756 4160 808
rect 4212 756 4218 808
rect 4522 756 4528 808
rect 4580 756 4586 808
rect 4890 756 4896 808
rect 4948 756 4954 808
rect 5276 805 5304 904
rect 7098 892 7104 904
rect 7156 892 7162 944
rect 7377 935 7435 941
rect 7377 901 7389 935
rect 7423 932 7435 935
rect 8849 935 8907 941
rect 7423 904 8708 932
rect 7423 901 7435 904
rect 7377 895 7435 901
rect 7009 867 7067 873
rect 7009 864 7021 867
rect 5644 836 7021 864
rect 5644 805 5672 836
rect 7009 833 7021 836
rect 7055 833 7067 867
rect 7009 827 7067 833
rect 7745 867 7803 873
rect 7745 833 7757 867
rect 7791 864 7803 867
rect 7926 864 7932 876
rect 7791 836 7932 864
rect 7791 833 7803 836
rect 7745 827 7803 833
rect 7926 824 7932 836
rect 7984 824 7990 876
rect 5261 799 5319 805
rect 5261 765 5273 799
rect 5307 765 5319 799
rect 5261 759 5319 765
rect 5629 799 5687 805
rect 5629 765 5641 799
rect 5675 765 5687 799
rect 5629 759 5687 765
rect 5902 756 5908 808
rect 5960 756 5966 808
rect 6178 756 6184 808
rect 6236 796 6242 808
rect 6365 799 6423 805
rect 6365 796 6377 799
rect 6236 768 6377 796
rect 6236 756 6242 768
rect 6365 765 6377 768
rect 6411 765 6423 799
rect 6365 759 6423 765
rect 7098 756 7104 808
rect 7156 756 7162 808
rect 7190 756 7196 808
rect 7248 756 7254 808
rect 7469 799 7527 805
rect 7469 765 7481 799
rect 7515 796 7527 799
rect 7834 796 7840 808
rect 7515 768 7840 796
rect 7515 765 7527 768
rect 7469 759 7527 765
rect 7834 756 7840 768
rect 7892 756 7898 808
rect 8021 799 8079 805
rect 8021 765 8033 799
rect 8067 796 8079 799
rect 8110 796 8116 808
rect 8067 768 8116 796
rect 8067 765 8079 768
rect 8021 759 8079 765
rect 8110 756 8116 768
rect 8168 756 8174 808
rect 8680 805 8708 904
rect 8849 901 8861 935
rect 8895 932 8907 935
rect 9582 932 9588 944
rect 8895 904 9588 932
rect 8895 901 8907 904
rect 8849 895 8907 901
rect 9582 892 9588 904
rect 9640 892 9646 944
rect 10321 935 10379 941
rect 10321 901 10333 935
rect 10367 932 10379 935
rect 10962 932 10968 944
rect 10367 904 10968 932
rect 10367 901 10379 904
rect 10321 895 10379 901
rect 10962 892 10968 904
rect 11020 892 11026 944
rect 11422 892 11428 944
rect 11480 932 11486 944
rect 11701 935 11759 941
rect 11701 932 11713 935
rect 11480 904 11713 932
rect 11480 892 11486 904
rect 11701 901 11713 904
rect 11747 901 11759 935
rect 11701 895 11759 901
rect 14918 892 14924 944
rect 14976 932 14982 944
rect 15473 935 15531 941
rect 15473 932 15485 935
rect 14976 904 15485 932
rect 14976 892 14982 904
rect 15473 901 15485 904
rect 15519 901 15531 935
rect 15473 895 15531 901
rect 9306 824 9312 876
rect 9364 864 9370 876
rect 10686 864 10692 876
rect 9364 836 10692 864
rect 9364 824 9370 836
rect 10686 824 10692 836
rect 10744 824 10750 876
rect 11517 867 11575 873
rect 10796 836 11192 864
rect 8573 799 8631 805
rect 8573 765 8585 799
rect 8619 765 8631 799
rect 8573 759 8631 765
rect 8665 799 8723 805
rect 8665 765 8677 799
rect 8711 765 8723 799
rect 8665 759 8723 765
rect 4982 728 4988 740
rect 3804 700 4988 728
rect 4982 688 4988 700
rect 5040 688 5046 740
rect 5534 728 5540 740
rect 5092 700 5540 728
rect 1029 663 1087 669
rect 1029 629 1041 663
rect 1075 660 1087 663
rect 1118 660 1124 672
rect 1075 632 1124 660
rect 1075 629 1087 632
rect 1029 623 1087 629
rect 1118 620 1124 632
rect 1176 620 1182 672
rect 1397 663 1455 669
rect 1397 629 1409 663
rect 1443 660 1455 663
rect 1486 660 1492 672
rect 1443 632 1492 660
rect 1443 629 1455 632
rect 1397 623 1455 629
rect 1486 620 1492 632
rect 1544 620 1550 672
rect 1765 663 1823 669
rect 1765 629 1777 663
rect 1811 660 1823 663
rect 1854 660 1860 672
rect 1811 632 1860 660
rect 1811 629 1823 632
rect 1765 623 1823 629
rect 1854 620 1860 632
rect 1912 620 1918 672
rect 2869 663 2927 669
rect 2869 629 2881 663
rect 2915 660 2927 663
rect 3694 660 3700 672
rect 2915 632 3700 660
rect 2915 629 2927 632
rect 2869 623 2927 629
rect 3694 620 3700 632
rect 3752 620 3758 672
rect 3973 663 4031 669
rect 3973 629 3985 663
rect 4019 660 4031 663
rect 4246 660 4252 672
rect 4019 632 4252 660
rect 4019 629 4031 632
rect 3973 623 4031 629
rect 4246 620 4252 632
rect 4304 620 4310 672
rect 4341 663 4399 669
rect 4341 629 4353 663
rect 4387 660 4399 663
rect 4798 660 4804 672
rect 4387 632 4804 660
rect 4387 629 4399 632
rect 4341 623 4399 629
rect 4798 620 4804 632
rect 4856 620 4862 672
rect 5092 669 5120 700
rect 5534 688 5540 700
rect 5592 688 5598 740
rect 6089 731 6147 737
rect 6089 697 6101 731
rect 6135 728 6147 731
rect 6730 728 6736 740
rect 6135 700 6736 728
rect 6135 697 6147 700
rect 6089 691 6147 697
rect 6730 688 6736 700
rect 6788 688 6794 740
rect 8588 728 8616 759
rect 8846 756 8852 808
rect 8904 796 8910 808
rect 9033 799 9091 805
rect 9033 796 9045 799
rect 8904 768 9045 796
rect 8904 756 8910 768
rect 9033 765 9045 768
rect 9079 765 9091 799
rect 9033 759 9091 765
rect 9401 799 9459 805
rect 9401 765 9413 799
rect 9447 765 9459 799
rect 9401 759 9459 765
rect 9122 728 9128 740
rect 7668 700 8524 728
rect 8588 700 9128 728
rect 5077 663 5135 669
rect 5077 629 5089 663
rect 5123 629 5135 663
rect 5077 623 5135 629
rect 5445 663 5503 669
rect 5445 629 5457 663
rect 5491 660 5503 663
rect 5810 660 5816 672
rect 5491 632 5816 660
rect 5491 629 5503 632
rect 5445 623 5503 629
rect 5810 620 5816 632
rect 5868 620 5874 672
rect 7668 669 7696 700
rect 7653 663 7711 669
rect 7653 629 7665 663
rect 7699 629 7711 663
rect 7653 623 7711 629
rect 7742 620 7748 672
rect 7800 620 7806 672
rect 8496 660 8524 700
rect 9122 688 9128 700
rect 9180 688 9186 740
rect 9416 660 9444 759
rect 9766 756 9772 808
rect 9824 756 9830 808
rect 10134 756 10140 808
rect 10192 756 10198 808
rect 10796 805 10824 836
rect 10781 799 10839 805
rect 10781 765 10793 799
rect 10827 765 10839 799
rect 10781 759 10839 765
rect 11054 756 11060 808
rect 11112 756 11118 808
rect 11164 796 11192 836
rect 11517 833 11529 867
rect 11563 864 11575 867
rect 13170 864 13176 876
rect 11563 836 11744 864
rect 11563 833 11575 836
rect 11517 827 11575 833
rect 11716 808 11744 836
rect 11808 836 13176 864
rect 11164 768 11468 796
rect 10612 700 11284 728
rect 8496 632 9444 660
rect 9585 663 9643 669
rect 9585 629 9597 663
rect 9631 660 9643 663
rect 9858 660 9864 672
rect 9631 632 9864 660
rect 9631 629 9643 632
rect 9585 623 9643 629
rect 9858 620 9864 632
rect 9916 620 9922 672
rect 9953 663 10011 669
rect 9953 629 9965 663
rect 9999 660 10011 663
rect 10226 660 10232 672
rect 9999 632 10232 660
rect 9999 629 10011 632
rect 9953 623 10011 629
rect 10226 620 10232 632
rect 10284 620 10290 672
rect 10612 669 10640 700
rect 10597 663 10655 669
rect 10597 629 10609 663
rect 10643 629 10655 663
rect 10597 623 10655 629
rect 11146 620 11152 672
rect 11204 620 11210 672
rect 11256 660 11284 700
rect 11330 688 11336 740
rect 11388 688 11394 740
rect 11440 728 11468 768
rect 11698 756 11704 808
rect 11756 756 11762 808
rect 11808 805 11836 836
rect 13170 824 13176 836
rect 13228 824 13234 876
rect 14277 867 14335 873
rect 14277 833 14289 867
rect 14323 864 14335 867
rect 14366 864 14372 876
rect 14323 836 14372 864
rect 14323 833 14335 836
rect 14277 827 14335 833
rect 14366 824 14372 836
rect 14424 824 14430 876
rect 16776 864 16804 972
rect 20254 960 20260 972
rect 20312 960 20318 1012
rect 21818 960 21824 1012
rect 21876 960 21882 1012
rect 22925 1003 22983 1009
rect 22925 1000 22937 1003
rect 21928 972 22937 1000
rect 15304 836 16804 864
rect 17604 904 19104 932
rect 11793 799 11851 805
rect 11793 765 11805 799
rect 11839 765 11851 799
rect 11793 759 11851 765
rect 11882 756 11888 808
rect 11940 756 11946 808
rect 12529 799 12587 805
rect 12529 765 12541 799
rect 12575 765 12587 799
rect 12529 759 12587 765
rect 11514 728 11520 740
rect 11440 700 11520 728
rect 11514 688 11520 700
rect 11572 688 11578 740
rect 12544 728 12572 759
rect 12618 756 12624 808
rect 12676 756 12682 808
rect 13262 756 13268 808
rect 13320 756 13326 808
rect 13814 756 13820 808
rect 13872 756 13878 808
rect 14185 799 14243 805
rect 14185 765 14197 799
rect 14231 796 14243 799
rect 14458 796 14464 808
rect 14231 768 14464 796
rect 14231 765 14243 768
rect 14185 759 14243 765
rect 14458 756 14464 768
rect 14516 756 14522 808
rect 14550 756 14556 808
rect 14608 756 14614 808
rect 14642 756 14648 808
rect 14700 756 14706 808
rect 15304 805 15332 836
rect 15948 805 15976 836
rect 15289 799 15347 805
rect 15289 765 15301 799
rect 15335 765 15347 799
rect 15289 759 15347 765
rect 15657 799 15715 805
rect 15657 765 15669 799
rect 15703 796 15715 799
rect 15841 799 15899 805
rect 15841 796 15853 799
rect 15703 768 15853 796
rect 15703 765 15715 768
rect 15657 759 15715 765
rect 15841 765 15853 768
rect 15887 765 15899 799
rect 15841 759 15899 765
rect 15933 799 15991 805
rect 15933 765 15945 799
rect 15979 765 15991 799
rect 15933 759 15991 765
rect 16206 756 16212 808
rect 16264 796 16270 808
rect 16485 799 16543 805
rect 16485 796 16497 799
rect 16264 768 16497 796
rect 16264 756 16270 768
rect 16485 765 16497 768
rect 16531 765 16543 799
rect 16485 759 16543 765
rect 16669 799 16727 805
rect 16669 765 16681 799
rect 16715 796 16727 799
rect 16758 796 16764 808
rect 16715 768 16764 796
rect 16715 765 16727 768
rect 16669 759 16727 765
rect 16758 756 16764 768
rect 16816 756 16822 808
rect 17604 796 17632 904
rect 17678 824 17684 876
rect 17736 864 17742 876
rect 19076 864 19104 904
rect 19150 892 19156 944
rect 19208 932 19214 944
rect 19613 935 19671 941
rect 19613 932 19625 935
rect 19208 904 19625 932
rect 19208 892 19214 904
rect 19613 901 19625 904
rect 19659 901 19671 935
rect 19613 895 19671 901
rect 19794 892 19800 944
rect 19852 932 19858 944
rect 19889 935 19947 941
rect 19889 932 19901 935
rect 19852 904 19901 932
rect 19852 892 19858 904
rect 19889 901 19901 904
rect 19935 901 19947 935
rect 19889 895 19947 901
rect 20438 892 20444 944
rect 20496 932 20502 944
rect 20901 935 20959 941
rect 20901 932 20913 935
rect 20496 904 20913 932
rect 20496 892 20502 904
rect 20901 901 20913 904
rect 20947 901 20959 935
rect 20901 895 20959 901
rect 20990 892 20996 944
rect 21048 932 21054 944
rect 21048 904 21404 932
rect 21048 892 21054 904
rect 19978 864 19984 876
rect 17736 836 18184 864
rect 19076 836 19984 864
rect 17736 824 17742 836
rect 17773 799 17831 805
rect 17773 796 17785 799
rect 17604 768 17785 796
rect 17773 765 17785 768
rect 17819 765 17831 799
rect 17773 759 17831 765
rect 17862 756 17868 808
rect 17920 756 17926 808
rect 18156 805 18184 836
rect 19978 824 19984 836
rect 20036 824 20042 876
rect 20257 867 20315 873
rect 20257 833 20269 867
rect 20303 864 20315 867
rect 20303 836 20484 864
rect 20303 833 20315 836
rect 20257 827 20315 833
rect 18141 799 18199 805
rect 18141 765 18153 799
rect 18187 765 18199 799
rect 18141 759 18199 765
rect 18693 799 18751 805
rect 18693 765 18705 799
rect 18739 765 18751 799
rect 18693 759 18751 765
rect 12710 728 12716 740
rect 12544 700 12716 728
rect 12710 688 12716 700
rect 12768 728 12774 740
rect 14277 731 14335 737
rect 14277 728 14289 731
rect 12768 700 14289 728
rect 12768 688 12774 700
rect 14277 697 14289 700
rect 14323 697 14335 731
rect 14277 691 14335 697
rect 14366 688 14372 740
rect 14424 728 14430 740
rect 18708 728 18736 759
rect 19058 756 19064 808
rect 19116 756 19122 808
rect 19242 756 19248 808
rect 19300 796 19306 808
rect 19429 799 19487 805
rect 19429 796 19441 799
rect 19300 768 19441 796
rect 19300 756 19306 768
rect 19429 765 19441 768
rect 19475 765 19487 799
rect 19429 759 19487 765
rect 19794 756 19800 808
rect 19852 756 19858 808
rect 20073 799 20131 805
rect 20073 765 20085 799
rect 20119 796 20131 799
rect 20162 796 20168 808
rect 20119 768 20168 796
rect 20119 765 20131 768
rect 20073 759 20131 765
rect 20162 756 20168 768
rect 20220 756 20226 808
rect 20346 756 20352 808
rect 20404 756 20410 808
rect 20456 796 20484 836
rect 20530 824 20536 876
rect 20588 864 20594 876
rect 21376 864 21404 904
rect 21726 892 21732 944
rect 21784 932 21790 944
rect 21928 932 21956 972
rect 22925 969 22937 972
rect 22971 969 22983 1003
rect 22925 963 22983 969
rect 22189 935 22247 941
rect 22189 932 22201 935
rect 21784 904 21956 932
rect 22066 904 22201 932
rect 21784 892 21790 904
rect 22066 864 22094 904
rect 22189 901 22201 904
rect 22235 901 22247 935
rect 22189 895 22247 901
rect 20588 836 21312 864
rect 21376 836 22094 864
rect 20588 824 20594 836
rect 20456 768 20668 796
rect 14424 700 15148 728
rect 14424 688 14430 700
rect 11422 660 11428 672
rect 11256 632 11428 660
rect 11422 620 11428 632
rect 11480 620 11486 672
rect 11790 620 11796 672
rect 11848 660 11854 672
rect 12069 663 12127 669
rect 12069 660 12081 663
rect 11848 632 12081 660
rect 11848 620 11854 632
rect 12069 629 12081 632
rect 12115 629 12127 663
rect 12069 623 12127 629
rect 12158 620 12164 672
rect 12216 660 12222 672
rect 12345 663 12403 669
rect 12345 660 12357 663
rect 12216 632 12357 660
rect 12216 620 12222 632
rect 12345 629 12357 632
rect 12391 629 12403 663
rect 12345 623 12403 629
rect 12526 620 12532 672
rect 12584 660 12590 672
rect 12805 663 12863 669
rect 12805 660 12817 663
rect 12584 632 12817 660
rect 12584 620 12590 632
rect 12805 629 12817 632
rect 12851 629 12863 663
rect 12805 623 12863 629
rect 12894 620 12900 672
rect 12952 660 12958 672
rect 13081 663 13139 669
rect 13081 660 13093 663
rect 12952 632 13093 660
rect 12952 620 12958 632
rect 13081 629 13093 632
rect 13127 629 13139 663
rect 13081 623 13139 629
rect 13262 620 13268 672
rect 13320 660 13326 672
rect 13633 663 13691 669
rect 13633 660 13645 663
rect 13320 632 13645 660
rect 13320 620 13326 632
rect 13633 629 13645 632
rect 13679 629 13691 663
rect 13633 623 13691 629
rect 13722 620 13728 672
rect 13780 660 13786 672
rect 14001 663 14059 669
rect 14001 660 14013 663
rect 13780 632 14013 660
rect 13780 620 13786 632
rect 14001 629 14013 632
rect 14047 629 14059 663
rect 14001 623 14059 629
rect 14090 620 14096 672
rect 14148 660 14154 672
rect 15120 669 15148 700
rect 18064 700 18736 728
rect 14829 663 14887 669
rect 14829 660 14841 663
rect 14148 632 14841 660
rect 14148 620 14154 632
rect 14829 629 14841 632
rect 14875 629 14887 663
rect 14829 623 14887 629
rect 15105 663 15163 669
rect 15105 629 15117 663
rect 15151 629 15163 663
rect 15105 623 15163 629
rect 17678 620 17684 672
rect 17736 620 17742 672
rect 18064 669 18092 700
rect 18782 688 18788 740
rect 18840 728 18846 740
rect 18840 700 19288 728
rect 18840 688 18846 700
rect 18049 663 18107 669
rect 18049 629 18061 663
rect 18095 629 18107 663
rect 18049 623 18107 629
rect 18138 620 18144 672
rect 18196 660 18202 672
rect 18325 663 18383 669
rect 18325 660 18337 663
rect 18196 632 18337 660
rect 18196 620 18202 632
rect 18325 629 18337 632
rect 18371 629 18383 663
rect 18325 623 18383 629
rect 18414 620 18420 672
rect 18472 660 18478 672
rect 19260 669 19288 700
rect 19518 688 19524 740
rect 19576 728 19582 740
rect 20640 728 20668 768
rect 20714 756 20720 808
rect 20772 756 20778 808
rect 21284 805 21312 836
rect 21269 799 21327 805
rect 21269 765 21281 799
rect 21315 765 21327 799
rect 21269 759 21327 765
rect 21637 799 21695 805
rect 21637 765 21649 799
rect 21683 765 21695 799
rect 21637 759 21695 765
rect 21652 728 21680 759
rect 21910 756 21916 808
rect 21968 796 21974 808
rect 22005 799 22063 805
rect 22005 796 22017 799
rect 21968 768 22017 796
rect 21968 756 21974 768
rect 22005 765 22017 768
rect 22051 765 22063 799
rect 22005 759 22063 765
rect 22186 756 22192 808
rect 22244 796 22250 808
rect 22373 799 22431 805
rect 22373 796 22385 799
rect 22244 768 22385 796
rect 22244 756 22250 768
rect 22373 765 22385 768
rect 22419 765 22431 799
rect 22373 759 22431 765
rect 22462 756 22468 808
rect 22520 796 22526 808
rect 22741 799 22799 805
rect 22741 796 22753 799
rect 22520 768 22753 796
rect 22520 756 22526 768
rect 22741 765 22753 768
rect 22787 796 22799 799
rect 23106 796 23112 808
rect 22787 768 23112 796
rect 22787 765 22799 768
rect 22741 759 22799 765
rect 23106 756 23112 768
rect 23164 756 23170 808
rect 19576 700 20576 728
rect 20640 700 21680 728
rect 22066 700 22600 728
rect 19576 688 19582 700
rect 20548 669 20576 700
rect 18877 663 18935 669
rect 18877 660 18889 663
rect 18472 632 18889 660
rect 18472 620 18478 632
rect 18877 629 18889 632
rect 18923 629 18935 663
rect 18877 623 18935 629
rect 19245 663 19303 669
rect 19245 629 19257 663
rect 19291 629 19303 663
rect 19245 623 19303 629
rect 20533 663 20591 669
rect 20533 629 20545 663
rect 20579 629 20591 663
rect 20533 623 20591 629
rect 20622 620 20628 672
rect 20680 660 20686 672
rect 21453 663 21511 669
rect 21453 660 21465 663
rect 20680 632 21465 660
rect 20680 620 20686 632
rect 21453 629 21465 632
rect 21499 629 21511 663
rect 21453 623 21511 629
rect 21542 620 21548 672
rect 21600 660 21606 672
rect 22066 660 22094 700
rect 22572 669 22600 700
rect 21600 632 22094 660
rect 22557 663 22615 669
rect 21600 620 21606 632
rect 22557 629 22569 663
rect 22603 629 22615 663
rect 22557 623 22615 629
rect 552 570 23368 592
rect 552 518 4366 570
rect 4418 518 4430 570
rect 4482 518 4494 570
rect 4546 518 4558 570
rect 4610 518 4622 570
rect 4674 518 4686 570
rect 4738 518 10366 570
rect 10418 518 10430 570
rect 10482 518 10494 570
rect 10546 518 10558 570
rect 10610 518 10622 570
rect 10674 518 10686 570
rect 10738 518 16366 570
rect 16418 518 16430 570
rect 16482 518 16494 570
rect 16546 518 16558 570
rect 16610 518 16622 570
rect 16674 518 16686 570
rect 16738 518 22366 570
rect 22418 518 22430 570
rect 22482 518 22494 570
rect 22546 518 22558 570
rect 22610 518 22622 570
rect 22674 518 22686 570
rect 22738 518 23368 570
rect 552 496 23368 518
rect 7190 416 7196 468
rect 7248 456 7254 468
rect 9674 456 9680 468
rect 7248 428 9680 456
rect 7248 416 7254 428
rect 9674 416 9680 428
rect 9732 416 9738 468
rect 9858 416 9864 468
rect 9916 456 9922 468
rect 10410 456 10416 468
rect 9916 428 10416 456
rect 9916 416 9922 428
rect 10410 416 10416 428
rect 10468 416 10474 468
rect 10594 416 10600 468
rect 10652 416 10658 468
rect 11146 416 11152 468
rect 11204 456 11210 468
rect 12066 456 12072 468
rect 11204 428 12072 456
rect 11204 416 11210 428
rect 12066 416 12072 428
rect 12124 416 12130 468
rect 17770 456 17776 468
rect 12176 428 17776 456
rect 1210 348 1216 400
rect 1268 388 1274 400
rect 7742 388 7748 400
rect 1268 360 7748 388
rect 1268 348 1274 360
rect 7742 348 7748 360
rect 7800 348 7806 400
rect 9306 388 9312 400
rect 7852 360 9312 388
rect 3050 280 3056 332
rect 3108 320 3114 332
rect 7852 320 7880 360
rect 9306 348 9312 360
rect 9364 348 9370 400
rect 10226 348 10232 400
rect 10284 388 10290 400
rect 10612 388 10640 416
rect 10284 360 10640 388
rect 10284 348 10290 360
rect 10778 348 10784 400
rect 10836 388 10842 400
rect 12176 388 12204 428
rect 17770 416 17776 428
rect 17828 416 17834 468
rect 17862 416 17868 468
rect 17920 456 17926 468
rect 18690 456 18696 468
rect 17920 428 18696 456
rect 17920 416 17926 428
rect 18690 416 18696 428
rect 18748 456 18754 468
rect 19794 456 19800 468
rect 18748 428 19800 456
rect 18748 416 18754 428
rect 19794 416 19800 428
rect 19852 416 19858 468
rect 19978 416 19984 468
rect 20036 456 20042 468
rect 20438 456 20444 468
rect 20036 428 20444 456
rect 20036 416 20042 428
rect 20438 416 20444 428
rect 20496 416 20502 468
rect 10836 360 12204 388
rect 10836 348 10842 360
rect 12986 348 12992 400
rect 13044 388 13050 400
rect 15102 388 15108 400
rect 13044 360 15108 388
rect 13044 348 13050 360
rect 15102 348 15108 360
rect 15160 348 15166 400
rect 17678 348 17684 400
rect 17736 388 17742 400
rect 22186 388 22192 400
rect 17736 360 22192 388
rect 17736 348 17742 360
rect 22186 348 22192 360
rect 22244 348 22250 400
rect 3108 292 7880 320
rect 3108 280 3114 292
rect 8110 280 8116 332
rect 8168 320 8174 332
rect 10042 320 10048 332
rect 8168 292 10048 320
rect 8168 280 8174 292
rect 10042 280 10048 292
rect 10100 280 10106 332
rect 14274 320 14280 332
rect 11624 292 14280 320
rect 3418 212 3424 264
rect 3476 252 3482 264
rect 11624 252 11652 292
rect 14274 280 14280 292
rect 14332 280 14338 332
rect 14550 280 14556 332
rect 14608 320 14614 332
rect 15562 320 15568 332
rect 14608 292 15568 320
rect 14608 280 14614 292
rect 15562 280 15568 292
rect 15620 280 15626 332
rect 18874 280 18880 332
rect 18932 320 18938 332
rect 20898 320 20904 332
rect 18932 292 20904 320
rect 18932 280 18938 292
rect 20898 280 20904 292
rect 20956 280 20962 332
rect 3476 224 11652 252
rect 3476 212 3482 224
rect 11698 212 11704 264
rect 11756 252 11762 264
rect 11756 224 13676 252
rect 11756 212 11762 224
rect 1946 144 1952 196
rect 2004 184 2010 196
rect 2004 156 2774 184
rect 2004 144 2010 156
rect 2746 48 2774 156
rect 4982 144 4988 196
rect 5040 184 5046 196
rect 12986 184 12992 196
rect 5040 156 12992 184
rect 5040 144 5046 156
rect 12986 144 12992 156
rect 13044 144 13050 196
rect 9122 76 9128 128
rect 9180 116 9186 128
rect 12066 116 12072 128
rect 9180 88 12072 116
rect 9180 76 9186 88
rect 12066 76 12072 88
rect 12124 76 12130 128
rect 13648 116 13676 224
rect 16850 212 16856 264
rect 16908 252 16914 264
rect 20806 252 20812 264
rect 16908 224 20812 252
rect 16908 212 16914 224
rect 20806 212 20812 224
rect 20864 212 20870 264
rect 18966 144 18972 196
rect 19024 184 19030 196
rect 23382 184 23388 196
rect 19024 156 23388 184
rect 19024 144 19030 156
rect 23382 144 23388 156
rect 23440 144 23446 196
rect 13648 88 14964 116
rect 12250 48 12256 60
rect 2746 20 12256 48
rect 12250 8 12256 20
rect 12308 8 12314 60
rect 14936 48 14964 88
rect 15194 76 15200 128
rect 15252 116 15258 128
rect 20070 116 20076 128
rect 15252 88 20076 116
rect 15252 76 15258 88
rect 20070 76 20076 88
rect 20128 76 20134 128
rect 20162 48 20168 60
rect 14936 20 20168 48
rect 20162 8 20168 20
rect 20220 8 20226 60
<< via1 >>
rect 2228 23604 2280 23656
rect 17960 23672 18012 23724
rect 4160 23536 4212 23588
rect 17224 23604 17276 23656
rect 6092 23468 6144 23520
rect 20076 23468 20128 23520
rect 4366 23366 4418 23418
rect 4430 23366 4482 23418
rect 4494 23366 4546 23418
rect 4558 23366 4610 23418
rect 4622 23366 4674 23418
rect 4686 23366 4738 23418
rect 10366 23366 10418 23418
rect 10430 23366 10482 23418
rect 10494 23366 10546 23418
rect 10558 23366 10610 23418
rect 10622 23366 10674 23418
rect 10686 23366 10738 23418
rect 16366 23366 16418 23418
rect 16430 23366 16482 23418
rect 16494 23366 16546 23418
rect 16558 23366 16610 23418
rect 16622 23366 16674 23418
rect 16686 23366 16738 23418
rect 22366 23366 22418 23418
rect 22430 23366 22482 23418
rect 22494 23366 22546 23418
rect 22558 23366 22610 23418
rect 22622 23366 22674 23418
rect 22686 23366 22738 23418
rect 3056 23264 3108 23316
rect 8300 23264 8352 23316
rect 10232 23264 10284 23316
rect 11060 23264 11112 23316
rect 11612 23264 11664 23316
rect 11796 23307 11848 23316
rect 11796 23273 11805 23307
rect 11805 23273 11839 23307
rect 11839 23273 11848 23307
rect 11796 23264 11848 23273
rect 2228 23171 2280 23180
rect 2228 23137 2237 23171
rect 2237 23137 2271 23171
rect 2271 23137 2280 23171
rect 2228 23128 2280 23137
rect 2412 23171 2464 23180
rect 2412 23137 2421 23171
rect 2421 23137 2455 23171
rect 2455 23137 2464 23171
rect 2412 23128 2464 23137
rect 3240 23171 3292 23180
rect 3240 23137 3249 23171
rect 3249 23137 3283 23171
rect 3283 23137 3292 23171
rect 3240 23128 3292 23137
rect 3332 23128 3384 23180
rect 5448 23128 5500 23180
rect 5724 23128 5776 23180
rect 5540 23060 5592 23112
rect 9404 23196 9456 23248
rect 15844 23264 15896 23316
rect 6736 23171 6788 23180
rect 6736 23137 6770 23171
rect 6770 23137 6788 23171
rect 6736 23128 6788 23137
rect 8208 23128 8260 23180
rect 9220 23128 9272 23180
rect 10048 23128 10100 23180
rect 10784 23171 10836 23180
rect 10784 23137 10793 23171
rect 10793 23137 10827 23171
rect 10827 23137 10836 23171
rect 10784 23128 10836 23137
rect 10968 23171 11020 23180
rect 10968 23137 10977 23171
rect 10977 23137 11011 23171
rect 11011 23137 11020 23171
rect 10968 23128 11020 23137
rect 11244 23171 11296 23180
rect 11244 23137 11253 23171
rect 11253 23137 11287 23171
rect 11287 23137 11296 23171
rect 11244 23128 11296 23137
rect 11336 23128 11388 23180
rect 11796 23128 11848 23180
rect 18236 23196 18288 23248
rect 18788 23196 18840 23248
rect 20076 23307 20128 23316
rect 20076 23273 20085 23307
rect 20085 23273 20119 23307
rect 20119 23273 20128 23307
rect 20076 23264 20128 23273
rect 21548 23196 21600 23248
rect 6368 23060 6420 23112
rect 14832 23128 14884 23180
rect 15660 23171 15712 23180
rect 15660 23137 15678 23171
rect 15678 23137 15712 23171
rect 15660 23128 15712 23137
rect 16212 23128 16264 23180
rect 20260 23171 20312 23180
rect 20260 23137 20269 23171
rect 20269 23137 20303 23171
rect 20303 23137 20312 23171
rect 20260 23128 20312 23137
rect 23388 23128 23440 23180
rect 5080 22992 5132 23044
rect 10140 22992 10192 23044
rect 13820 23103 13872 23112
rect 13820 23069 13829 23103
rect 13829 23069 13863 23103
rect 13863 23069 13872 23103
rect 13820 23060 13872 23069
rect 15936 23103 15988 23112
rect 15936 23069 15945 23103
rect 15945 23069 15979 23103
rect 15979 23069 15988 23103
rect 15936 23060 15988 23069
rect 18696 23103 18748 23112
rect 18696 23069 18705 23103
rect 18705 23069 18739 23103
rect 18739 23069 18748 23103
rect 18696 23060 18748 23069
rect 20812 23060 20864 23112
rect 22836 23060 22888 23112
rect 16028 22992 16080 23044
rect 17960 23035 18012 23044
rect 17960 23001 17969 23035
rect 17969 23001 18003 23035
rect 18003 23001 18012 23035
rect 17960 22992 18012 23001
rect 1768 22924 1820 22976
rect 3976 22924 4028 22976
rect 4896 22967 4948 22976
rect 4896 22933 4905 22967
rect 4905 22933 4939 22967
rect 4939 22933 4948 22967
rect 4896 22924 4948 22933
rect 5448 22924 5500 22976
rect 8116 22924 8168 22976
rect 8576 22967 8628 22976
rect 8576 22933 8585 22967
rect 8585 22933 8619 22967
rect 8619 22933 8628 22967
rect 8576 22924 8628 22933
rect 13176 22924 13228 22976
rect 14464 22967 14516 22976
rect 14464 22933 14473 22967
rect 14473 22933 14507 22967
rect 14507 22933 14516 22967
rect 14464 22924 14516 22933
rect 18880 22924 18932 22976
rect 21364 22924 21416 22976
rect 21640 22924 21692 22976
rect 1366 22822 1418 22874
rect 1430 22822 1482 22874
rect 1494 22822 1546 22874
rect 1558 22822 1610 22874
rect 1622 22822 1674 22874
rect 1686 22822 1738 22874
rect 7366 22822 7418 22874
rect 7430 22822 7482 22874
rect 7494 22822 7546 22874
rect 7558 22822 7610 22874
rect 7622 22822 7674 22874
rect 7686 22822 7738 22874
rect 13366 22822 13418 22874
rect 13430 22822 13482 22874
rect 13494 22822 13546 22874
rect 13558 22822 13610 22874
rect 13622 22822 13674 22874
rect 13686 22822 13738 22874
rect 19366 22822 19418 22874
rect 19430 22822 19482 22874
rect 19494 22822 19546 22874
rect 19558 22822 19610 22874
rect 19622 22822 19674 22874
rect 19686 22822 19738 22874
rect 5540 22763 5592 22772
rect 5540 22729 5549 22763
rect 5549 22729 5583 22763
rect 5583 22729 5592 22763
rect 5540 22720 5592 22729
rect 5724 22763 5776 22772
rect 5724 22729 5733 22763
rect 5733 22729 5767 22763
rect 5767 22729 5776 22763
rect 5724 22720 5776 22729
rect 6736 22720 6788 22772
rect 9220 22763 9272 22772
rect 9220 22729 9229 22763
rect 9229 22729 9263 22763
rect 9263 22729 9272 22763
rect 9220 22720 9272 22729
rect 9496 22763 9548 22772
rect 9496 22729 9505 22763
rect 9505 22729 9539 22763
rect 9539 22729 9548 22763
rect 9496 22720 9548 22729
rect 9956 22720 10008 22772
rect 4804 22652 4856 22704
rect 5632 22652 5684 22704
rect 1492 22559 1544 22568
rect 1492 22525 1501 22559
rect 1501 22525 1535 22559
rect 1535 22525 1544 22559
rect 1492 22516 1544 22525
rect 1768 22559 1820 22568
rect 1768 22525 1777 22559
rect 1777 22525 1811 22559
rect 1811 22525 1820 22559
rect 1768 22516 1820 22525
rect 2964 22627 3016 22636
rect 2964 22593 2973 22627
rect 2973 22593 3007 22627
rect 3007 22593 3016 22627
rect 2964 22584 3016 22593
rect 4252 22584 4304 22636
rect 3700 22559 3752 22568
rect 3700 22525 3709 22559
rect 3709 22525 3743 22559
rect 3743 22525 3752 22559
rect 3700 22516 3752 22525
rect 3976 22559 4028 22568
rect 3976 22525 3985 22559
rect 3985 22525 4019 22559
rect 4019 22525 4028 22559
rect 3976 22516 4028 22525
rect 4160 22559 4212 22568
rect 4160 22525 4169 22559
rect 4169 22525 4203 22559
rect 4203 22525 4212 22559
rect 4160 22516 4212 22525
rect 4896 22516 4948 22568
rect 6092 22584 6144 22636
rect 8576 22652 8628 22704
rect 11244 22720 11296 22772
rect 7840 22584 7892 22636
rect 8116 22627 8168 22636
rect 8116 22593 8125 22627
rect 8125 22593 8159 22627
rect 8159 22593 8168 22627
rect 8116 22584 8168 22593
rect 1768 22380 1820 22432
rect 5080 22448 5132 22500
rect 5540 22448 5592 22500
rect 6092 22491 6144 22500
rect 6092 22457 6101 22491
rect 6101 22457 6135 22491
rect 6135 22457 6144 22491
rect 6092 22448 6144 22457
rect 5264 22380 5316 22432
rect 5356 22423 5408 22432
rect 5356 22389 5365 22423
rect 5365 22389 5399 22423
rect 5399 22389 5408 22423
rect 5356 22380 5408 22389
rect 6184 22423 6236 22432
rect 6184 22389 6193 22423
rect 6193 22389 6227 22423
rect 6227 22389 6236 22423
rect 6184 22380 6236 22389
rect 7288 22516 7340 22568
rect 9220 22516 9272 22568
rect 9312 22559 9364 22568
rect 9312 22525 9321 22559
rect 9321 22525 9355 22559
rect 9355 22525 9364 22559
rect 9312 22516 9364 22525
rect 9680 22559 9732 22568
rect 9680 22525 9689 22559
rect 9689 22525 9723 22559
rect 9723 22525 9732 22559
rect 9680 22516 9732 22525
rect 10140 22516 10192 22568
rect 7748 22448 7800 22500
rect 11520 22559 11572 22568
rect 11520 22525 11529 22559
rect 11529 22525 11563 22559
rect 11563 22525 11572 22559
rect 11520 22516 11572 22525
rect 12624 22516 12676 22568
rect 13820 22652 13872 22704
rect 14372 22695 14424 22704
rect 14372 22661 14381 22695
rect 14381 22661 14415 22695
rect 14415 22661 14424 22695
rect 14372 22652 14424 22661
rect 15016 22652 15068 22704
rect 15476 22652 15528 22704
rect 7196 22423 7248 22432
rect 7196 22389 7205 22423
rect 7205 22389 7239 22423
rect 7239 22389 7248 22423
rect 7196 22380 7248 22389
rect 10232 22380 10284 22432
rect 11244 22380 11296 22432
rect 11980 22380 12032 22432
rect 12256 22380 12308 22432
rect 13176 22516 13228 22568
rect 13452 22516 13504 22568
rect 17132 22720 17184 22772
rect 19708 22720 19760 22772
rect 20076 22720 20128 22772
rect 14464 22516 14516 22568
rect 15200 22516 15252 22568
rect 16120 22516 16172 22568
rect 19064 22652 19116 22704
rect 17316 22584 17368 22636
rect 17960 22584 18012 22636
rect 19800 22652 19852 22704
rect 20904 22652 20956 22704
rect 13636 22448 13688 22500
rect 14556 22448 14608 22500
rect 15936 22448 15988 22500
rect 20444 22516 20496 22568
rect 14280 22380 14332 22432
rect 15108 22380 15160 22432
rect 15384 22380 15436 22432
rect 15568 22380 15620 22432
rect 17040 22423 17092 22432
rect 17040 22389 17049 22423
rect 17049 22389 17083 22423
rect 17083 22389 17092 22423
rect 17040 22380 17092 22389
rect 20260 22448 20312 22500
rect 20628 22491 20680 22500
rect 20628 22457 20637 22491
rect 20637 22457 20671 22491
rect 20671 22457 20680 22491
rect 20628 22448 20680 22457
rect 20720 22491 20772 22500
rect 20720 22457 20729 22491
rect 20729 22457 20763 22491
rect 20763 22457 20772 22491
rect 20720 22448 20772 22457
rect 21088 22516 21140 22568
rect 22192 22516 22244 22568
rect 22836 22516 22888 22568
rect 21640 22448 21692 22500
rect 23020 22448 23072 22500
rect 19340 22380 19392 22432
rect 19708 22380 19760 22432
rect 21088 22423 21140 22432
rect 21088 22389 21097 22423
rect 21097 22389 21131 22423
rect 21131 22389 21140 22423
rect 21088 22380 21140 22389
rect 4366 22278 4418 22330
rect 4430 22278 4482 22330
rect 4494 22278 4546 22330
rect 4558 22278 4610 22330
rect 4622 22278 4674 22330
rect 4686 22278 4738 22330
rect 10366 22278 10418 22330
rect 10430 22278 10482 22330
rect 10494 22278 10546 22330
rect 10558 22278 10610 22330
rect 10622 22278 10674 22330
rect 10686 22278 10738 22330
rect 16366 22278 16418 22330
rect 16430 22278 16482 22330
rect 16494 22278 16546 22330
rect 16558 22278 16610 22330
rect 16622 22278 16674 22330
rect 16686 22278 16738 22330
rect 22366 22278 22418 22330
rect 22430 22278 22482 22330
rect 22494 22278 22546 22330
rect 22558 22278 22610 22330
rect 22622 22278 22674 22330
rect 22686 22278 22738 22330
rect 1492 22176 1544 22228
rect 2412 22176 2464 22228
rect 2228 22108 2280 22160
rect 3332 22176 3384 22228
rect 4804 22219 4856 22228
rect 4804 22185 4813 22219
rect 4813 22185 4847 22219
rect 4847 22185 4856 22219
rect 4804 22176 4856 22185
rect 3516 22108 3568 22160
rect 3700 22151 3752 22160
rect 3700 22117 3709 22151
rect 3709 22117 3743 22151
rect 3743 22117 3752 22151
rect 5448 22176 5500 22228
rect 5540 22176 5592 22228
rect 3700 22108 3752 22117
rect 1860 22083 1912 22092
rect 1860 22049 1869 22083
rect 1869 22049 1903 22083
rect 1903 22049 1912 22083
rect 1860 22040 1912 22049
rect 2044 22040 2096 22092
rect 2228 21972 2280 22024
rect 2964 22083 3016 22092
rect 2964 22049 2973 22083
rect 2973 22049 3007 22083
rect 3007 22049 3016 22083
rect 2964 22040 3016 22049
rect 3424 22040 3476 22092
rect 3884 22083 3936 22092
rect 2872 21972 2924 22024
rect 3056 22015 3108 22024
rect 3056 21981 3065 22015
rect 3065 21981 3099 22015
rect 3099 21981 3108 22015
rect 3056 21972 3108 21981
rect 3884 22049 3893 22083
rect 3893 22049 3927 22083
rect 3927 22049 3936 22083
rect 3884 22040 3936 22049
rect 7196 22176 7248 22228
rect 4068 21972 4120 22024
rect 4252 21972 4304 22024
rect 4712 22040 4764 22092
rect 5172 22040 5224 22092
rect 5264 22083 5316 22092
rect 5264 22049 5273 22083
rect 5273 22049 5307 22083
rect 5307 22049 5316 22083
rect 5264 22040 5316 22049
rect 5448 22083 5500 22092
rect 5448 22049 5457 22083
rect 5457 22049 5491 22083
rect 5491 22049 5500 22083
rect 5448 22040 5500 22049
rect 6460 22108 6512 22160
rect 7748 22108 7800 22160
rect 8668 22176 8720 22228
rect 9680 22176 9732 22228
rect 5080 21904 5132 21956
rect 1952 21836 2004 21888
rect 3332 21836 3384 21888
rect 3884 21836 3936 21888
rect 4712 21836 4764 21888
rect 4896 21879 4948 21888
rect 4896 21845 4905 21879
rect 4905 21845 4939 21879
rect 4939 21845 4948 21879
rect 4896 21836 4948 21845
rect 7196 22040 7248 22092
rect 8484 22108 8536 22160
rect 9128 22108 9180 22160
rect 9404 22108 9456 22160
rect 10048 22108 10100 22160
rect 10968 22176 11020 22228
rect 6460 21972 6512 22024
rect 5816 21904 5868 21956
rect 8116 21972 8168 22024
rect 8392 22083 8444 22092
rect 8392 22049 8401 22083
rect 8401 22049 8435 22083
rect 8435 22049 8444 22083
rect 8392 22040 8444 22049
rect 7932 21904 7984 21956
rect 8024 21947 8076 21956
rect 8024 21913 8033 21947
rect 8033 21913 8067 21947
rect 8067 21913 8076 21947
rect 8024 21904 8076 21913
rect 9496 22015 9548 22024
rect 9496 21981 9505 22015
rect 9505 21981 9539 22015
rect 9539 21981 9548 22015
rect 9496 21972 9548 21981
rect 9588 22015 9640 22024
rect 9588 21981 9597 22015
rect 9597 21981 9631 22015
rect 9631 21981 9640 22015
rect 9588 21972 9640 21981
rect 9680 22015 9732 22024
rect 9680 21981 9689 22015
rect 9689 21981 9723 22015
rect 9723 21981 9732 22015
rect 9680 21972 9732 21981
rect 10324 22040 10376 22092
rect 10784 22083 10836 22092
rect 10784 22049 10793 22083
rect 10793 22049 10827 22083
rect 10827 22049 10836 22083
rect 10784 22040 10836 22049
rect 11520 22176 11572 22228
rect 15660 22176 15712 22228
rect 15844 22176 15896 22228
rect 16028 22176 16080 22228
rect 16212 22176 16264 22228
rect 17224 22176 17276 22228
rect 11244 22151 11296 22160
rect 11244 22117 11253 22151
rect 11253 22117 11287 22151
rect 11287 22117 11296 22151
rect 11244 22108 11296 22117
rect 11428 22083 11480 22092
rect 11428 22049 11437 22083
rect 11437 22049 11471 22083
rect 11471 22049 11480 22083
rect 11428 22040 11480 22049
rect 12256 22108 12308 22160
rect 13452 22108 13504 22160
rect 13636 22151 13688 22160
rect 13636 22117 13645 22151
rect 13645 22117 13679 22151
rect 13679 22117 13688 22151
rect 13636 22108 13688 22117
rect 12532 22040 12584 22092
rect 13728 22040 13780 22092
rect 14372 22108 14424 22160
rect 14832 22151 14884 22160
rect 14832 22117 14841 22151
rect 14841 22117 14875 22151
rect 14875 22117 14884 22151
rect 14832 22108 14884 22117
rect 15016 22151 15068 22160
rect 15016 22117 15025 22151
rect 15025 22117 15059 22151
rect 15059 22117 15068 22151
rect 15016 22108 15068 22117
rect 17960 22108 18012 22160
rect 20168 22176 20220 22228
rect 20260 22219 20312 22228
rect 20260 22185 20269 22219
rect 20269 22185 20303 22219
rect 20303 22185 20312 22219
rect 20260 22176 20312 22185
rect 19432 22108 19484 22160
rect 20628 22176 20680 22228
rect 20720 22108 20772 22160
rect 14188 22083 14240 22092
rect 14188 22049 14197 22083
rect 14197 22049 14231 22083
rect 14231 22049 14240 22083
rect 14188 22040 14240 22049
rect 15292 22040 15344 22092
rect 15384 22083 15436 22092
rect 15384 22049 15393 22083
rect 15393 22049 15427 22083
rect 15427 22049 15436 22083
rect 15384 22040 15436 22049
rect 15660 22083 15712 22092
rect 15660 22049 15669 22083
rect 15669 22049 15703 22083
rect 15703 22049 15712 22083
rect 15660 22040 15712 22049
rect 16120 22083 16172 22092
rect 16120 22049 16129 22083
rect 16129 22049 16163 22083
rect 16163 22049 16172 22083
rect 16120 22040 16172 22049
rect 16856 22083 16908 22092
rect 16856 22049 16865 22083
rect 16865 22049 16899 22083
rect 16899 22049 16908 22083
rect 16856 22040 16908 22049
rect 8576 21947 8628 21956
rect 8576 21913 8585 21947
rect 8585 21913 8619 21947
rect 8619 21913 8628 21947
rect 8576 21904 8628 21913
rect 9220 21947 9272 21956
rect 9220 21913 9229 21947
rect 9229 21913 9263 21947
rect 9263 21913 9272 21947
rect 9220 21904 9272 21913
rect 6184 21836 6236 21888
rect 6552 21836 6604 21888
rect 7104 21836 7156 21888
rect 8392 21836 8444 21888
rect 9036 21879 9088 21888
rect 9036 21845 9045 21879
rect 9045 21845 9079 21879
rect 9079 21845 9088 21879
rect 9036 21836 9088 21845
rect 9404 21836 9456 21888
rect 14280 22015 14332 22024
rect 14280 21981 14289 22015
rect 14289 21981 14323 22015
rect 14323 21981 14332 22015
rect 14280 21972 14332 21981
rect 17868 22040 17920 22092
rect 18604 22040 18656 22092
rect 18696 22083 18748 22092
rect 18696 22049 18705 22083
rect 18705 22049 18739 22083
rect 18739 22049 18748 22083
rect 18696 22040 18748 22049
rect 19156 22040 19208 22092
rect 17132 22015 17184 22024
rect 17132 21981 17141 22015
rect 17141 21981 17175 22015
rect 17175 21981 17184 22015
rect 17132 21972 17184 21981
rect 17316 21972 17368 22024
rect 18972 22015 19024 22024
rect 18972 21981 18981 22015
rect 18981 21981 19015 22015
rect 19015 21981 19024 22015
rect 18972 21972 19024 21981
rect 19984 22083 20036 22092
rect 19984 22049 19993 22083
rect 19993 22049 20027 22083
rect 20027 22049 20036 22083
rect 19984 22040 20036 22049
rect 20168 22083 20220 22092
rect 20168 22049 20177 22083
rect 20177 22049 20211 22083
rect 20211 22049 20220 22083
rect 20168 22040 20220 22049
rect 20260 22040 20312 22092
rect 21548 22083 21600 22092
rect 21548 22049 21582 22083
rect 21582 22049 21600 22083
rect 9864 21904 9916 21956
rect 12716 21904 12768 21956
rect 13268 21904 13320 21956
rect 20352 21972 20404 22024
rect 20536 21972 20588 22024
rect 12072 21879 12124 21888
rect 12072 21845 12081 21879
rect 12081 21845 12115 21879
rect 12115 21845 12124 21879
rect 12072 21836 12124 21845
rect 12532 21879 12584 21888
rect 12532 21845 12541 21879
rect 12541 21845 12575 21879
rect 12575 21845 12584 21879
rect 12532 21836 12584 21845
rect 12624 21836 12676 21888
rect 15016 21836 15068 21888
rect 16396 21836 16448 21888
rect 16856 21836 16908 21888
rect 19800 21904 19852 21956
rect 21548 22040 21600 22049
rect 22928 22151 22980 22160
rect 22928 22117 22937 22151
rect 22937 22117 22971 22151
rect 22971 22117 22980 22151
rect 22928 22108 22980 22117
rect 21272 22015 21324 22024
rect 21272 21981 21281 22015
rect 21281 21981 21315 22015
rect 21315 21981 21324 22015
rect 21272 21972 21324 21981
rect 19432 21836 19484 21888
rect 20812 21836 20864 21888
rect 21180 21836 21232 21888
rect 21272 21836 21324 21888
rect 22192 21836 22244 21888
rect 22284 21836 22336 21888
rect 1366 21734 1418 21786
rect 1430 21734 1482 21786
rect 1494 21734 1546 21786
rect 1558 21734 1610 21786
rect 1622 21734 1674 21786
rect 1686 21734 1738 21786
rect 7366 21734 7418 21786
rect 7430 21734 7482 21786
rect 7494 21734 7546 21786
rect 7558 21734 7610 21786
rect 7622 21734 7674 21786
rect 7686 21734 7738 21786
rect 13366 21734 13418 21786
rect 13430 21734 13482 21786
rect 13494 21734 13546 21786
rect 13558 21734 13610 21786
rect 13622 21734 13674 21786
rect 13686 21734 13738 21786
rect 19366 21734 19418 21786
rect 19430 21734 19482 21786
rect 19494 21734 19546 21786
rect 19558 21734 19610 21786
rect 19622 21734 19674 21786
rect 19686 21734 19738 21786
rect 1860 21632 1912 21684
rect 3424 21675 3476 21684
rect 3424 21641 3433 21675
rect 3433 21641 3467 21675
rect 3467 21641 3476 21675
rect 3424 21632 3476 21641
rect 5172 21632 5224 21684
rect 5908 21675 5960 21684
rect 5908 21641 5917 21675
rect 5917 21641 5951 21675
rect 5951 21641 5960 21675
rect 5908 21632 5960 21641
rect 3240 21564 3292 21616
rect 2780 21539 2832 21548
rect 2780 21505 2789 21539
rect 2789 21505 2823 21539
rect 2823 21505 2832 21539
rect 2780 21496 2832 21505
rect 2964 21539 3016 21548
rect 2964 21505 2973 21539
rect 2973 21505 3007 21539
rect 3007 21505 3016 21539
rect 5264 21564 5316 21616
rect 2964 21496 3016 21505
rect 1952 21471 2004 21480
rect 1952 21437 1970 21471
rect 1970 21437 2004 21471
rect 1952 21428 2004 21437
rect 2504 21471 2556 21480
rect 2504 21437 2513 21471
rect 2513 21437 2547 21471
rect 2547 21437 2556 21471
rect 2504 21428 2556 21437
rect 3148 21428 3200 21480
rect 2136 21360 2188 21412
rect 2872 21360 2924 21412
rect 3332 21360 3384 21412
rect 3884 21471 3936 21480
rect 3884 21437 3893 21471
rect 3893 21437 3927 21471
rect 3927 21437 3936 21471
rect 3884 21428 3936 21437
rect 4252 21428 4304 21480
rect 4896 21496 4948 21548
rect 6828 21632 6880 21684
rect 6644 21564 6696 21616
rect 7472 21675 7524 21684
rect 7472 21641 7481 21675
rect 7481 21641 7515 21675
rect 7515 21641 7524 21675
rect 7472 21632 7524 21641
rect 8852 21632 8904 21684
rect 8024 21564 8076 21616
rect 9312 21564 9364 21616
rect 2044 21292 2096 21344
rect 2596 21292 2648 21344
rect 2964 21292 3016 21344
rect 5172 21471 5224 21480
rect 5172 21437 5181 21471
rect 5181 21437 5215 21471
rect 5215 21437 5224 21471
rect 5172 21428 5224 21437
rect 5632 21428 5684 21480
rect 7932 21496 7984 21548
rect 6184 21471 6236 21480
rect 6184 21437 6193 21471
rect 6193 21437 6227 21471
rect 6227 21437 6236 21471
rect 6184 21428 6236 21437
rect 6644 21471 6696 21480
rect 6644 21437 6653 21471
rect 6653 21437 6687 21471
rect 6687 21437 6696 21471
rect 6644 21428 6696 21437
rect 6920 21471 6972 21480
rect 6920 21437 6929 21471
rect 6929 21437 6963 21471
rect 6963 21437 6972 21471
rect 6920 21428 6972 21437
rect 7012 21471 7064 21480
rect 7012 21437 7021 21471
rect 7021 21437 7055 21471
rect 7055 21437 7064 21471
rect 7012 21428 7064 21437
rect 7196 21428 7248 21480
rect 7380 21471 7432 21480
rect 7380 21437 7389 21471
rect 7389 21437 7423 21471
rect 7423 21437 7432 21471
rect 7380 21428 7432 21437
rect 7656 21471 7708 21480
rect 7656 21437 7665 21471
rect 7665 21437 7699 21471
rect 7699 21437 7708 21471
rect 7656 21428 7708 21437
rect 8392 21428 8444 21480
rect 8852 21496 8904 21548
rect 9496 21607 9548 21616
rect 9496 21573 9505 21607
rect 9505 21573 9539 21607
rect 9539 21573 9548 21607
rect 9496 21564 9548 21573
rect 10048 21632 10100 21684
rect 14188 21632 14240 21684
rect 15384 21632 15436 21684
rect 15752 21632 15804 21684
rect 19248 21632 19300 21684
rect 19524 21632 19576 21684
rect 16028 21564 16080 21616
rect 20812 21632 20864 21684
rect 20168 21564 20220 21616
rect 8944 21428 8996 21480
rect 9312 21471 9364 21480
rect 9312 21437 9321 21471
rect 9321 21437 9355 21471
rect 9355 21437 9364 21471
rect 9312 21428 9364 21437
rect 9864 21428 9916 21480
rect 10324 21428 10376 21480
rect 11980 21496 12032 21548
rect 10784 21428 10836 21480
rect 11428 21428 11480 21480
rect 11520 21428 11572 21480
rect 12624 21428 12676 21480
rect 13176 21471 13228 21480
rect 13176 21437 13185 21471
rect 13185 21437 13219 21471
rect 13219 21437 13228 21471
rect 13176 21428 13228 21437
rect 4896 21335 4948 21344
rect 4896 21301 4905 21335
rect 4905 21301 4939 21335
rect 4939 21301 4948 21335
rect 4896 21292 4948 21301
rect 5080 21335 5132 21344
rect 5080 21301 5089 21335
rect 5089 21301 5123 21335
rect 5123 21301 5132 21335
rect 5080 21292 5132 21301
rect 5816 21292 5868 21344
rect 5908 21292 5960 21344
rect 7472 21292 7524 21344
rect 8300 21292 8352 21344
rect 9680 21292 9732 21344
rect 9864 21292 9916 21344
rect 11980 21360 12032 21412
rect 10784 21292 10836 21344
rect 11428 21335 11480 21344
rect 11428 21301 11437 21335
rect 11437 21301 11471 21335
rect 11471 21301 11480 21335
rect 11428 21292 11480 21301
rect 11704 21335 11756 21344
rect 11704 21301 11713 21335
rect 11713 21301 11747 21335
rect 11747 21301 11756 21335
rect 11704 21292 11756 21301
rect 12716 21292 12768 21344
rect 12808 21335 12860 21344
rect 12808 21301 12817 21335
rect 12817 21301 12851 21335
rect 12851 21301 12860 21335
rect 12808 21292 12860 21301
rect 13912 21335 13964 21344
rect 13912 21301 13921 21335
rect 13921 21301 13955 21335
rect 13955 21301 13964 21335
rect 13912 21292 13964 21301
rect 14188 21471 14240 21480
rect 14188 21437 14197 21471
rect 14197 21437 14231 21471
rect 14231 21437 14240 21471
rect 14188 21428 14240 21437
rect 14280 21471 14332 21480
rect 14280 21437 14289 21471
rect 14289 21437 14323 21471
rect 14323 21437 14332 21471
rect 14280 21428 14332 21437
rect 14372 21471 14424 21480
rect 14372 21437 14381 21471
rect 14381 21437 14415 21471
rect 14415 21437 14424 21471
rect 14372 21428 14424 21437
rect 14464 21471 14516 21480
rect 14464 21437 14473 21471
rect 14473 21437 14507 21471
rect 14507 21437 14516 21471
rect 14464 21428 14516 21437
rect 15292 21496 15344 21548
rect 15568 21496 15620 21548
rect 14740 21428 14792 21480
rect 14096 21360 14148 21412
rect 15200 21360 15252 21412
rect 15384 21360 15436 21412
rect 15844 21360 15896 21412
rect 16672 21471 16724 21480
rect 16672 21437 16681 21471
rect 16681 21437 16715 21471
rect 16715 21437 16724 21471
rect 16672 21428 16724 21437
rect 19064 21496 19116 21548
rect 19248 21496 19300 21548
rect 19892 21428 19944 21480
rect 20076 21471 20128 21480
rect 20076 21437 20085 21471
rect 20085 21437 20119 21471
rect 20119 21437 20128 21471
rect 20076 21428 20128 21437
rect 20168 21471 20220 21480
rect 20168 21437 20177 21471
rect 20177 21437 20211 21471
rect 20211 21437 20220 21471
rect 20168 21428 20220 21437
rect 21088 21564 21140 21616
rect 21456 21564 21508 21616
rect 16120 21292 16172 21344
rect 16396 21292 16448 21344
rect 17776 21360 17828 21412
rect 19248 21360 19300 21412
rect 19524 21360 19576 21412
rect 19708 21360 19760 21412
rect 16948 21292 17000 21344
rect 17500 21292 17552 21344
rect 18420 21335 18472 21344
rect 18420 21301 18429 21335
rect 18429 21301 18463 21335
rect 18463 21301 18472 21335
rect 18420 21292 18472 21301
rect 18880 21335 18932 21344
rect 18880 21301 18889 21335
rect 18889 21301 18923 21335
rect 18923 21301 18932 21335
rect 18880 21292 18932 21301
rect 19432 21335 19484 21344
rect 19432 21301 19441 21335
rect 19441 21301 19475 21335
rect 19475 21301 19484 21335
rect 19432 21292 19484 21301
rect 19984 21360 20036 21412
rect 20536 21428 20588 21480
rect 22836 21496 22888 21548
rect 21364 21428 21416 21480
rect 20812 21403 20864 21412
rect 20812 21369 20821 21403
rect 20821 21369 20855 21403
rect 20855 21369 20864 21403
rect 20812 21360 20864 21369
rect 22008 21360 22060 21412
rect 22284 21360 22336 21412
rect 21456 21292 21508 21344
rect 4366 21190 4418 21242
rect 4430 21190 4482 21242
rect 4494 21190 4546 21242
rect 4558 21190 4610 21242
rect 4622 21190 4674 21242
rect 4686 21190 4738 21242
rect 10366 21190 10418 21242
rect 10430 21190 10482 21242
rect 10494 21190 10546 21242
rect 10558 21190 10610 21242
rect 10622 21190 10674 21242
rect 10686 21190 10738 21242
rect 16366 21190 16418 21242
rect 16430 21190 16482 21242
rect 16494 21190 16546 21242
rect 16558 21190 16610 21242
rect 16622 21190 16674 21242
rect 16686 21190 16738 21242
rect 22366 21190 22418 21242
rect 22430 21190 22482 21242
rect 22494 21190 22546 21242
rect 22558 21190 22610 21242
rect 22622 21190 22674 21242
rect 22686 21190 22738 21242
rect 2228 21088 2280 21140
rect 1860 20995 1912 21004
rect 1860 20961 1869 20995
rect 1869 20961 1903 20995
rect 1903 20961 1912 20995
rect 1860 20952 1912 20961
rect 2136 21063 2188 21072
rect 2136 21029 2145 21063
rect 2145 21029 2179 21063
rect 2179 21029 2188 21063
rect 2136 21020 2188 21029
rect 2504 21131 2556 21140
rect 2504 21097 2513 21131
rect 2513 21097 2547 21131
rect 2547 21097 2556 21131
rect 2504 21088 2556 21097
rect 2780 21088 2832 21140
rect 5632 21131 5684 21140
rect 5632 21097 5641 21131
rect 5641 21097 5675 21131
rect 5675 21097 5684 21131
rect 5632 21088 5684 21097
rect 6276 21131 6328 21140
rect 6276 21097 6285 21131
rect 6285 21097 6319 21131
rect 6319 21097 6328 21131
rect 6276 21088 6328 21097
rect 6920 21088 6972 21140
rect 7840 21131 7892 21140
rect 7840 21097 7849 21131
rect 7849 21097 7883 21131
rect 7883 21097 7892 21131
rect 7840 21088 7892 21097
rect 9588 21088 9640 21140
rect 9772 21088 9824 21140
rect 2964 21063 3016 21072
rect 2228 20952 2280 21004
rect 2964 21029 2973 21063
rect 2973 21029 3007 21063
rect 3007 21029 3016 21063
rect 2964 21020 3016 21029
rect 3516 20952 3568 21004
rect 4344 21020 4396 21072
rect 4896 21020 4948 21072
rect 4160 20884 4212 20936
rect 3148 20859 3200 20868
rect 3148 20825 3157 20859
rect 3157 20825 3191 20859
rect 3191 20825 3200 20859
rect 3148 20816 3200 20825
rect 4620 20995 4672 21004
rect 4620 20961 4629 20995
rect 4629 20961 4663 20995
rect 4663 20961 4672 20995
rect 4620 20952 4672 20961
rect 4712 20995 4764 21004
rect 4712 20961 4721 20995
rect 4721 20961 4755 20995
rect 4755 20961 4764 20995
rect 4712 20952 4764 20961
rect 4804 20884 4856 20936
rect 4988 20995 5040 21004
rect 4988 20961 4997 20995
rect 4997 20961 5031 20995
rect 5031 20961 5040 20995
rect 4988 20952 5040 20961
rect 5264 20995 5316 21004
rect 5264 20961 5273 20995
rect 5273 20961 5307 20995
rect 5307 20961 5316 20995
rect 5264 20952 5316 20961
rect 5540 20952 5592 21004
rect 5816 20995 5868 21004
rect 5816 20961 5825 20995
rect 5825 20961 5859 20995
rect 5859 20961 5868 20995
rect 5816 20952 5868 20961
rect 6092 20995 6144 21004
rect 6092 20961 6101 20995
rect 6101 20961 6135 20995
rect 6135 20961 6144 20995
rect 6092 20952 6144 20961
rect 6460 20995 6512 21004
rect 6460 20961 6469 20995
rect 6469 20961 6503 20995
rect 6503 20961 6512 20995
rect 6460 20952 6512 20961
rect 7104 20952 7156 21004
rect 7840 20952 7892 21004
rect 7932 20995 7984 21004
rect 7932 20961 7941 20995
rect 7941 20961 7975 20995
rect 7975 20961 7984 20995
rect 7932 20952 7984 20961
rect 8116 20995 8168 21004
rect 8116 20961 8125 20995
rect 8125 20961 8159 20995
rect 8159 20961 8168 20995
rect 8116 20952 8168 20961
rect 4988 20816 5040 20868
rect 7012 20884 7064 20936
rect 7288 20884 7340 20936
rect 8668 20927 8720 20936
rect 8668 20893 8677 20927
rect 8677 20893 8711 20927
rect 8711 20893 8720 20927
rect 8668 20884 8720 20893
rect 9680 21020 9732 21072
rect 9864 20995 9916 21004
rect 9864 20961 9873 20995
rect 9873 20961 9907 20995
rect 9907 20961 9916 20995
rect 9864 20952 9916 20961
rect 9588 20884 9640 20936
rect 9772 20927 9824 20936
rect 9772 20893 9781 20927
rect 9781 20893 9815 20927
rect 9815 20893 9824 20927
rect 9772 20884 9824 20893
rect 10784 21020 10836 21072
rect 10048 20952 10100 21004
rect 10692 20952 10744 21004
rect 11244 20995 11296 21004
rect 11244 20961 11253 20995
rect 11253 20961 11287 20995
rect 11287 20961 11296 20995
rect 11244 20952 11296 20961
rect 11704 21088 11756 21140
rect 12164 21131 12216 21140
rect 12164 21097 12173 21131
rect 12173 21097 12207 21131
rect 12207 21097 12216 21131
rect 12164 21088 12216 21097
rect 11796 21020 11848 21072
rect 11980 20995 12032 21004
rect 11980 20961 11989 20995
rect 11989 20961 12023 20995
rect 12023 20961 12032 20995
rect 11980 20952 12032 20961
rect 12072 20995 12124 21004
rect 12072 20961 12081 20995
rect 12081 20961 12115 20995
rect 12115 20961 12124 20995
rect 12072 20952 12124 20961
rect 13268 20995 13320 21004
rect 14096 21020 14148 21072
rect 15384 21088 15436 21140
rect 13268 20961 13286 20995
rect 13286 20961 13320 20995
rect 13268 20952 13320 20961
rect 13820 20995 13872 21004
rect 13820 20961 13829 20995
rect 13829 20961 13863 20995
rect 13863 20961 13872 20995
rect 13820 20952 13872 20961
rect 14740 21020 14792 21072
rect 15752 21088 15804 21140
rect 19064 21088 19116 21140
rect 19984 21088 20036 21140
rect 14832 20995 14884 21004
rect 14832 20961 14841 20995
rect 14841 20961 14875 20995
rect 14875 20961 14884 20995
rect 14832 20952 14884 20961
rect 17592 21020 17644 21072
rect 18604 21020 18656 21072
rect 20076 21020 20128 21072
rect 20444 21088 20496 21140
rect 20812 21063 20864 21072
rect 20812 21029 20821 21063
rect 20821 21029 20855 21063
rect 20855 21029 20864 21063
rect 20812 21020 20864 21029
rect 20904 21063 20956 21072
rect 20904 21029 20913 21063
rect 20913 21029 20947 21063
rect 20947 21029 20956 21063
rect 20904 21020 20956 21029
rect 20996 21020 21048 21072
rect 16396 20995 16448 21004
rect 16396 20961 16430 20995
rect 16430 20961 16448 20995
rect 16396 20952 16448 20961
rect 16764 20952 16816 21004
rect 20720 20995 20772 21004
rect 20720 20961 20729 20995
rect 20729 20961 20763 20995
rect 20763 20961 20772 20995
rect 20720 20952 20772 20961
rect 21088 20995 21140 21004
rect 21088 20961 21097 20995
rect 21097 20961 21131 20995
rect 21131 20961 21140 20995
rect 21088 20952 21140 20961
rect 22744 20995 22796 21004
rect 22744 20961 22762 20995
rect 22762 20961 22796 20995
rect 22744 20952 22796 20961
rect 22928 20952 22980 21004
rect 10324 20884 10376 20936
rect 11060 20884 11112 20936
rect 8392 20816 8444 20868
rect 4068 20791 4120 20800
rect 4068 20757 4077 20791
rect 4077 20757 4111 20791
rect 4111 20757 4120 20791
rect 4068 20748 4120 20757
rect 6184 20748 6236 20800
rect 6828 20791 6880 20800
rect 6828 20757 6837 20791
rect 6837 20757 6871 20791
rect 6871 20757 6880 20791
rect 6828 20748 6880 20757
rect 7104 20748 7156 20800
rect 7656 20748 7708 20800
rect 9496 20791 9548 20800
rect 9496 20757 9505 20791
rect 9505 20757 9539 20791
rect 9539 20757 9548 20791
rect 9496 20748 9548 20757
rect 12072 20816 12124 20868
rect 14188 20927 14240 20936
rect 14188 20893 14197 20927
rect 14197 20893 14231 20927
rect 14231 20893 14240 20927
rect 14188 20884 14240 20893
rect 15200 20884 15252 20936
rect 17592 20927 17644 20936
rect 17592 20893 17601 20927
rect 17601 20893 17635 20927
rect 17635 20893 17644 20927
rect 17592 20884 17644 20893
rect 17868 20927 17920 20936
rect 17868 20893 17877 20927
rect 17877 20893 17911 20927
rect 17911 20893 17920 20927
rect 17868 20884 17920 20893
rect 21272 20884 21324 20936
rect 21640 20884 21692 20936
rect 14096 20816 14148 20868
rect 12164 20748 12216 20800
rect 12532 20748 12584 20800
rect 14372 20748 14424 20800
rect 15292 20791 15344 20800
rect 15292 20757 15301 20791
rect 15301 20757 15335 20791
rect 15335 20757 15344 20791
rect 15292 20748 15344 20757
rect 17500 20859 17552 20868
rect 17500 20825 17509 20859
rect 17509 20825 17543 20859
rect 17543 20825 17552 20859
rect 17500 20816 17552 20825
rect 18696 20816 18748 20868
rect 20168 20816 20220 20868
rect 21088 20816 21140 20868
rect 20352 20748 20404 20800
rect 22100 20748 22152 20800
rect 22376 20748 22428 20800
rect 1366 20646 1418 20698
rect 1430 20646 1482 20698
rect 1494 20646 1546 20698
rect 1558 20646 1610 20698
rect 1622 20646 1674 20698
rect 1686 20646 1738 20698
rect 7366 20646 7418 20698
rect 7430 20646 7482 20698
rect 7494 20646 7546 20698
rect 7558 20646 7610 20698
rect 7622 20646 7674 20698
rect 7686 20646 7738 20698
rect 13366 20646 13418 20698
rect 13430 20646 13482 20698
rect 13494 20646 13546 20698
rect 13558 20646 13610 20698
rect 13622 20646 13674 20698
rect 13686 20646 13738 20698
rect 19366 20646 19418 20698
rect 19430 20646 19482 20698
rect 19494 20646 19546 20698
rect 19558 20646 19610 20698
rect 19622 20646 19674 20698
rect 19686 20646 19738 20698
rect 1860 20544 1912 20596
rect 2688 20544 2740 20596
rect 6368 20587 6420 20596
rect 6368 20553 6377 20587
rect 6377 20553 6411 20587
rect 6411 20553 6420 20587
rect 6368 20544 6420 20553
rect 6644 20544 6696 20596
rect 7196 20587 7248 20596
rect 7196 20553 7205 20587
rect 7205 20553 7239 20587
rect 7239 20553 7248 20587
rect 7196 20544 7248 20553
rect 7932 20587 7984 20596
rect 7932 20553 7941 20587
rect 7941 20553 7975 20587
rect 7975 20553 7984 20587
rect 7932 20544 7984 20553
rect 8576 20544 8628 20596
rect 9772 20544 9824 20596
rect 10232 20544 10284 20596
rect 10692 20544 10744 20596
rect 11428 20587 11480 20596
rect 11428 20553 11437 20587
rect 11437 20553 11471 20587
rect 11471 20553 11480 20587
rect 11428 20544 11480 20553
rect 12808 20544 12860 20596
rect 5540 20476 5592 20528
rect 6920 20476 6972 20528
rect 3240 20451 3292 20460
rect 3240 20417 3249 20451
rect 3249 20417 3283 20451
rect 3283 20417 3292 20451
rect 3240 20408 3292 20417
rect 4620 20408 4672 20460
rect 4896 20408 4948 20460
rect 1860 20383 1912 20392
rect 1860 20349 1869 20383
rect 1869 20349 1903 20383
rect 1903 20349 1912 20383
rect 1860 20340 1912 20349
rect 2044 20383 2096 20392
rect 2044 20349 2053 20383
rect 2053 20349 2087 20383
rect 2087 20349 2096 20383
rect 2044 20340 2096 20349
rect 2504 20383 2556 20392
rect 2504 20349 2513 20383
rect 2513 20349 2547 20383
rect 2547 20349 2556 20383
rect 2504 20340 2556 20349
rect 2780 20340 2832 20392
rect 4068 20340 4120 20392
rect 6920 20383 6972 20392
rect 6920 20349 6929 20383
rect 6929 20349 6963 20383
rect 6963 20349 6972 20383
rect 6920 20340 6972 20349
rect 7380 20383 7432 20392
rect 7380 20349 7389 20383
rect 7389 20349 7423 20383
rect 7423 20349 7432 20383
rect 7380 20340 7432 20349
rect 2596 20272 2648 20324
rect 5540 20272 5592 20324
rect 6184 20272 6236 20324
rect 1400 20247 1452 20256
rect 1400 20213 1409 20247
rect 1409 20213 1443 20247
rect 1443 20213 1452 20247
rect 1400 20204 1452 20213
rect 2044 20204 2096 20256
rect 2688 20247 2740 20256
rect 2688 20213 2697 20247
rect 2697 20213 2731 20247
rect 2731 20213 2740 20247
rect 2688 20204 2740 20213
rect 4344 20204 4396 20256
rect 5356 20204 5408 20256
rect 7012 20204 7064 20256
rect 7656 20204 7708 20256
rect 8024 20383 8076 20392
rect 8024 20349 8033 20383
rect 8033 20349 8067 20383
rect 8067 20349 8076 20383
rect 8024 20340 8076 20349
rect 8116 20272 8168 20324
rect 8392 20340 8444 20392
rect 8576 20383 8628 20392
rect 8576 20349 8585 20383
rect 8585 20349 8619 20383
rect 8619 20349 8628 20383
rect 8576 20340 8628 20349
rect 8760 20383 8812 20392
rect 8760 20349 8769 20383
rect 8769 20349 8803 20383
rect 8803 20349 8812 20383
rect 8760 20340 8812 20349
rect 9496 20340 9548 20392
rect 9864 20340 9916 20392
rect 9956 20383 10008 20392
rect 9956 20349 9965 20383
rect 9965 20349 9999 20383
rect 9999 20349 10008 20383
rect 9956 20340 10008 20349
rect 10324 20383 10376 20392
rect 10324 20349 10333 20383
rect 10333 20349 10367 20383
rect 10367 20349 10376 20383
rect 10324 20340 10376 20349
rect 10416 20383 10468 20392
rect 10416 20349 10425 20383
rect 10425 20349 10459 20383
rect 10459 20349 10468 20383
rect 10416 20340 10468 20349
rect 11520 20476 11572 20528
rect 11796 20451 11848 20460
rect 11796 20417 11805 20451
rect 11805 20417 11839 20451
rect 11839 20417 11848 20451
rect 11796 20408 11848 20417
rect 13268 20544 13320 20596
rect 14464 20544 14516 20596
rect 14556 20587 14608 20596
rect 14556 20553 14565 20587
rect 14565 20553 14599 20587
rect 14599 20553 14608 20587
rect 14556 20544 14608 20553
rect 14832 20544 14884 20596
rect 15660 20544 15712 20596
rect 16396 20544 16448 20596
rect 17316 20544 17368 20596
rect 17868 20544 17920 20596
rect 18144 20544 18196 20596
rect 22284 20544 22336 20596
rect 13820 20408 13872 20460
rect 11244 20340 11296 20392
rect 11520 20340 11572 20392
rect 8484 20204 8536 20256
rect 12072 20315 12124 20324
rect 9772 20247 9824 20256
rect 9772 20213 9781 20247
rect 9781 20213 9815 20247
rect 9815 20213 9824 20247
rect 9772 20204 9824 20213
rect 12072 20281 12106 20315
rect 12106 20281 12124 20315
rect 12072 20272 12124 20281
rect 14096 20383 14148 20392
rect 14096 20349 14105 20383
rect 14105 20349 14139 20383
rect 14139 20349 14148 20383
rect 14096 20340 14148 20349
rect 14924 20408 14976 20460
rect 16212 20451 16264 20460
rect 16212 20417 16221 20451
rect 16221 20417 16255 20451
rect 16255 20417 16264 20451
rect 16212 20408 16264 20417
rect 11060 20204 11112 20256
rect 11428 20247 11480 20256
rect 11428 20213 11437 20247
rect 11437 20213 11471 20247
rect 11471 20213 11480 20247
rect 11428 20204 11480 20213
rect 14280 20272 14332 20324
rect 14740 20340 14792 20392
rect 15292 20383 15344 20392
rect 15292 20349 15301 20383
rect 15301 20349 15335 20383
rect 15335 20349 15344 20383
rect 15292 20340 15344 20349
rect 15660 20340 15712 20392
rect 15752 20340 15804 20392
rect 16856 20476 16908 20528
rect 17224 20476 17276 20528
rect 16948 20451 17000 20460
rect 16948 20417 16957 20451
rect 16957 20417 16991 20451
rect 16991 20417 17000 20451
rect 16948 20408 17000 20417
rect 20720 20476 20772 20528
rect 20812 20519 20864 20528
rect 20812 20485 20821 20519
rect 20821 20485 20855 20519
rect 20855 20485 20864 20519
rect 20812 20476 20864 20485
rect 21824 20476 21876 20528
rect 22100 20476 22152 20528
rect 16856 20383 16908 20392
rect 16856 20349 16865 20383
rect 16865 20349 16899 20383
rect 16899 20349 16908 20383
rect 16856 20340 16908 20349
rect 17040 20272 17092 20324
rect 12624 20204 12676 20256
rect 15292 20204 15344 20256
rect 15568 20204 15620 20256
rect 18512 20383 18564 20392
rect 18512 20349 18521 20383
rect 18521 20349 18555 20383
rect 18555 20349 18564 20383
rect 18512 20340 18564 20349
rect 21180 20408 21232 20460
rect 18696 20315 18748 20324
rect 18696 20281 18705 20315
rect 18705 20281 18739 20315
rect 18739 20281 18748 20315
rect 18696 20272 18748 20281
rect 18880 20315 18932 20324
rect 18880 20281 18889 20315
rect 18889 20281 18923 20315
rect 18923 20281 18932 20315
rect 18880 20272 18932 20281
rect 17960 20204 18012 20256
rect 19340 20204 19392 20256
rect 19524 20247 19576 20256
rect 19524 20213 19533 20247
rect 19533 20213 19567 20247
rect 19567 20213 19576 20247
rect 19524 20204 19576 20213
rect 19892 20247 19944 20256
rect 19892 20213 19901 20247
rect 19901 20213 19935 20247
rect 19935 20213 19944 20247
rect 19892 20204 19944 20213
rect 20904 20340 20956 20392
rect 20996 20383 21048 20392
rect 20996 20349 21005 20383
rect 21005 20349 21039 20383
rect 21039 20349 21048 20383
rect 20996 20340 21048 20349
rect 21272 20340 21324 20392
rect 21364 20383 21416 20392
rect 21364 20349 21373 20383
rect 21373 20349 21407 20383
rect 21407 20349 21416 20383
rect 21364 20340 21416 20349
rect 21548 20340 21600 20392
rect 21824 20340 21876 20392
rect 22560 20408 22612 20460
rect 20444 20315 20496 20324
rect 20444 20281 20453 20315
rect 20453 20281 20487 20315
rect 20487 20281 20496 20315
rect 20444 20272 20496 20281
rect 20536 20315 20588 20324
rect 20536 20281 20545 20315
rect 20545 20281 20579 20315
rect 20579 20281 20588 20315
rect 20536 20272 20588 20281
rect 21456 20272 21508 20324
rect 22376 20383 22428 20392
rect 22376 20349 22385 20383
rect 22385 20349 22419 20383
rect 22419 20349 22428 20383
rect 22376 20340 22428 20349
rect 23480 20340 23532 20392
rect 22560 20272 22612 20324
rect 23296 20272 23348 20324
rect 20720 20204 20772 20256
rect 21916 20204 21968 20256
rect 23020 20204 23072 20256
rect 4366 20102 4418 20154
rect 4430 20102 4482 20154
rect 4494 20102 4546 20154
rect 4558 20102 4610 20154
rect 4622 20102 4674 20154
rect 4686 20102 4738 20154
rect 10366 20102 10418 20154
rect 10430 20102 10482 20154
rect 10494 20102 10546 20154
rect 10558 20102 10610 20154
rect 10622 20102 10674 20154
rect 10686 20102 10738 20154
rect 16366 20102 16418 20154
rect 16430 20102 16482 20154
rect 16494 20102 16546 20154
rect 16558 20102 16610 20154
rect 16622 20102 16674 20154
rect 16686 20102 16738 20154
rect 22366 20102 22418 20154
rect 22430 20102 22482 20154
rect 22494 20102 22546 20154
rect 22558 20102 22610 20154
rect 22622 20102 22674 20154
rect 22686 20102 22738 20154
rect 1952 20000 2004 20052
rect 2688 20000 2740 20052
rect 4804 20000 4856 20052
rect 5264 20000 5316 20052
rect 5816 20043 5868 20052
rect 5816 20009 5825 20043
rect 5825 20009 5859 20043
rect 5859 20009 5868 20043
rect 5816 20000 5868 20009
rect 6184 20043 6236 20052
rect 6184 20009 6193 20043
rect 6193 20009 6227 20043
rect 6227 20009 6236 20043
rect 6184 20000 6236 20009
rect 7932 20000 7984 20052
rect 2504 19975 2556 19984
rect 2504 19941 2513 19975
rect 2513 19941 2547 19975
rect 2547 19941 2556 19975
rect 2504 19932 2556 19941
rect 2964 19932 3016 19984
rect 4252 19932 4304 19984
rect 5356 19932 5408 19984
rect 1400 19864 1452 19916
rect 2044 19907 2096 19916
rect 2044 19873 2053 19907
rect 2053 19873 2087 19907
rect 2087 19873 2096 19907
rect 2044 19864 2096 19873
rect 2780 19864 2832 19916
rect 3240 19864 3292 19916
rect 3424 19907 3476 19916
rect 3424 19873 3458 19907
rect 3458 19873 3476 19907
rect 3424 19864 3476 19873
rect 5080 19864 5132 19916
rect 5448 19907 5500 19916
rect 5448 19873 5457 19907
rect 5457 19873 5491 19907
rect 5491 19873 5500 19907
rect 5448 19864 5500 19873
rect 6184 19864 6236 19916
rect 1768 19796 1820 19848
rect 4988 19796 5040 19848
rect 1860 19660 1912 19712
rect 3516 19660 3568 19712
rect 4528 19703 4580 19712
rect 4528 19669 4537 19703
rect 4537 19669 4571 19703
rect 4571 19669 4580 19703
rect 4528 19660 4580 19669
rect 5908 19796 5960 19848
rect 7288 19864 7340 19916
rect 7656 19864 7708 19916
rect 7932 19907 7984 19916
rect 7932 19873 7941 19907
rect 7941 19873 7975 19907
rect 7975 19873 7984 19907
rect 7932 19864 7984 19873
rect 8208 19864 8260 19916
rect 9772 20000 9824 20052
rect 10140 20000 10192 20052
rect 10416 20000 10468 20052
rect 8852 19932 8904 19984
rect 10876 19932 10928 19984
rect 11428 20043 11480 20052
rect 11428 20009 11437 20043
rect 11437 20009 11471 20043
rect 11471 20009 11480 20043
rect 11428 20000 11480 20009
rect 11520 20043 11572 20052
rect 11520 20009 11529 20043
rect 11529 20009 11563 20043
rect 11563 20009 11572 20043
rect 11520 20000 11572 20009
rect 11796 20000 11848 20052
rect 8484 19796 8536 19848
rect 8852 19796 8904 19848
rect 9864 19864 9916 19916
rect 10968 19907 11020 19916
rect 10968 19873 10977 19907
rect 10977 19873 11011 19907
rect 11011 19873 11020 19907
rect 10968 19864 11020 19873
rect 13084 20000 13136 20052
rect 14372 20000 14424 20052
rect 15936 20043 15988 20052
rect 15936 20009 15945 20043
rect 15945 20009 15979 20043
rect 15979 20009 15988 20043
rect 15936 20000 15988 20009
rect 16028 20000 16080 20052
rect 9772 19796 9824 19848
rect 12072 19864 12124 19916
rect 11888 19796 11940 19848
rect 12532 19907 12584 19916
rect 12532 19873 12566 19907
rect 12566 19873 12584 19907
rect 12532 19864 12584 19873
rect 14740 19932 14792 19984
rect 16948 20000 17000 20052
rect 17592 20000 17644 20052
rect 19524 20000 19576 20052
rect 20352 20000 20404 20052
rect 20444 20000 20496 20052
rect 21272 20000 21324 20052
rect 21364 20000 21416 20052
rect 13820 19864 13872 19916
rect 15108 19864 15160 19916
rect 15568 19864 15620 19916
rect 14832 19796 14884 19848
rect 15844 19864 15896 19916
rect 17040 19932 17092 19984
rect 18696 19932 18748 19984
rect 16764 19864 16816 19916
rect 20168 19864 20220 19916
rect 23388 19932 23440 19984
rect 20628 19907 20680 19916
rect 20628 19873 20637 19907
rect 20637 19873 20671 19907
rect 20671 19873 20680 19907
rect 20628 19864 20680 19873
rect 20812 19864 20864 19916
rect 21088 19907 21140 19916
rect 21088 19873 21097 19907
rect 21097 19873 21131 19907
rect 21131 19873 21140 19907
rect 21088 19864 21140 19873
rect 21364 19864 21416 19916
rect 21640 19907 21692 19916
rect 21640 19873 21649 19907
rect 21649 19873 21683 19907
rect 21683 19873 21692 19907
rect 21640 19864 21692 19873
rect 21732 19864 21784 19916
rect 7748 19728 7800 19780
rect 9036 19728 9088 19780
rect 9404 19728 9456 19780
rect 6736 19660 6788 19712
rect 7104 19703 7156 19712
rect 7104 19669 7113 19703
rect 7113 19669 7147 19703
rect 7147 19669 7156 19703
rect 7104 19660 7156 19669
rect 7196 19703 7248 19712
rect 7196 19669 7205 19703
rect 7205 19669 7239 19703
rect 7239 19669 7248 19703
rect 7196 19660 7248 19669
rect 8484 19703 8536 19712
rect 8484 19669 8493 19703
rect 8493 19669 8527 19703
rect 8527 19669 8536 19703
rect 8484 19660 8536 19669
rect 8944 19660 8996 19712
rect 9680 19660 9732 19712
rect 10416 19660 10468 19712
rect 12072 19703 12124 19712
rect 12072 19669 12081 19703
rect 12081 19669 12115 19703
rect 12115 19669 12124 19703
rect 12072 19660 12124 19669
rect 14924 19728 14976 19780
rect 16120 19728 16172 19780
rect 14740 19660 14792 19712
rect 15108 19703 15160 19712
rect 15108 19669 15117 19703
rect 15117 19669 15151 19703
rect 15151 19669 15160 19703
rect 15108 19660 15160 19669
rect 15568 19660 15620 19712
rect 16212 19660 16264 19712
rect 16304 19703 16356 19712
rect 16304 19669 16313 19703
rect 16313 19669 16347 19703
rect 16347 19669 16356 19703
rect 16304 19660 16356 19669
rect 16580 19703 16632 19712
rect 16580 19669 16589 19703
rect 16589 19669 16623 19703
rect 16623 19669 16632 19703
rect 16580 19660 16632 19669
rect 17592 19660 17644 19712
rect 18144 19703 18196 19712
rect 18144 19669 18153 19703
rect 18153 19669 18187 19703
rect 18187 19669 18196 19703
rect 18144 19660 18196 19669
rect 18696 19728 18748 19780
rect 18972 19839 19024 19848
rect 18972 19805 18981 19839
rect 18981 19805 19015 19839
rect 19015 19805 19024 19839
rect 18972 19796 19024 19805
rect 19064 19839 19116 19848
rect 19064 19805 19073 19839
rect 19073 19805 19107 19839
rect 19107 19805 19116 19839
rect 19064 19796 19116 19805
rect 19156 19796 19208 19848
rect 19800 19796 19852 19848
rect 20536 19839 20588 19848
rect 20536 19805 20545 19839
rect 20545 19805 20579 19839
rect 20579 19805 20588 19839
rect 20536 19796 20588 19805
rect 21180 19796 21232 19848
rect 20260 19728 20312 19780
rect 20812 19771 20864 19780
rect 20812 19737 20821 19771
rect 20821 19737 20855 19771
rect 20855 19737 20864 19771
rect 20812 19728 20864 19737
rect 20536 19660 20588 19712
rect 1366 19558 1418 19610
rect 1430 19558 1482 19610
rect 1494 19558 1546 19610
rect 1558 19558 1610 19610
rect 1622 19558 1674 19610
rect 1686 19558 1738 19610
rect 7366 19558 7418 19610
rect 7430 19558 7482 19610
rect 7494 19558 7546 19610
rect 7558 19558 7610 19610
rect 7622 19558 7674 19610
rect 7686 19558 7738 19610
rect 13366 19558 13418 19610
rect 13430 19558 13482 19610
rect 13494 19558 13546 19610
rect 13558 19558 13610 19610
rect 13622 19558 13674 19610
rect 13686 19558 13738 19610
rect 19366 19558 19418 19610
rect 19430 19558 19482 19610
rect 19494 19558 19546 19610
rect 19558 19558 19610 19610
rect 19622 19558 19674 19610
rect 19686 19558 19738 19610
rect 3332 19456 3384 19508
rect 3424 19456 3476 19508
rect 4988 19456 5040 19508
rect 2504 19431 2556 19440
rect 2504 19397 2513 19431
rect 2513 19397 2547 19431
rect 2547 19397 2556 19431
rect 2504 19388 2556 19397
rect 572 19320 624 19372
rect 5264 19388 5316 19440
rect 1768 19252 1820 19304
rect 1860 19295 1912 19304
rect 1860 19261 1869 19295
rect 1869 19261 1903 19295
rect 1903 19261 1912 19295
rect 1860 19252 1912 19261
rect 2228 19295 2280 19304
rect 2228 19261 2237 19295
rect 2237 19261 2271 19295
rect 2271 19261 2280 19295
rect 2228 19252 2280 19261
rect 2412 19295 2464 19304
rect 2412 19261 2421 19295
rect 2421 19261 2455 19295
rect 2455 19261 2464 19295
rect 2412 19252 2464 19261
rect 3424 19295 3476 19304
rect 3424 19261 3433 19295
rect 3433 19261 3467 19295
rect 3467 19261 3476 19295
rect 3424 19252 3476 19261
rect 3516 19252 3568 19304
rect 3792 19295 3844 19304
rect 3792 19261 3801 19295
rect 3801 19261 3835 19295
rect 3835 19261 3844 19295
rect 3792 19252 3844 19261
rect 3976 19295 4028 19304
rect 3976 19261 3985 19295
rect 3985 19261 4019 19295
rect 4019 19261 4028 19295
rect 3976 19252 4028 19261
rect 4068 19252 4120 19304
rect 2964 19184 3016 19236
rect 4528 19252 4580 19304
rect 5448 19456 5500 19508
rect 5540 19456 5592 19508
rect 8668 19456 8720 19508
rect 8852 19456 8904 19508
rect 9772 19456 9824 19508
rect 10416 19499 10468 19508
rect 10416 19465 10425 19499
rect 10425 19465 10459 19499
rect 10459 19465 10468 19499
rect 10416 19456 10468 19465
rect 12808 19456 12860 19508
rect 7932 19320 7984 19372
rect 8208 19320 8260 19372
rect 9404 19363 9456 19372
rect 9404 19329 9413 19363
rect 9413 19329 9447 19363
rect 9447 19329 9456 19363
rect 9404 19320 9456 19329
rect 9588 19320 9640 19372
rect 9680 19320 9732 19372
rect 10784 19388 10836 19440
rect 11888 19388 11940 19440
rect 13820 19456 13872 19508
rect 14372 19499 14424 19508
rect 14372 19465 14381 19499
rect 14381 19465 14415 19499
rect 14415 19465 14424 19499
rect 14372 19456 14424 19465
rect 14832 19456 14884 19508
rect 15292 19456 15344 19508
rect 20444 19456 20496 19508
rect 20720 19499 20772 19508
rect 20720 19465 20729 19499
rect 20729 19465 20763 19499
rect 20763 19465 20772 19499
rect 20720 19456 20772 19465
rect 6828 19295 6880 19304
rect 6828 19261 6837 19295
rect 6837 19261 6871 19295
rect 6871 19261 6880 19295
rect 6828 19252 6880 19261
rect 3056 19159 3108 19168
rect 3056 19125 3065 19159
rect 3065 19125 3099 19159
rect 3099 19125 3108 19159
rect 3056 19116 3108 19125
rect 4252 19159 4304 19168
rect 4252 19125 4261 19159
rect 4261 19125 4295 19159
rect 4295 19125 4304 19159
rect 4252 19116 4304 19125
rect 5816 19184 5868 19236
rect 6368 19184 6420 19236
rect 6920 19184 6972 19236
rect 7196 19184 7248 19236
rect 9864 19252 9916 19304
rect 9956 19295 10008 19304
rect 9956 19261 9965 19295
rect 9965 19261 9999 19295
rect 9999 19261 10008 19295
rect 9956 19252 10008 19261
rect 10048 19295 10100 19304
rect 10048 19261 10057 19295
rect 10057 19261 10091 19295
rect 10091 19261 10100 19295
rect 10048 19252 10100 19261
rect 8668 19184 8720 19236
rect 4804 19116 4856 19168
rect 5172 19116 5224 19168
rect 8208 19159 8260 19168
rect 8208 19125 8217 19159
rect 8217 19125 8251 19159
rect 8251 19125 8260 19159
rect 8208 19116 8260 19125
rect 8760 19159 8812 19168
rect 8760 19125 8785 19159
rect 8785 19125 8812 19159
rect 8760 19116 8812 19125
rect 9036 19159 9088 19168
rect 9036 19125 9045 19159
rect 9045 19125 9079 19159
rect 9079 19125 9088 19159
rect 9036 19116 9088 19125
rect 9220 19184 9272 19236
rect 10140 19184 10192 19236
rect 10508 19320 10560 19372
rect 11796 19320 11848 19372
rect 9864 19116 9916 19168
rect 11152 19116 11204 19168
rect 11796 19227 11848 19236
rect 11796 19193 11805 19227
rect 11805 19193 11839 19227
rect 11839 19193 11848 19227
rect 11796 19184 11848 19193
rect 11888 19227 11940 19236
rect 11888 19193 11897 19227
rect 11897 19193 11931 19227
rect 11931 19193 11940 19227
rect 11888 19184 11940 19193
rect 12072 19227 12124 19236
rect 12072 19193 12097 19227
rect 12097 19193 12124 19227
rect 12072 19184 12124 19193
rect 11980 19116 12032 19168
rect 12440 19116 12492 19168
rect 12900 19159 12952 19168
rect 12900 19125 12909 19159
rect 12909 19125 12943 19159
rect 12943 19125 12952 19159
rect 12900 19116 12952 19125
rect 14004 19295 14056 19304
rect 14004 19261 14013 19295
rect 14013 19261 14047 19295
rect 14047 19261 14056 19295
rect 14004 19252 14056 19261
rect 15200 19252 15252 19304
rect 20260 19388 20312 19440
rect 16120 19295 16172 19304
rect 16120 19261 16129 19295
rect 16129 19261 16163 19295
rect 16163 19261 16172 19295
rect 18144 19320 18196 19372
rect 16120 19252 16172 19261
rect 14924 19227 14976 19236
rect 14372 19159 14424 19168
rect 14372 19125 14381 19159
rect 14381 19125 14415 19159
rect 14415 19125 14424 19159
rect 14372 19116 14424 19125
rect 14924 19193 14958 19227
rect 14958 19193 14976 19227
rect 14924 19184 14976 19193
rect 15568 19184 15620 19236
rect 15752 19184 15804 19236
rect 16488 19184 16540 19236
rect 17868 19295 17920 19304
rect 17868 19261 17877 19295
rect 17877 19261 17911 19295
rect 17911 19261 17920 19295
rect 17868 19252 17920 19261
rect 18512 19252 18564 19304
rect 20260 19252 20312 19304
rect 20536 19320 20588 19372
rect 21180 19320 21232 19372
rect 22008 19456 22060 19508
rect 21824 19388 21876 19440
rect 21732 19320 21784 19372
rect 20628 19252 20680 19304
rect 20720 19252 20772 19304
rect 20996 19295 21048 19304
rect 20996 19261 21005 19295
rect 21005 19261 21039 19295
rect 21039 19261 21048 19295
rect 20996 19252 21048 19261
rect 21088 19252 21140 19304
rect 21548 19252 21600 19304
rect 16580 19116 16632 19168
rect 16856 19116 16908 19168
rect 17684 19116 17736 19168
rect 18788 19184 18840 19236
rect 18972 19227 19024 19236
rect 18972 19193 19006 19227
rect 19006 19193 19024 19227
rect 18972 19184 19024 19193
rect 19064 19184 19116 19236
rect 19248 19116 19300 19168
rect 19432 19116 19484 19168
rect 19708 19116 19760 19168
rect 21364 19116 21416 19168
rect 21732 19184 21784 19236
rect 22100 19295 22152 19304
rect 22100 19261 22109 19295
rect 22109 19261 22143 19295
rect 22143 19261 22152 19295
rect 22100 19252 22152 19261
rect 22468 19252 22520 19304
rect 22008 19116 22060 19168
rect 22192 19116 22244 19168
rect 22376 19116 22428 19168
rect 23112 19116 23164 19168
rect 4366 19014 4418 19066
rect 4430 19014 4482 19066
rect 4494 19014 4546 19066
rect 4558 19014 4610 19066
rect 4622 19014 4674 19066
rect 4686 19014 4738 19066
rect 10366 19014 10418 19066
rect 10430 19014 10482 19066
rect 10494 19014 10546 19066
rect 10558 19014 10610 19066
rect 10622 19014 10674 19066
rect 10686 19014 10738 19066
rect 16366 19014 16418 19066
rect 16430 19014 16482 19066
rect 16494 19014 16546 19066
rect 16558 19014 16610 19066
rect 16622 19014 16674 19066
rect 16686 19014 16738 19066
rect 22366 19014 22418 19066
rect 22430 19014 22482 19066
rect 22494 19014 22546 19066
rect 22558 19014 22610 19066
rect 22622 19014 22674 19066
rect 22686 19014 22738 19066
rect 2412 18776 2464 18828
rect 3056 18912 3108 18964
rect 3240 18912 3292 18964
rect 3976 18912 4028 18964
rect 6184 18955 6236 18964
rect 6184 18921 6193 18955
rect 6193 18921 6227 18955
rect 6227 18921 6236 18955
rect 6184 18912 6236 18921
rect 7288 18912 7340 18964
rect 9312 18912 9364 18964
rect 10048 18912 10100 18964
rect 4896 18844 4948 18896
rect 5264 18844 5316 18896
rect 1952 18751 2004 18760
rect 1952 18717 1961 18751
rect 1961 18717 1995 18751
rect 1995 18717 2004 18751
rect 1952 18708 2004 18717
rect 2596 18708 2648 18760
rect 4988 18776 5040 18828
rect 5172 18776 5224 18828
rect 5632 18776 5684 18828
rect 5816 18819 5868 18828
rect 5816 18785 5831 18819
rect 5831 18785 5865 18819
rect 5865 18785 5868 18819
rect 5816 18776 5868 18785
rect 7840 18844 7892 18896
rect 8484 18887 8536 18896
rect 8484 18853 8493 18887
rect 8493 18853 8527 18887
rect 8527 18853 8536 18887
rect 8484 18844 8536 18853
rect 8668 18844 8720 18896
rect 4252 18708 4304 18760
rect 4804 18708 4856 18760
rect 8300 18819 8352 18828
rect 8300 18785 8309 18819
rect 8309 18785 8343 18819
rect 8343 18785 8352 18819
rect 8300 18776 8352 18785
rect 8576 18776 8628 18828
rect 10140 18844 10192 18896
rect 8944 18776 8996 18828
rect 9220 18776 9272 18828
rect 9956 18776 10008 18828
rect 10508 18819 10560 18828
rect 12532 18912 12584 18964
rect 12900 18955 12952 18964
rect 12900 18921 12909 18955
rect 12909 18921 12943 18955
rect 12943 18921 12952 18955
rect 12900 18912 12952 18921
rect 13452 18912 13504 18964
rect 14004 18912 14056 18964
rect 14372 18955 14424 18964
rect 14372 18921 14381 18955
rect 14381 18921 14415 18955
rect 14415 18921 14424 18955
rect 14372 18912 14424 18921
rect 15292 18887 15344 18896
rect 15292 18853 15301 18887
rect 15301 18853 15335 18887
rect 15335 18853 15344 18887
rect 15292 18844 15344 18853
rect 10508 18785 10526 18819
rect 10526 18785 10560 18819
rect 10508 18776 10560 18785
rect 10968 18776 11020 18828
rect 11060 18776 11112 18828
rect 11980 18819 12032 18828
rect 11980 18785 11989 18819
rect 11989 18785 12023 18819
rect 12023 18785 12032 18819
rect 11980 18776 12032 18785
rect 12072 18819 12124 18828
rect 12072 18785 12081 18819
rect 12081 18785 12115 18819
rect 12115 18785 12124 18819
rect 12072 18776 12124 18785
rect 12348 18819 12400 18828
rect 12348 18785 12357 18819
rect 12357 18785 12391 18819
rect 12391 18785 12400 18819
rect 12348 18776 12400 18785
rect 12440 18819 12492 18828
rect 12440 18785 12449 18819
rect 12449 18785 12483 18819
rect 12483 18785 12492 18819
rect 12440 18776 12492 18785
rect 12532 18776 12584 18828
rect 13176 18776 13228 18828
rect 13452 18776 13504 18828
rect 13912 18776 13964 18828
rect 6460 18708 6512 18760
rect 7196 18751 7248 18760
rect 7196 18717 7205 18751
rect 7205 18717 7239 18751
rect 7239 18717 7248 18751
rect 7196 18708 7248 18717
rect 9404 18708 9456 18760
rect 5264 18683 5316 18692
rect 5264 18649 5273 18683
rect 5273 18649 5307 18683
rect 5307 18649 5316 18683
rect 5264 18640 5316 18649
rect 5448 18640 5500 18692
rect 8024 18640 8076 18692
rect 4896 18615 4948 18624
rect 4896 18581 4905 18615
rect 4905 18581 4939 18615
rect 4939 18581 4948 18615
rect 4896 18572 4948 18581
rect 5724 18572 5776 18624
rect 6092 18572 6144 18624
rect 6184 18572 6236 18624
rect 8576 18572 8628 18624
rect 9312 18572 9364 18624
rect 9404 18615 9456 18624
rect 9404 18581 9413 18615
rect 9413 18581 9447 18615
rect 9447 18581 9456 18615
rect 9404 18572 9456 18581
rect 10416 18572 10468 18624
rect 11520 18683 11572 18692
rect 11520 18649 11529 18683
rect 11529 18649 11563 18683
rect 11563 18649 11572 18683
rect 11520 18640 11572 18649
rect 11796 18640 11848 18692
rect 12072 18640 12124 18692
rect 13820 18708 13872 18760
rect 14372 18776 14424 18828
rect 12808 18572 12860 18624
rect 13176 18572 13228 18624
rect 15752 18955 15804 18964
rect 15752 18921 15761 18955
rect 15761 18921 15795 18955
rect 15795 18921 15804 18955
rect 15752 18912 15804 18921
rect 16856 18912 16908 18964
rect 17040 18955 17092 18964
rect 17040 18921 17049 18955
rect 17049 18921 17083 18955
rect 17083 18921 17092 18955
rect 17040 18912 17092 18921
rect 17776 18912 17828 18964
rect 17960 18955 18012 18964
rect 17960 18921 17969 18955
rect 17969 18921 18003 18955
rect 18003 18921 18012 18955
rect 17960 18912 18012 18921
rect 16948 18776 17000 18828
rect 17316 18819 17368 18828
rect 17316 18785 17325 18819
rect 17325 18785 17359 18819
rect 17359 18785 17368 18819
rect 17316 18776 17368 18785
rect 17592 18819 17644 18828
rect 17592 18785 17601 18819
rect 17601 18785 17635 18819
rect 17635 18785 17644 18819
rect 17592 18776 17644 18785
rect 18972 18912 19024 18964
rect 18328 18844 18380 18896
rect 20444 18912 20496 18964
rect 20904 18912 20956 18964
rect 21732 18912 21784 18964
rect 22284 18912 22336 18964
rect 22928 18912 22980 18964
rect 19248 18844 19300 18896
rect 19432 18819 19484 18828
rect 15936 18708 15988 18760
rect 19432 18785 19441 18819
rect 19441 18785 19475 18819
rect 19475 18785 19484 18819
rect 19432 18776 19484 18785
rect 18972 18708 19024 18760
rect 19892 18819 19944 18828
rect 19892 18785 19901 18819
rect 19901 18785 19935 18819
rect 19935 18785 19944 18819
rect 19892 18776 19944 18785
rect 20536 18819 20588 18828
rect 20536 18785 20545 18819
rect 20545 18785 20579 18819
rect 20579 18785 20588 18819
rect 20536 18776 20588 18785
rect 21088 18844 21140 18896
rect 22100 18844 22152 18896
rect 21180 18776 21232 18828
rect 20168 18708 20220 18760
rect 20444 18751 20496 18760
rect 20444 18717 20453 18751
rect 20453 18717 20487 18751
rect 20487 18717 20496 18751
rect 20444 18708 20496 18717
rect 20996 18708 21048 18760
rect 20076 18640 20128 18692
rect 22928 18776 22980 18828
rect 16948 18572 17000 18624
rect 17592 18572 17644 18624
rect 17868 18572 17920 18624
rect 19984 18572 20036 18624
rect 21732 18572 21784 18624
rect 1366 18470 1418 18522
rect 1430 18470 1482 18522
rect 1494 18470 1546 18522
rect 1558 18470 1610 18522
rect 1622 18470 1674 18522
rect 1686 18470 1738 18522
rect 7366 18470 7418 18522
rect 7430 18470 7482 18522
rect 7494 18470 7546 18522
rect 7558 18470 7610 18522
rect 7622 18470 7674 18522
rect 7686 18470 7738 18522
rect 13366 18470 13418 18522
rect 13430 18470 13482 18522
rect 13494 18470 13546 18522
rect 13558 18470 13610 18522
rect 13622 18470 13674 18522
rect 13686 18470 13738 18522
rect 19366 18470 19418 18522
rect 19430 18470 19482 18522
rect 19494 18470 19546 18522
rect 19558 18470 19610 18522
rect 19622 18470 19674 18522
rect 19686 18470 19738 18522
rect 2320 18368 2372 18420
rect 3976 18368 4028 18420
rect 6460 18411 6512 18420
rect 6460 18377 6469 18411
rect 6469 18377 6503 18411
rect 6503 18377 6512 18411
rect 6460 18368 6512 18377
rect 2044 18300 2096 18352
rect 4896 18300 4948 18352
rect 5816 18300 5868 18352
rect 5908 18343 5960 18352
rect 5908 18309 5917 18343
rect 5917 18309 5951 18343
rect 5951 18309 5960 18343
rect 5908 18300 5960 18309
rect 7288 18368 7340 18420
rect 8760 18368 8812 18420
rect 1952 18164 2004 18216
rect 2964 18232 3016 18284
rect 4160 18232 4212 18284
rect 2780 18164 2832 18216
rect 2228 18096 2280 18148
rect 2688 18096 2740 18148
rect 4068 18164 4120 18216
rect 5172 18232 5224 18284
rect 5264 18232 5316 18284
rect 4252 18139 4304 18148
rect 4252 18105 4261 18139
rect 4261 18105 4295 18139
rect 4295 18105 4304 18139
rect 4252 18096 4304 18105
rect 1768 18071 1820 18080
rect 1768 18037 1777 18071
rect 1777 18037 1811 18071
rect 1811 18037 1820 18071
rect 1768 18028 1820 18037
rect 3056 18028 3108 18080
rect 3884 18028 3936 18080
rect 4804 18028 4856 18080
rect 4896 18071 4948 18080
rect 4896 18037 4905 18071
rect 4905 18037 4939 18071
rect 4939 18037 4948 18071
rect 4896 18028 4948 18037
rect 4988 18028 5040 18080
rect 6092 18164 6144 18216
rect 6184 18207 6236 18216
rect 6184 18173 6193 18207
rect 6193 18173 6227 18207
rect 6227 18173 6236 18207
rect 6184 18164 6236 18173
rect 6920 18164 6972 18216
rect 7196 18164 7248 18216
rect 6368 18096 6420 18148
rect 6828 18096 6880 18148
rect 7380 18207 7432 18216
rect 7380 18173 7389 18207
rect 7389 18173 7423 18207
rect 7423 18173 7432 18207
rect 7380 18164 7432 18173
rect 7472 18207 7524 18216
rect 7472 18173 7481 18207
rect 7481 18173 7515 18207
rect 7515 18173 7524 18207
rect 7472 18164 7524 18173
rect 7656 18164 7708 18216
rect 8392 18300 8444 18352
rect 7932 18207 7984 18216
rect 7932 18173 7941 18207
rect 7941 18173 7975 18207
rect 7975 18173 7984 18207
rect 7932 18164 7984 18173
rect 8024 18207 8076 18216
rect 8024 18173 8033 18207
rect 8033 18173 8067 18207
rect 8067 18173 8076 18207
rect 8024 18164 8076 18173
rect 9680 18300 9732 18352
rect 10508 18368 10560 18420
rect 11704 18368 11756 18420
rect 11428 18300 11480 18352
rect 9496 18164 9548 18216
rect 11336 18232 11388 18284
rect 5724 18071 5776 18080
rect 5724 18037 5733 18071
rect 5733 18037 5767 18071
rect 5767 18037 5776 18071
rect 5724 18028 5776 18037
rect 5816 18028 5868 18080
rect 6276 18028 6328 18080
rect 6920 18028 6972 18080
rect 7196 18028 7248 18080
rect 8760 18096 8812 18148
rect 9588 18139 9640 18148
rect 9588 18105 9597 18139
rect 9597 18105 9631 18139
rect 9631 18105 9640 18139
rect 9588 18096 9640 18105
rect 10416 18164 10468 18216
rect 11704 18207 11756 18216
rect 11704 18173 11713 18207
rect 11713 18173 11747 18207
rect 11747 18173 11756 18207
rect 11704 18164 11756 18173
rect 10140 18096 10192 18148
rect 11060 18096 11112 18148
rect 12348 18368 12400 18420
rect 14188 18368 14240 18420
rect 14740 18300 14792 18352
rect 15292 18368 15344 18420
rect 17592 18368 17644 18420
rect 16120 18232 16172 18284
rect 16856 18232 16908 18284
rect 14188 18207 14240 18216
rect 14188 18173 14197 18207
rect 14197 18173 14231 18207
rect 14231 18173 14240 18207
rect 14188 18164 14240 18173
rect 15108 18207 15160 18216
rect 15108 18173 15117 18207
rect 15117 18173 15151 18207
rect 15151 18173 15160 18207
rect 15108 18164 15160 18173
rect 15568 18164 15620 18216
rect 17040 18164 17092 18216
rect 18052 18232 18104 18284
rect 17500 18164 17552 18216
rect 18420 18368 18472 18420
rect 18880 18300 18932 18352
rect 21088 18411 21140 18420
rect 21088 18377 21097 18411
rect 21097 18377 21131 18411
rect 21131 18377 21140 18411
rect 21088 18368 21140 18377
rect 21364 18300 21416 18352
rect 18512 18207 18564 18216
rect 18512 18173 18521 18207
rect 18521 18173 18555 18207
rect 18555 18173 18564 18207
rect 18512 18164 18564 18173
rect 18788 18232 18840 18284
rect 19984 18164 20036 18216
rect 20076 18164 20128 18216
rect 21456 18232 21508 18284
rect 8024 18028 8076 18080
rect 8944 18028 8996 18080
rect 9128 18028 9180 18080
rect 9772 18071 9824 18080
rect 9772 18037 9781 18071
rect 9781 18037 9815 18071
rect 9815 18037 9824 18071
rect 9772 18028 9824 18037
rect 11520 18028 11572 18080
rect 13820 18096 13872 18148
rect 13912 18139 13964 18148
rect 13912 18105 13921 18139
rect 13921 18105 13955 18139
rect 13955 18105 13964 18139
rect 13912 18096 13964 18105
rect 15200 18096 15252 18148
rect 17316 18096 17368 18148
rect 17960 18096 18012 18148
rect 12992 18028 13044 18080
rect 14372 18071 14424 18080
rect 14372 18037 14381 18071
rect 14381 18037 14415 18071
rect 14415 18037 14424 18071
rect 14372 18028 14424 18037
rect 14832 18028 14884 18080
rect 15752 18028 15804 18080
rect 15844 18028 15896 18080
rect 18420 18028 18472 18080
rect 18696 18139 18748 18148
rect 18696 18105 18705 18139
rect 18705 18105 18739 18139
rect 18739 18105 18748 18139
rect 18696 18096 18748 18105
rect 18880 18139 18932 18148
rect 18880 18105 18889 18139
rect 18889 18105 18923 18139
rect 18923 18105 18932 18139
rect 18880 18096 18932 18105
rect 19156 18071 19208 18080
rect 19156 18037 19165 18071
rect 19165 18037 19199 18071
rect 19199 18037 19208 18071
rect 19156 18028 19208 18037
rect 20904 18028 20956 18080
rect 21456 18071 21508 18080
rect 21456 18037 21465 18071
rect 21465 18037 21499 18071
rect 21499 18037 21508 18071
rect 21456 18028 21508 18037
rect 21548 18071 21600 18080
rect 21548 18037 21557 18071
rect 21557 18037 21591 18071
rect 21591 18037 21600 18071
rect 21548 18028 21600 18037
rect 23388 18028 23440 18080
rect 4366 17926 4418 17978
rect 4430 17926 4482 17978
rect 4494 17926 4546 17978
rect 4558 17926 4610 17978
rect 4622 17926 4674 17978
rect 4686 17926 4738 17978
rect 10366 17926 10418 17978
rect 10430 17926 10482 17978
rect 10494 17926 10546 17978
rect 10558 17926 10610 17978
rect 10622 17926 10674 17978
rect 10686 17926 10738 17978
rect 16366 17926 16418 17978
rect 16430 17926 16482 17978
rect 16494 17926 16546 17978
rect 16558 17926 16610 17978
rect 16622 17926 16674 17978
rect 16686 17926 16738 17978
rect 22366 17926 22418 17978
rect 22430 17926 22482 17978
rect 22494 17926 22546 17978
rect 22558 17926 22610 17978
rect 22622 17926 22674 17978
rect 22686 17926 22738 17978
rect 2320 17867 2372 17876
rect 2320 17833 2329 17867
rect 2329 17833 2363 17867
rect 2363 17833 2372 17867
rect 2320 17824 2372 17833
rect 2688 17867 2740 17876
rect 2688 17833 2697 17867
rect 2697 17833 2731 17867
rect 2731 17833 2740 17867
rect 2688 17824 2740 17833
rect 4160 17867 4212 17876
rect 4160 17833 4169 17867
rect 4169 17833 4203 17867
rect 4203 17833 4212 17867
rect 4160 17824 4212 17833
rect 5448 17824 5500 17876
rect 5724 17824 5776 17876
rect 6184 17867 6236 17876
rect 6184 17833 6193 17867
rect 6193 17833 6227 17867
rect 6227 17833 6236 17867
rect 6184 17824 6236 17833
rect 6368 17867 6420 17876
rect 6368 17833 6377 17867
rect 6377 17833 6411 17867
rect 6411 17833 6420 17867
rect 6368 17824 6420 17833
rect 6552 17824 6604 17876
rect 7840 17824 7892 17876
rect 7932 17824 7984 17876
rect 8760 17867 8812 17876
rect 8760 17833 8769 17867
rect 8769 17833 8803 17867
rect 8803 17833 8812 17867
rect 8760 17824 8812 17833
rect 9036 17824 9088 17876
rect 3884 17756 3936 17808
rect 5264 17799 5316 17808
rect 5264 17765 5273 17799
rect 5273 17765 5307 17799
rect 5307 17765 5316 17799
rect 5264 17756 5316 17765
rect 1216 17731 1268 17740
rect 1216 17697 1250 17731
rect 1250 17697 1268 17731
rect 1216 17688 1268 17697
rect 2872 17688 2924 17740
rect 3056 17731 3108 17740
rect 3056 17697 3090 17731
rect 3090 17697 3108 17731
rect 3056 17688 3108 17697
rect 848 17620 900 17672
rect 2688 17663 2740 17672
rect 2688 17629 2697 17663
rect 2697 17629 2731 17663
rect 2731 17629 2740 17663
rect 2688 17620 2740 17629
rect 2504 17527 2556 17536
rect 2504 17493 2513 17527
rect 2513 17493 2547 17527
rect 2547 17493 2556 17527
rect 2504 17484 2556 17493
rect 3884 17620 3936 17672
rect 4804 17688 4856 17740
rect 5356 17620 5408 17672
rect 3700 17484 3752 17536
rect 3792 17484 3844 17536
rect 6092 17688 6144 17740
rect 6828 17756 6880 17808
rect 7380 17799 7432 17808
rect 7380 17765 7389 17799
rect 7389 17765 7423 17799
rect 7423 17765 7432 17799
rect 7380 17756 7432 17765
rect 8024 17756 8076 17808
rect 8208 17756 8260 17808
rect 6368 17663 6420 17672
rect 6368 17629 6377 17663
rect 6377 17629 6411 17663
rect 6411 17629 6420 17663
rect 6368 17620 6420 17629
rect 6736 17595 6788 17604
rect 6736 17561 6745 17595
rect 6745 17561 6779 17595
rect 6779 17561 6788 17595
rect 6736 17552 6788 17561
rect 6092 17484 6144 17536
rect 8392 17731 8444 17740
rect 8392 17697 8401 17731
rect 8401 17697 8435 17731
rect 8435 17697 8444 17731
rect 8392 17688 8444 17697
rect 8484 17731 8536 17740
rect 8484 17697 8493 17731
rect 8493 17697 8527 17731
rect 8527 17697 8536 17731
rect 8484 17688 8536 17697
rect 8944 17731 8996 17740
rect 8944 17697 8953 17731
rect 8953 17697 8987 17731
rect 8987 17697 8996 17731
rect 8944 17688 8996 17697
rect 9312 17824 9364 17876
rect 13820 17824 13872 17876
rect 13176 17756 13228 17808
rect 14464 17756 14516 17808
rect 9680 17731 9732 17740
rect 9680 17697 9714 17731
rect 9714 17697 9732 17731
rect 9680 17688 9732 17697
rect 10968 17731 11020 17740
rect 10968 17697 10977 17731
rect 10977 17697 11011 17731
rect 11011 17697 11020 17731
rect 10968 17688 11020 17697
rect 11060 17688 11112 17740
rect 12716 17688 12768 17740
rect 12900 17731 12952 17740
rect 12900 17697 12909 17731
rect 12909 17697 12943 17731
rect 12943 17697 12952 17731
rect 12900 17688 12952 17697
rect 12992 17688 13044 17740
rect 7564 17663 7616 17672
rect 7564 17629 7573 17663
rect 7573 17629 7607 17663
rect 7607 17629 7616 17663
rect 7564 17620 7616 17629
rect 7932 17663 7984 17672
rect 7932 17629 7941 17663
rect 7941 17629 7975 17663
rect 7975 17629 7984 17663
rect 7932 17620 7984 17629
rect 8024 17663 8076 17672
rect 8024 17629 8033 17663
rect 8033 17629 8067 17663
rect 8067 17629 8076 17663
rect 8024 17620 8076 17629
rect 7840 17552 7892 17604
rect 12808 17663 12860 17672
rect 12808 17629 12817 17663
rect 12817 17629 12851 17663
rect 12851 17629 12860 17663
rect 12808 17620 12860 17629
rect 7196 17484 7248 17536
rect 7288 17484 7340 17536
rect 11980 17552 12032 17604
rect 14188 17688 14240 17740
rect 16948 17824 17000 17876
rect 17960 17867 18012 17876
rect 17960 17833 17987 17867
rect 17987 17833 18012 17867
rect 17960 17824 18012 17833
rect 18696 17824 18748 17876
rect 13912 17552 13964 17604
rect 12348 17527 12400 17536
rect 12348 17493 12357 17527
rect 12357 17493 12391 17527
rect 12391 17493 12400 17527
rect 12348 17484 12400 17493
rect 12440 17527 12492 17536
rect 12440 17493 12449 17527
rect 12449 17493 12483 17527
rect 12483 17493 12492 17527
rect 12440 17484 12492 17493
rect 12624 17484 12676 17536
rect 12992 17484 13044 17536
rect 14280 17484 14332 17536
rect 14556 17552 14608 17604
rect 15568 17731 15620 17740
rect 15568 17697 15577 17731
rect 15577 17697 15611 17731
rect 15611 17697 15620 17731
rect 15568 17688 15620 17697
rect 15752 17688 15804 17740
rect 15844 17731 15896 17740
rect 15844 17697 15853 17731
rect 15853 17697 15887 17731
rect 15887 17697 15896 17731
rect 15844 17688 15896 17697
rect 17040 17756 17092 17808
rect 18144 17799 18196 17808
rect 18144 17765 18153 17799
rect 18153 17765 18187 17799
rect 18187 17765 18196 17799
rect 18144 17756 18196 17765
rect 19156 17756 19208 17808
rect 19248 17756 19300 17808
rect 16948 17731 17000 17740
rect 16948 17697 16957 17731
rect 16957 17697 16991 17731
rect 16991 17697 17000 17731
rect 16948 17688 17000 17697
rect 18788 17731 18840 17740
rect 18788 17697 18797 17731
rect 18797 17697 18831 17731
rect 18831 17697 18840 17731
rect 18788 17688 18840 17697
rect 20720 17731 20772 17740
rect 20720 17697 20729 17731
rect 20729 17697 20763 17731
rect 20763 17697 20772 17731
rect 20720 17688 20772 17697
rect 20076 17620 20128 17672
rect 20812 17620 20864 17672
rect 17776 17552 17828 17604
rect 16028 17484 16080 17536
rect 17960 17527 18012 17536
rect 17960 17493 17969 17527
rect 17969 17493 18003 17527
rect 18003 17493 18012 17527
rect 17960 17484 18012 17493
rect 18512 17484 18564 17536
rect 19984 17484 20036 17536
rect 20076 17484 20128 17536
rect 22192 17824 22244 17876
rect 23296 17824 23348 17876
rect 22008 17756 22060 17808
rect 21364 17688 21416 17740
rect 21732 17688 21784 17740
rect 1366 17382 1418 17434
rect 1430 17382 1482 17434
rect 1494 17382 1546 17434
rect 1558 17382 1610 17434
rect 1622 17382 1674 17434
rect 1686 17382 1738 17434
rect 7366 17382 7418 17434
rect 7430 17382 7482 17434
rect 7494 17382 7546 17434
rect 7558 17382 7610 17434
rect 7622 17382 7674 17434
rect 7686 17382 7738 17434
rect 13366 17382 13418 17434
rect 13430 17382 13482 17434
rect 13494 17382 13546 17434
rect 13558 17382 13610 17434
rect 13622 17382 13674 17434
rect 13686 17382 13738 17434
rect 19366 17382 19418 17434
rect 19430 17382 19482 17434
rect 19494 17382 19546 17434
rect 19558 17382 19610 17434
rect 19622 17382 19674 17434
rect 19686 17382 19738 17434
rect 1216 17280 1268 17332
rect 2504 17280 2556 17332
rect 2780 17280 2832 17332
rect 2872 17323 2924 17332
rect 2872 17289 2881 17323
rect 2881 17289 2915 17323
rect 2915 17289 2924 17323
rect 2872 17280 2924 17289
rect 3056 17280 3108 17332
rect 6184 17323 6236 17332
rect 6184 17289 6193 17323
rect 6193 17289 6227 17323
rect 6227 17289 6236 17323
rect 6184 17280 6236 17289
rect 6368 17280 6420 17332
rect 5632 17212 5684 17264
rect 7104 17280 7156 17332
rect 7196 17280 7248 17332
rect 3608 17144 3660 17196
rect 1676 17076 1728 17128
rect 1952 17119 2004 17128
rect 1952 17085 1961 17119
rect 1961 17085 1995 17119
rect 1995 17085 2004 17119
rect 1952 17076 2004 17085
rect 2044 17119 2096 17128
rect 2044 17085 2053 17119
rect 2053 17085 2087 17119
rect 2087 17085 2096 17119
rect 2044 17076 2096 17085
rect 2872 17076 2924 17128
rect 2964 17076 3016 17128
rect 5540 17144 5592 17196
rect 6828 17212 6880 17264
rect 7932 17280 7984 17332
rect 8668 17280 8720 17332
rect 9588 17323 9640 17332
rect 9588 17289 9597 17323
rect 9597 17289 9631 17323
rect 9631 17289 9640 17323
rect 9588 17280 9640 17289
rect 11060 17280 11112 17332
rect 11428 17280 11480 17332
rect 11704 17280 11756 17332
rect 13820 17280 13872 17332
rect 13912 17280 13964 17332
rect 15568 17280 15620 17332
rect 16672 17280 16724 17332
rect 16948 17280 17000 17332
rect 18052 17280 18104 17332
rect 19892 17280 19944 17332
rect 21272 17280 21324 17332
rect 23388 17280 23440 17332
rect 2504 17008 2556 17060
rect 5080 17119 5132 17128
rect 5080 17085 5089 17119
rect 5089 17085 5123 17119
rect 5123 17085 5132 17119
rect 5080 17076 5132 17085
rect 5816 17076 5868 17128
rect 6368 17119 6420 17128
rect 6368 17085 6377 17119
rect 6377 17085 6411 17119
rect 6411 17085 6420 17119
rect 6368 17076 6420 17085
rect 1124 16983 1176 16992
rect 1124 16949 1133 16983
rect 1133 16949 1167 16983
rect 1167 16949 1176 16983
rect 1124 16940 1176 16949
rect 2872 16983 2924 16992
rect 2872 16949 2899 16983
rect 2899 16949 2924 16983
rect 2872 16940 2924 16949
rect 3700 16983 3752 16992
rect 3700 16949 3709 16983
rect 3709 16949 3743 16983
rect 3743 16949 3752 16983
rect 3700 16940 3752 16949
rect 5448 17051 5500 17060
rect 5448 17017 5457 17051
rect 5457 17017 5491 17051
rect 5491 17017 5500 17051
rect 5448 17008 5500 17017
rect 6276 17008 6328 17060
rect 9772 17212 9824 17264
rect 9312 17144 9364 17196
rect 6092 16940 6144 16992
rect 6736 16940 6788 16992
rect 7012 17051 7064 17060
rect 7012 17017 7021 17051
rect 7021 17017 7055 17051
rect 7055 17017 7064 17051
rect 7012 17008 7064 17017
rect 8576 16940 8628 16992
rect 8760 16983 8812 16992
rect 8760 16949 8769 16983
rect 8769 16949 8803 16983
rect 8803 16949 8812 16983
rect 8760 16940 8812 16949
rect 9588 17076 9640 17128
rect 10876 17144 10928 17196
rect 16764 17212 16816 17264
rect 18420 17212 18472 17264
rect 21364 17212 21416 17264
rect 12440 17144 12492 17196
rect 13176 17144 13228 17196
rect 9128 17008 9180 17060
rect 9956 17051 10008 17060
rect 9956 17017 9965 17051
rect 9965 17017 9999 17051
rect 9999 17017 10008 17051
rect 9956 17008 10008 17017
rect 9312 16940 9364 16992
rect 9588 16940 9640 16992
rect 13268 17076 13320 17128
rect 13912 17076 13964 17128
rect 14372 17076 14424 17128
rect 14924 17144 14976 17196
rect 16672 17144 16724 17196
rect 10784 17008 10836 17060
rect 11336 17051 11388 17060
rect 11336 17017 11361 17051
rect 11361 17017 11388 17051
rect 11336 17008 11388 17017
rect 12716 17008 12768 17060
rect 12992 17008 13044 17060
rect 13084 17008 13136 17060
rect 13636 17008 13688 17060
rect 14004 17051 14056 17060
rect 14004 17017 14013 17051
rect 14013 17017 14047 17051
rect 14047 17017 14056 17051
rect 14004 17008 14056 17017
rect 14740 17008 14792 17060
rect 15476 17076 15528 17128
rect 15752 17076 15804 17128
rect 14372 16983 14424 16992
rect 14372 16949 14381 16983
rect 14381 16949 14415 16983
rect 14415 16949 14424 16983
rect 14372 16940 14424 16949
rect 14556 16940 14608 16992
rect 15568 16983 15620 16992
rect 15568 16949 15577 16983
rect 15577 16949 15611 16983
rect 15611 16949 15620 16983
rect 15568 16940 15620 16949
rect 15936 16940 15988 16992
rect 16672 16983 16724 16992
rect 16672 16949 16681 16983
rect 16681 16949 16715 16983
rect 16715 16949 16724 16983
rect 16672 16940 16724 16949
rect 16856 16983 16908 16992
rect 16856 16949 16883 16983
rect 16883 16949 16908 16983
rect 16856 16940 16908 16949
rect 17408 17008 17460 17060
rect 17684 17051 17736 17060
rect 17684 17017 17693 17051
rect 17693 17017 17727 17051
rect 17727 17017 17736 17051
rect 17684 17008 17736 17017
rect 17224 16940 17276 16992
rect 18052 17076 18104 17128
rect 18328 17076 18380 17128
rect 18420 17119 18472 17128
rect 18420 17085 18429 17119
rect 18429 17085 18463 17119
rect 18463 17085 18472 17119
rect 18420 17076 18472 17085
rect 20812 17144 20864 17196
rect 21732 17076 21784 17128
rect 22192 17076 22244 17128
rect 19156 17051 19208 17060
rect 19156 17017 19165 17051
rect 19165 17017 19199 17051
rect 19199 17017 19208 17051
rect 19156 17008 19208 17017
rect 19340 17051 19392 17060
rect 19340 17017 19349 17051
rect 19349 17017 19383 17051
rect 19383 17017 19392 17051
rect 19340 17008 19392 17017
rect 19984 17008 20036 17060
rect 18328 16940 18380 16992
rect 18788 16940 18840 16992
rect 18880 16983 18932 16992
rect 18880 16949 18889 16983
rect 18889 16949 18923 16983
rect 18923 16949 18932 16983
rect 18880 16940 18932 16949
rect 4366 16838 4418 16890
rect 4430 16838 4482 16890
rect 4494 16838 4546 16890
rect 4558 16838 4610 16890
rect 4622 16838 4674 16890
rect 4686 16838 4738 16890
rect 10366 16838 10418 16890
rect 10430 16838 10482 16890
rect 10494 16838 10546 16890
rect 10558 16838 10610 16890
rect 10622 16838 10674 16890
rect 10686 16838 10738 16890
rect 16366 16838 16418 16890
rect 16430 16838 16482 16890
rect 16494 16838 16546 16890
rect 16558 16838 16610 16890
rect 16622 16838 16674 16890
rect 16686 16838 16738 16890
rect 22366 16838 22418 16890
rect 22430 16838 22482 16890
rect 22494 16838 22546 16890
rect 22558 16838 22610 16890
rect 22622 16838 22674 16890
rect 22686 16838 22738 16890
rect 848 16600 900 16652
rect 3884 16779 3936 16788
rect 3884 16745 3893 16779
rect 3893 16745 3927 16779
rect 3927 16745 3936 16779
rect 3884 16736 3936 16745
rect 3976 16736 4028 16788
rect 4344 16736 4396 16788
rect 4528 16736 4580 16788
rect 5080 16736 5132 16788
rect 5264 16736 5316 16788
rect 6644 16736 6696 16788
rect 7288 16736 7340 16788
rect 7840 16779 7892 16788
rect 7840 16745 7849 16779
rect 7849 16745 7883 16779
rect 7883 16745 7892 16779
rect 7840 16736 7892 16745
rect 8484 16736 8536 16788
rect 3700 16668 3752 16720
rect 2412 16643 2464 16652
rect 2412 16609 2421 16643
rect 2421 16609 2455 16643
rect 2455 16609 2464 16643
rect 2412 16600 2464 16609
rect 2504 16600 2556 16652
rect 2688 16643 2740 16652
rect 2688 16609 2697 16643
rect 2697 16609 2731 16643
rect 2731 16609 2740 16643
rect 2688 16600 2740 16609
rect 2320 16439 2372 16448
rect 2320 16405 2329 16439
rect 2329 16405 2363 16439
rect 2363 16405 2372 16439
rect 2320 16396 2372 16405
rect 2688 16396 2740 16448
rect 3516 16643 3568 16652
rect 3516 16609 3525 16643
rect 3525 16609 3559 16643
rect 3559 16609 3568 16643
rect 3516 16600 3568 16609
rect 3608 16643 3660 16652
rect 3608 16609 3617 16643
rect 3617 16609 3651 16643
rect 3651 16609 3660 16643
rect 3608 16600 3660 16609
rect 3792 16643 3844 16652
rect 3792 16609 3801 16643
rect 3801 16609 3835 16643
rect 3835 16609 3844 16643
rect 3792 16600 3844 16609
rect 4068 16643 4120 16652
rect 4068 16609 4077 16643
rect 4077 16609 4111 16643
rect 4111 16609 4120 16643
rect 4068 16600 4120 16609
rect 4252 16600 4304 16652
rect 5172 16600 5224 16652
rect 5632 16643 5684 16652
rect 5632 16609 5641 16643
rect 5641 16609 5675 16643
rect 5675 16609 5684 16643
rect 5632 16600 5684 16609
rect 5908 16600 5960 16652
rect 7012 16600 7064 16652
rect 7472 16643 7524 16652
rect 7472 16609 7481 16643
rect 7481 16609 7515 16643
rect 7515 16609 7524 16643
rect 7472 16600 7524 16609
rect 7748 16643 7800 16652
rect 7748 16609 7757 16643
rect 7757 16609 7791 16643
rect 7791 16609 7800 16643
rect 7748 16600 7800 16609
rect 9036 16736 9088 16788
rect 9956 16736 10008 16788
rect 8944 16668 8996 16720
rect 9312 16643 9364 16652
rect 9312 16609 9346 16643
rect 9346 16609 9364 16643
rect 9312 16600 9364 16609
rect 3332 16464 3384 16516
rect 8484 16532 8536 16584
rect 4804 16464 4856 16516
rect 3792 16396 3844 16448
rect 6460 16396 6512 16448
rect 6552 16396 6604 16448
rect 7748 16464 7800 16516
rect 12348 16736 12400 16788
rect 10600 16643 10652 16652
rect 10600 16609 10609 16643
rect 10609 16609 10643 16643
rect 10643 16609 10652 16643
rect 10600 16600 10652 16609
rect 10784 16643 10836 16652
rect 10784 16609 10793 16643
rect 10793 16609 10827 16643
rect 10827 16609 10836 16643
rect 10784 16600 10836 16609
rect 11336 16600 11388 16652
rect 11980 16643 12032 16652
rect 11980 16609 11989 16643
rect 11989 16609 12023 16643
rect 12023 16609 12032 16643
rect 11980 16600 12032 16609
rect 12256 16668 12308 16720
rect 13728 16736 13780 16788
rect 14372 16736 14424 16788
rect 12164 16643 12216 16652
rect 12164 16609 12173 16643
rect 12173 16609 12207 16643
rect 12207 16609 12216 16643
rect 12164 16600 12216 16609
rect 12348 16643 12400 16652
rect 12348 16609 12357 16643
rect 12357 16609 12391 16643
rect 12391 16609 12400 16643
rect 12348 16600 12400 16609
rect 12992 16600 13044 16652
rect 14924 16668 14976 16720
rect 13636 16643 13688 16652
rect 13636 16609 13645 16643
rect 13645 16609 13679 16643
rect 13679 16609 13688 16643
rect 13636 16600 13688 16609
rect 14004 16600 14056 16652
rect 14556 16643 14608 16652
rect 14556 16609 14565 16643
rect 14565 16609 14599 16643
rect 14599 16609 14608 16643
rect 14556 16600 14608 16609
rect 14832 16600 14884 16652
rect 15476 16736 15528 16788
rect 15568 16643 15620 16652
rect 15568 16609 15577 16643
rect 15577 16609 15611 16643
rect 15611 16609 15620 16643
rect 15568 16600 15620 16609
rect 10140 16532 10192 16584
rect 10692 16532 10744 16584
rect 13268 16532 13320 16584
rect 13728 16532 13780 16584
rect 16764 16668 16816 16720
rect 17132 16668 17184 16720
rect 15936 16600 15988 16652
rect 16212 16643 16264 16652
rect 16212 16609 16221 16643
rect 16221 16609 16255 16643
rect 16255 16609 16264 16643
rect 16212 16600 16264 16609
rect 17040 16643 17092 16652
rect 17040 16609 17049 16643
rect 17049 16609 17083 16643
rect 17083 16609 17092 16643
rect 17040 16600 17092 16609
rect 17224 16643 17276 16652
rect 17224 16609 17233 16643
rect 17233 16609 17267 16643
rect 17267 16609 17276 16643
rect 17224 16600 17276 16609
rect 17408 16643 17460 16652
rect 17408 16609 17417 16643
rect 17417 16609 17451 16643
rect 17451 16609 17460 16643
rect 17408 16600 17460 16609
rect 18420 16736 18472 16788
rect 18880 16668 18932 16720
rect 18788 16600 18840 16652
rect 21088 16736 21140 16788
rect 21180 16736 21232 16788
rect 22192 16736 22244 16788
rect 22744 16736 22796 16788
rect 23204 16736 23256 16788
rect 19892 16711 19944 16720
rect 19892 16677 19901 16711
rect 19901 16677 19935 16711
rect 19935 16677 19944 16711
rect 19892 16668 19944 16677
rect 20076 16711 20128 16720
rect 20076 16677 20085 16711
rect 20085 16677 20119 16711
rect 20119 16677 20128 16711
rect 20076 16668 20128 16677
rect 7104 16396 7156 16448
rect 9680 16396 9732 16448
rect 10416 16439 10468 16448
rect 10416 16405 10425 16439
rect 10425 16405 10459 16439
rect 10459 16405 10468 16439
rect 10416 16396 10468 16405
rect 10968 16396 11020 16448
rect 11520 16439 11572 16448
rect 11520 16405 11529 16439
rect 11529 16405 11563 16439
rect 11563 16405 11572 16439
rect 11520 16396 11572 16405
rect 11612 16439 11664 16448
rect 11612 16405 11621 16439
rect 11621 16405 11655 16439
rect 11655 16405 11664 16439
rect 11612 16396 11664 16405
rect 11980 16396 12032 16448
rect 12164 16396 12216 16448
rect 12808 16464 12860 16516
rect 12900 16507 12952 16516
rect 12900 16473 12909 16507
rect 12909 16473 12943 16507
rect 12943 16473 12952 16507
rect 12900 16464 12952 16473
rect 12992 16464 13044 16516
rect 18328 16507 18380 16516
rect 18328 16473 18337 16507
rect 18337 16473 18371 16507
rect 18371 16473 18380 16507
rect 18328 16464 18380 16473
rect 18512 16464 18564 16516
rect 19156 16464 19208 16516
rect 20720 16600 20772 16652
rect 21088 16600 21140 16652
rect 21732 16600 21784 16652
rect 22376 16600 22428 16652
rect 12716 16439 12768 16448
rect 12716 16405 12725 16439
rect 12725 16405 12759 16439
rect 12759 16405 12768 16439
rect 12716 16396 12768 16405
rect 13084 16396 13136 16448
rect 13360 16396 13412 16448
rect 15936 16439 15988 16448
rect 15936 16405 15945 16439
rect 15945 16405 15979 16439
rect 15979 16405 15988 16439
rect 15936 16396 15988 16405
rect 17500 16439 17552 16448
rect 17500 16405 17509 16439
rect 17509 16405 17543 16439
rect 17543 16405 17552 16439
rect 17500 16396 17552 16405
rect 19064 16439 19116 16448
rect 19064 16405 19073 16439
rect 19073 16405 19107 16439
rect 19107 16405 19116 16439
rect 19064 16396 19116 16405
rect 20076 16396 20128 16448
rect 20444 16439 20496 16448
rect 20444 16405 20453 16439
rect 20453 16405 20487 16439
rect 20487 16405 20496 16439
rect 20444 16396 20496 16405
rect 21088 16439 21140 16448
rect 21088 16405 21097 16439
rect 21097 16405 21131 16439
rect 21131 16405 21140 16439
rect 21088 16396 21140 16405
rect 1366 16294 1418 16346
rect 1430 16294 1482 16346
rect 1494 16294 1546 16346
rect 1558 16294 1610 16346
rect 1622 16294 1674 16346
rect 1686 16294 1738 16346
rect 7366 16294 7418 16346
rect 7430 16294 7482 16346
rect 7494 16294 7546 16346
rect 7558 16294 7610 16346
rect 7622 16294 7674 16346
rect 7686 16294 7738 16346
rect 13366 16294 13418 16346
rect 13430 16294 13482 16346
rect 13494 16294 13546 16346
rect 13558 16294 13610 16346
rect 13622 16294 13674 16346
rect 13686 16294 13738 16346
rect 19366 16294 19418 16346
rect 19430 16294 19482 16346
rect 19494 16294 19546 16346
rect 19558 16294 19610 16346
rect 19622 16294 19674 16346
rect 19686 16294 19738 16346
rect 2320 16192 2372 16244
rect 4988 16192 5040 16244
rect 5448 16192 5500 16244
rect 8208 16192 8260 16244
rect 8484 16192 8536 16244
rect 8760 16235 8812 16244
rect 8760 16201 8769 16235
rect 8769 16201 8803 16235
rect 8803 16201 8812 16235
rect 8760 16192 8812 16201
rect 2872 16124 2924 16176
rect 5632 16124 5684 16176
rect 6828 16124 6880 16176
rect 848 16099 900 16108
rect 848 16065 857 16099
rect 857 16065 891 16099
rect 891 16065 900 16099
rect 848 16056 900 16065
rect 2688 16056 2740 16108
rect 3056 16099 3108 16108
rect 3056 16065 3065 16099
rect 3065 16065 3099 16099
rect 3099 16065 3108 16099
rect 3056 16056 3108 16065
rect 4896 16099 4948 16108
rect 4896 16065 4905 16099
rect 4905 16065 4939 16099
rect 4939 16065 4948 16099
rect 4896 16056 4948 16065
rect 5724 16099 5776 16108
rect 5724 16065 5733 16099
rect 5733 16065 5767 16099
rect 5767 16065 5776 16099
rect 5724 16056 5776 16065
rect 1124 16031 1176 16040
rect 1124 15997 1158 16031
rect 1158 15997 1176 16031
rect 1124 15988 1176 15997
rect 2780 15988 2832 16040
rect 3240 16031 3292 16040
rect 3240 15997 3249 16031
rect 3249 15997 3283 16031
rect 3283 15997 3292 16031
rect 3240 15988 3292 15997
rect 3332 15988 3384 16040
rect 4988 15988 5040 16040
rect 2504 15852 2556 15904
rect 2780 15852 2832 15904
rect 4804 15920 4856 15972
rect 6184 15988 6236 16040
rect 4988 15895 5040 15904
rect 4988 15861 4997 15895
rect 4997 15861 5031 15895
rect 5031 15861 5040 15895
rect 4988 15852 5040 15861
rect 5264 15852 5316 15904
rect 5448 15895 5500 15904
rect 5448 15861 5457 15895
rect 5457 15861 5491 15895
rect 5491 15861 5500 15895
rect 5448 15852 5500 15861
rect 5724 15852 5776 15904
rect 6552 16031 6604 16040
rect 6552 15997 6561 16031
rect 6561 15997 6595 16031
rect 6595 15997 6604 16031
rect 6552 15988 6604 15997
rect 6736 16056 6788 16108
rect 6460 15920 6512 15972
rect 6920 15988 6972 16040
rect 7196 16056 7248 16108
rect 9680 16192 9732 16244
rect 9956 16192 10008 16244
rect 10600 16192 10652 16244
rect 10784 16192 10836 16244
rect 12256 16192 12308 16244
rect 15660 16192 15712 16244
rect 16212 16192 16264 16244
rect 18236 16192 18288 16244
rect 9772 16124 9824 16176
rect 17960 16124 18012 16176
rect 21180 16192 21232 16244
rect 22284 16192 22336 16244
rect 22928 16192 22980 16244
rect 20260 16124 20312 16176
rect 20996 16124 21048 16176
rect 21272 16124 21324 16176
rect 7840 15988 7892 16040
rect 8208 16031 8260 16040
rect 8208 15997 8217 16031
rect 8217 15997 8251 16031
rect 8251 15997 8260 16031
rect 8208 15988 8260 15997
rect 7196 15920 7248 15972
rect 9036 16031 9088 16040
rect 9036 15997 9045 16031
rect 9045 15997 9079 16031
rect 9079 15997 9088 16031
rect 9036 15988 9088 15997
rect 7288 15852 7340 15904
rect 9128 15920 9180 15972
rect 9680 15988 9732 16040
rect 10048 16031 10100 16040
rect 10048 15997 10057 16031
rect 10057 15997 10091 16031
rect 10091 15997 10100 16031
rect 10048 15988 10100 15997
rect 10232 16031 10284 16040
rect 10232 15997 10241 16031
rect 10241 15997 10275 16031
rect 10275 15997 10284 16031
rect 10232 15988 10284 15997
rect 10416 16056 10468 16108
rect 10140 15920 10192 15972
rect 7840 15852 7892 15904
rect 8024 15895 8076 15904
rect 8024 15861 8033 15895
rect 8033 15861 8067 15895
rect 8067 15861 8076 15895
rect 8024 15852 8076 15861
rect 8668 15852 8720 15904
rect 9404 15852 9456 15904
rect 11336 15895 11388 15904
rect 11336 15861 11345 15895
rect 11345 15861 11379 15895
rect 11379 15861 11388 15895
rect 11336 15852 11388 15861
rect 11796 16031 11848 16040
rect 11796 15997 11805 16031
rect 11805 15997 11839 16031
rect 11839 15997 11848 16031
rect 11796 15988 11848 15997
rect 12256 16056 12308 16108
rect 12716 16056 12768 16108
rect 12348 15988 12400 16040
rect 12992 16099 13044 16108
rect 12992 16065 13001 16099
rect 13001 16065 13035 16099
rect 13035 16065 13044 16099
rect 12992 16056 13044 16065
rect 13084 16056 13136 16108
rect 12256 15920 12308 15972
rect 13544 16031 13596 16040
rect 13544 15997 13553 16031
rect 13553 15997 13587 16031
rect 13587 15997 13596 16031
rect 13544 15988 13596 15997
rect 19064 16056 19116 16108
rect 22008 16124 22060 16176
rect 13820 15963 13872 15972
rect 13820 15929 13829 15963
rect 13829 15929 13863 15963
rect 13863 15929 13872 15963
rect 13820 15920 13872 15929
rect 16948 15988 17000 16040
rect 11980 15852 12032 15904
rect 15384 15920 15436 15972
rect 16120 15920 16172 15972
rect 14648 15852 14700 15904
rect 16212 15895 16264 15904
rect 16212 15861 16221 15895
rect 16221 15861 16255 15895
rect 16255 15861 16264 15895
rect 17408 15920 17460 15972
rect 19708 15988 19760 16040
rect 20076 16031 20128 16040
rect 20076 15997 20085 16031
rect 20085 15997 20119 16031
rect 20119 15997 20128 16031
rect 20076 15988 20128 15997
rect 20444 15988 20496 16040
rect 21364 16031 21416 16040
rect 21364 15997 21373 16031
rect 21373 15997 21407 16031
rect 21407 15997 21416 16031
rect 21364 15988 21416 15997
rect 22100 16056 22152 16108
rect 22192 16056 22244 16108
rect 21916 16031 21968 16040
rect 21916 15997 21925 16031
rect 21925 15997 21959 16031
rect 21959 15997 21968 16031
rect 21916 15988 21968 15997
rect 16212 15852 16264 15861
rect 17868 15852 17920 15904
rect 19432 15852 19484 15904
rect 22008 15920 22060 15972
rect 22376 15988 22428 16040
rect 22744 16031 22796 16040
rect 22744 15997 22753 16031
rect 22753 15997 22787 16031
rect 22787 15997 22796 16031
rect 22744 15988 22796 15997
rect 23112 15988 23164 16040
rect 23480 15920 23532 15972
rect 20352 15852 20404 15904
rect 21824 15852 21876 15904
rect 4366 15750 4418 15802
rect 4430 15750 4482 15802
rect 4494 15750 4546 15802
rect 4558 15750 4610 15802
rect 4622 15750 4674 15802
rect 4686 15750 4738 15802
rect 10366 15750 10418 15802
rect 10430 15750 10482 15802
rect 10494 15750 10546 15802
rect 10558 15750 10610 15802
rect 10622 15750 10674 15802
rect 10686 15750 10738 15802
rect 16366 15750 16418 15802
rect 16430 15750 16482 15802
rect 16494 15750 16546 15802
rect 16558 15750 16610 15802
rect 16622 15750 16674 15802
rect 16686 15750 16738 15802
rect 22366 15750 22418 15802
rect 22430 15750 22482 15802
rect 22494 15750 22546 15802
rect 22558 15750 22610 15802
rect 22622 15750 22674 15802
rect 22686 15750 22738 15802
rect 2964 15691 3016 15700
rect 2964 15657 2973 15691
rect 2973 15657 3007 15691
rect 3007 15657 3016 15691
rect 2964 15648 3016 15657
rect 3792 15691 3844 15700
rect 3792 15657 3801 15691
rect 3801 15657 3835 15691
rect 3835 15657 3844 15691
rect 3792 15648 3844 15657
rect 5448 15648 5500 15700
rect 6644 15648 6696 15700
rect 940 15580 992 15632
rect 1216 15623 1268 15632
rect 1216 15589 1225 15623
rect 1225 15589 1259 15623
rect 1259 15589 1268 15623
rect 1216 15580 1268 15589
rect 2780 15580 2832 15632
rect 3240 15580 3292 15632
rect 5540 15580 5592 15632
rect 1676 15555 1728 15564
rect 1676 15521 1685 15555
rect 1685 15521 1719 15555
rect 1719 15521 1728 15555
rect 1676 15512 1728 15521
rect 1952 15512 2004 15564
rect 2320 15512 2372 15564
rect 3608 15512 3660 15564
rect 6552 15512 6604 15564
rect 7104 15555 7156 15564
rect 7104 15521 7113 15555
rect 7113 15521 7147 15555
rect 7147 15521 7156 15555
rect 7104 15512 7156 15521
rect 7380 15648 7432 15700
rect 9496 15648 9548 15700
rect 8300 15580 8352 15632
rect 8484 15580 8536 15632
rect 9588 15580 9640 15632
rect 9956 15580 10008 15632
rect 7380 15555 7432 15564
rect 7380 15521 7389 15555
rect 7389 15521 7423 15555
rect 7423 15521 7432 15555
rect 7380 15512 7432 15521
rect 7932 15512 7984 15564
rect 9036 15512 9088 15564
rect 9680 15555 9732 15564
rect 9680 15521 9689 15555
rect 9689 15521 9723 15555
rect 9723 15521 9732 15555
rect 9680 15512 9732 15521
rect 9772 15512 9824 15564
rect 10048 15512 10100 15564
rect 10324 15512 10376 15564
rect 3332 15487 3384 15496
rect 3332 15453 3341 15487
rect 3341 15453 3375 15487
rect 3375 15453 3384 15487
rect 3332 15444 3384 15453
rect 1860 15376 1912 15428
rect 3148 15376 3200 15428
rect 5448 15444 5500 15496
rect 6276 15487 6328 15496
rect 6276 15453 6285 15487
rect 6285 15453 6319 15487
rect 6319 15453 6328 15487
rect 6276 15444 6328 15453
rect 9220 15487 9272 15496
rect 9220 15453 9229 15487
rect 9229 15453 9263 15487
rect 9263 15453 9272 15487
rect 9220 15444 9272 15453
rect 9312 15487 9364 15496
rect 9312 15453 9321 15487
rect 9321 15453 9355 15487
rect 9355 15453 9364 15487
rect 9312 15444 9364 15453
rect 9404 15487 9456 15496
rect 9404 15453 9413 15487
rect 9413 15453 9447 15487
rect 9447 15453 9456 15487
rect 9404 15444 9456 15453
rect 10140 15444 10192 15496
rect 10416 15444 10468 15496
rect 3056 15308 3108 15360
rect 6460 15376 6512 15428
rect 6920 15376 6972 15428
rect 8208 15376 8260 15428
rect 9588 15376 9640 15428
rect 10232 15376 10284 15428
rect 6368 15308 6420 15360
rect 8116 15351 8168 15360
rect 8116 15317 8125 15351
rect 8125 15317 8159 15351
rect 8159 15317 8168 15351
rect 8116 15308 8168 15317
rect 8300 15308 8352 15360
rect 8852 15308 8904 15360
rect 9404 15308 9456 15360
rect 11796 15648 11848 15700
rect 10968 15555 11020 15564
rect 10968 15521 10977 15555
rect 10977 15521 11011 15555
rect 11011 15521 11020 15555
rect 10968 15512 11020 15521
rect 12164 15580 12216 15632
rect 12440 15555 12492 15564
rect 12440 15521 12449 15555
rect 12449 15521 12483 15555
rect 12483 15521 12492 15555
rect 12440 15512 12492 15521
rect 10692 15444 10744 15496
rect 11336 15444 11388 15496
rect 11796 15444 11848 15496
rect 13544 15648 13596 15700
rect 13820 15648 13872 15700
rect 15200 15648 15252 15700
rect 17592 15648 17644 15700
rect 18052 15648 18104 15700
rect 16212 15580 16264 15632
rect 17408 15580 17460 15632
rect 13820 15555 13872 15564
rect 13820 15521 13829 15555
rect 13829 15521 13863 15555
rect 13863 15521 13872 15555
rect 13820 15512 13872 15521
rect 13912 15444 13964 15496
rect 14832 15512 14884 15564
rect 15016 15555 15068 15564
rect 15016 15521 15025 15555
rect 15025 15521 15059 15555
rect 15059 15521 15068 15555
rect 15016 15512 15068 15521
rect 15660 15555 15712 15564
rect 15660 15521 15669 15555
rect 15669 15521 15703 15555
rect 15703 15521 15712 15555
rect 15660 15512 15712 15521
rect 15752 15512 15804 15564
rect 10876 15376 10928 15428
rect 12256 15376 12308 15428
rect 14096 15376 14148 15428
rect 14924 15376 14976 15428
rect 15108 15376 15160 15428
rect 15476 15376 15528 15428
rect 16120 15444 16172 15496
rect 17132 15444 17184 15496
rect 12716 15308 12768 15360
rect 12992 15308 13044 15360
rect 15016 15308 15068 15360
rect 16488 15308 16540 15360
rect 16764 15308 16816 15360
rect 17408 15487 17460 15496
rect 17408 15453 17417 15487
rect 17417 15453 17451 15487
rect 17451 15453 17460 15487
rect 17408 15444 17460 15453
rect 17868 15555 17920 15564
rect 17868 15521 17877 15555
rect 17877 15521 17911 15555
rect 17911 15521 17920 15555
rect 17868 15512 17920 15521
rect 19432 15555 19484 15564
rect 18236 15444 18288 15496
rect 18696 15487 18748 15496
rect 18696 15453 18705 15487
rect 18705 15453 18739 15487
rect 18739 15453 18748 15487
rect 18696 15444 18748 15453
rect 19432 15521 19441 15555
rect 19441 15521 19475 15555
rect 19475 15521 19484 15555
rect 19432 15512 19484 15521
rect 19708 15512 19760 15564
rect 20168 15580 20220 15632
rect 22468 15648 22520 15700
rect 22836 15691 22888 15700
rect 22836 15657 22845 15691
rect 22845 15657 22879 15691
rect 22879 15657 22888 15691
rect 22836 15648 22888 15657
rect 20812 15512 20864 15564
rect 21088 15555 21140 15564
rect 21088 15521 21097 15555
rect 21097 15521 21131 15555
rect 21131 15521 21140 15555
rect 21088 15512 21140 15521
rect 19156 15376 19208 15428
rect 20444 15444 20496 15496
rect 20536 15376 20588 15428
rect 21088 15376 21140 15428
rect 21824 15555 21876 15564
rect 21824 15521 21833 15555
rect 21833 15521 21867 15555
rect 21867 15521 21876 15555
rect 21824 15512 21876 15521
rect 22008 15555 22060 15564
rect 22008 15521 22017 15555
rect 22017 15521 22051 15555
rect 22051 15521 22060 15555
rect 22008 15512 22060 15521
rect 22100 15512 22152 15564
rect 22284 15555 22336 15564
rect 22284 15521 22293 15555
rect 22293 15521 22327 15555
rect 22327 15521 22336 15555
rect 22284 15512 22336 15521
rect 23020 15555 23072 15564
rect 23020 15521 23029 15555
rect 23029 15521 23063 15555
rect 23063 15521 23072 15555
rect 23020 15512 23072 15521
rect 22284 15376 22336 15428
rect 19248 15308 19300 15360
rect 20260 15351 20312 15360
rect 20260 15317 20269 15351
rect 20269 15317 20303 15351
rect 20303 15317 20312 15351
rect 20260 15308 20312 15317
rect 20352 15308 20404 15360
rect 20720 15308 20772 15360
rect 22560 15351 22612 15360
rect 22560 15317 22569 15351
rect 22569 15317 22603 15351
rect 22603 15317 22612 15351
rect 22560 15308 22612 15317
rect 1366 15206 1418 15258
rect 1430 15206 1482 15258
rect 1494 15206 1546 15258
rect 1558 15206 1610 15258
rect 1622 15206 1674 15258
rect 1686 15206 1738 15258
rect 7366 15206 7418 15258
rect 7430 15206 7482 15258
rect 7494 15206 7546 15258
rect 7558 15206 7610 15258
rect 7622 15206 7674 15258
rect 7686 15206 7738 15258
rect 13366 15206 13418 15258
rect 13430 15206 13482 15258
rect 13494 15206 13546 15258
rect 13558 15206 13610 15258
rect 13622 15206 13674 15258
rect 13686 15206 13738 15258
rect 19366 15206 19418 15258
rect 19430 15206 19482 15258
rect 19494 15206 19546 15258
rect 19558 15206 19610 15258
rect 19622 15206 19674 15258
rect 19686 15206 19738 15258
rect 2504 15104 2556 15156
rect 1216 14900 1268 14952
rect 3240 15036 3292 15088
rect 4712 15104 4764 15156
rect 6552 15104 6604 15156
rect 7196 15104 7248 15156
rect 2504 15011 2556 15020
rect 2504 14977 2513 15011
rect 2513 14977 2547 15011
rect 2547 14977 2556 15011
rect 2504 14968 2556 14977
rect 2872 14968 2924 15020
rect 2596 14943 2648 14952
rect 2596 14909 2605 14943
rect 2605 14909 2639 14943
rect 2639 14909 2648 14943
rect 2596 14900 2648 14909
rect 4160 14968 4212 15020
rect 3424 14832 3476 14884
rect 1584 14764 1636 14816
rect 1952 14764 2004 14816
rect 3884 14832 3936 14884
rect 4068 14900 4120 14952
rect 4344 14900 4396 14952
rect 6460 15079 6512 15088
rect 6460 15045 6469 15079
rect 6469 15045 6503 15079
rect 6503 15045 6512 15079
rect 6460 15036 6512 15045
rect 4896 14968 4948 15020
rect 4804 14900 4856 14952
rect 5540 14900 5592 14952
rect 4436 14832 4488 14884
rect 4712 14875 4764 14884
rect 4712 14841 4721 14875
rect 4721 14841 4755 14875
rect 4755 14841 4764 14875
rect 4712 14832 4764 14841
rect 4896 14832 4948 14884
rect 5172 14832 5224 14884
rect 6184 14943 6236 14952
rect 6184 14909 6193 14943
rect 6193 14909 6227 14943
rect 6227 14909 6236 14943
rect 6184 14900 6236 14909
rect 3700 14807 3752 14816
rect 3700 14773 3709 14807
rect 3709 14773 3743 14807
rect 3743 14773 3752 14807
rect 3700 14764 3752 14773
rect 3792 14764 3844 14816
rect 6276 14832 6328 14884
rect 6920 14943 6972 14952
rect 6920 14909 6929 14943
rect 6929 14909 6963 14943
rect 6963 14909 6972 14943
rect 6920 14900 6972 14909
rect 7840 14900 7892 14952
rect 8484 15104 8536 15156
rect 9220 15104 9272 15156
rect 10324 15147 10376 15156
rect 10324 15113 10333 15147
rect 10333 15113 10367 15147
rect 10367 15113 10376 15147
rect 10324 15104 10376 15113
rect 10232 15036 10284 15088
rect 12164 15104 12216 15156
rect 12440 15104 12492 15156
rect 12624 15104 12676 15156
rect 15292 15104 15344 15156
rect 12716 15036 12768 15088
rect 12900 15036 12952 15088
rect 13268 15036 13320 15088
rect 13728 15036 13780 15088
rect 9312 15011 9364 15020
rect 9312 14977 9321 15011
rect 9321 14977 9355 15011
rect 9355 14977 9364 15011
rect 9312 14968 9364 14977
rect 7472 14832 7524 14884
rect 5908 14764 5960 14816
rect 6920 14764 6972 14816
rect 7012 14764 7064 14816
rect 7932 14764 7984 14816
rect 9128 14832 9180 14884
rect 10140 14900 10192 14952
rect 10692 14968 10744 15020
rect 11796 15011 11848 15020
rect 11796 14977 11805 15011
rect 11805 14977 11839 15011
rect 11839 14977 11848 15011
rect 11796 14968 11848 14977
rect 10600 14943 10652 14952
rect 10600 14909 10609 14943
rect 10609 14909 10643 14943
rect 10643 14909 10652 14943
rect 10600 14900 10652 14909
rect 10968 14900 11020 14952
rect 11060 14943 11112 14952
rect 11060 14909 11069 14943
rect 11069 14909 11103 14943
rect 11103 14909 11112 14943
rect 11060 14900 11112 14909
rect 12072 14943 12124 14952
rect 12072 14909 12081 14943
rect 12081 14909 12115 14943
rect 12115 14909 12124 14943
rect 12072 14900 12124 14909
rect 8760 14807 8812 14816
rect 8760 14773 8769 14807
rect 8769 14773 8803 14807
rect 8803 14773 8812 14807
rect 8760 14764 8812 14773
rect 9036 14764 9088 14816
rect 10416 14764 10468 14816
rect 10968 14764 11020 14816
rect 13820 14968 13872 15020
rect 15016 15011 15068 15020
rect 12900 14900 12952 14952
rect 12992 14943 13044 14952
rect 12992 14909 13001 14943
rect 13001 14909 13035 14943
rect 13035 14909 13044 14943
rect 12992 14900 13044 14909
rect 12808 14764 12860 14816
rect 12900 14807 12952 14816
rect 12900 14773 12909 14807
rect 12909 14773 12943 14807
rect 12943 14773 12952 14807
rect 12900 14764 12952 14773
rect 13268 14807 13320 14816
rect 13268 14773 13277 14807
rect 13277 14773 13311 14807
rect 13311 14773 13320 14807
rect 13268 14764 13320 14773
rect 14004 14943 14056 14952
rect 14004 14909 14013 14943
rect 14013 14909 14047 14943
rect 14047 14909 14056 14943
rect 14004 14900 14056 14909
rect 14372 14900 14424 14952
rect 13728 14875 13780 14884
rect 13728 14841 13737 14875
rect 13737 14841 13771 14875
rect 13771 14841 13780 14875
rect 13728 14832 13780 14841
rect 13912 14875 13964 14884
rect 13912 14841 13921 14875
rect 13921 14841 13955 14875
rect 13955 14841 13964 14875
rect 15016 14977 15025 15011
rect 15025 14977 15059 15011
rect 15059 14977 15068 15011
rect 15016 14968 15068 14977
rect 14832 14900 14884 14952
rect 15108 14943 15160 14952
rect 15108 14909 15117 14943
rect 15117 14909 15151 14943
rect 15151 14909 15160 14943
rect 15108 14900 15160 14909
rect 20720 15104 20772 15156
rect 16488 15036 16540 15088
rect 17684 14968 17736 15020
rect 18696 14968 18748 15020
rect 18972 15011 19024 15020
rect 18972 14977 18981 15011
rect 18981 14977 19015 15011
rect 19015 14977 19024 15011
rect 18972 14968 19024 14977
rect 19156 15011 19208 15020
rect 19156 14977 19165 15011
rect 19165 14977 19199 15011
rect 19199 14977 19208 15011
rect 19156 14968 19208 14977
rect 19340 15079 19392 15088
rect 19340 15045 19349 15079
rect 19349 15045 19383 15079
rect 19383 15045 19392 15079
rect 19340 15036 19392 15045
rect 19800 15036 19852 15088
rect 19984 15036 20036 15088
rect 17132 14943 17184 14952
rect 17132 14909 17141 14943
rect 17141 14909 17175 14943
rect 17175 14909 17184 14943
rect 17132 14900 17184 14909
rect 18144 14900 18196 14952
rect 19248 14900 19300 14952
rect 19524 14943 19576 14952
rect 19524 14909 19533 14943
rect 19533 14909 19567 14943
rect 19567 14909 19576 14943
rect 19524 14900 19576 14909
rect 13912 14832 13964 14841
rect 19340 14832 19392 14884
rect 20812 14900 20864 14952
rect 19800 14832 19852 14884
rect 14096 14764 14148 14816
rect 14188 14807 14240 14816
rect 14188 14773 14197 14807
rect 14197 14773 14231 14807
rect 14231 14773 14240 14807
rect 14188 14764 14240 14773
rect 14556 14764 14608 14816
rect 15108 14764 15160 14816
rect 16212 14807 16264 14816
rect 16212 14773 16221 14807
rect 16221 14773 16255 14807
rect 16255 14773 16264 14807
rect 16212 14764 16264 14773
rect 16304 14764 16356 14816
rect 17408 14764 17460 14816
rect 18696 14807 18748 14816
rect 18696 14773 18705 14807
rect 18705 14773 18739 14807
rect 18739 14773 18748 14807
rect 18696 14764 18748 14773
rect 19524 14764 19576 14816
rect 19984 14764 20036 14816
rect 20352 14764 20404 14816
rect 20444 14764 20496 14816
rect 22560 15011 22612 15020
rect 22560 14977 22569 15011
rect 22569 14977 22603 15011
rect 22603 14977 22612 15011
rect 22560 14968 22612 14977
rect 22284 14900 22336 14952
rect 22468 14943 22520 14952
rect 22468 14909 22477 14943
rect 22477 14909 22511 14943
rect 22511 14909 22520 14943
rect 22468 14900 22520 14909
rect 21364 14764 21416 14816
rect 21824 14764 21876 14816
rect 4366 14662 4418 14714
rect 4430 14662 4482 14714
rect 4494 14662 4546 14714
rect 4558 14662 4610 14714
rect 4622 14662 4674 14714
rect 4686 14662 4738 14714
rect 10366 14662 10418 14714
rect 10430 14662 10482 14714
rect 10494 14662 10546 14714
rect 10558 14662 10610 14714
rect 10622 14662 10674 14714
rect 10686 14662 10738 14714
rect 16366 14662 16418 14714
rect 16430 14662 16482 14714
rect 16494 14662 16546 14714
rect 16558 14662 16610 14714
rect 16622 14662 16674 14714
rect 16686 14662 16738 14714
rect 22366 14662 22418 14714
rect 22430 14662 22482 14714
rect 22494 14662 22546 14714
rect 22558 14662 22610 14714
rect 22622 14662 22674 14714
rect 22686 14662 22738 14714
rect 1860 14560 1912 14612
rect 3424 14603 3476 14612
rect 3424 14569 3433 14603
rect 3433 14569 3467 14603
rect 3467 14569 3476 14603
rect 3424 14560 3476 14569
rect 4068 14560 4120 14612
rect 4252 14603 4304 14612
rect 4252 14569 4261 14603
rect 4261 14569 4295 14603
rect 4295 14569 4304 14603
rect 4252 14560 4304 14569
rect 4896 14560 4948 14612
rect 6184 14560 6236 14612
rect 6552 14560 6604 14612
rect 8392 14560 8444 14612
rect 1768 14535 1820 14544
rect 1768 14501 1777 14535
rect 1777 14501 1811 14535
rect 1811 14501 1820 14535
rect 1768 14492 1820 14501
rect 1032 14467 1084 14476
rect 1032 14433 1041 14467
rect 1041 14433 1075 14467
rect 1075 14433 1084 14467
rect 1032 14424 1084 14433
rect 1124 14467 1176 14476
rect 1124 14433 1133 14467
rect 1133 14433 1167 14467
rect 1167 14433 1176 14467
rect 1124 14424 1176 14433
rect 1584 14467 1636 14476
rect 1584 14433 1593 14467
rect 1593 14433 1627 14467
rect 1627 14433 1636 14467
rect 1584 14424 1636 14433
rect 2044 14467 2096 14476
rect 2044 14433 2053 14467
rect 2053 14433 2087 14467
rect 2087 14433 2096 14467
rect 2044 14424 2096 14433
rect 2596 14492 2648 14544
rect 3700 14492 3752 14544
rect 4804 14492 4856 14544
rect 5448 14492 5500 14544
rect 6736 14492 6788 14544
rect 2964 14467 3016 14476
rect 2964 14433 2973 14467
rect 2973 14433 3007 14467
rect 3007 14433 3016 14467
rect 2964 14424 3016 14433
rect 3148 14424 3200 14476
rect 3884 14424 3936 14476
rect 4528 14467 4580 14476
rect 4528 14433 4537 14467
rect 4537 14433 4571 14467
rect 4571 14433 4580 14467
rect 4528 14424 4580 14433
rect 4620 14467 4672 14476
rect 4620 14433 4629 14467
rect 4629 14433 4663 14467
rect 4663 14433 4672 14467
rect 4620 14424 4672 14433
rect 5172 14424 5224 14476
rect 6092 14467 6144 14476
rect 6092 14433 6101 14467
rect 6101 14433 6135 14467
rect 6135 14433 6144 14467
rect 6092 14424 6144 14433
rect 7104 14424 7156 14476
rect 7932 14535 7984 14544
rect 7932 14501 7941 14535
rect 7941 14501 7975 14535
rect 7975 14501 7984 14535
rect 7932 14492 7984 14501
rect 9220 14560 9272 14612
rect 10048 14560 10100 14612
rect 11060 14560 11112 14612
rect 12256 14603 12308 14612
rect 12256 14569 12265 14603
rect 12265 14569 12299 14603
rect 12299 14569 12308 14603
rect 12256 14560 12308 14569
rect 7472 14467 7524 14476
rect 7472 14433 7481 14467
rect 7481 14433 7515 14467
rect 7515 14433 7524 14467
rect 7472 14424 7524 14433
rect 8208 14424 8260 14476
rect 8484 14424 8536 14476
rect 9312 14492 9364 14544
rect 8760 14424 8812 14476
rect 8852 14467 8904 14476
rect 8852 14433 8861 14467
rect 8861 14433 8895 14467
rect 8895 14433 8904 14467
rect 8852 14424 8904 14433
rect 9220 14467 9272 14476
rect 9220 14433 9229 14467
rect 9229 14433 9263 14467
rect 9263 14433 9272 14467
rect 9220 14424 9272 14433
rect 9404 14467 9456 14476
rect 9404 14433 9413 14467
rect 9413 14433 9447 14467
rect 9447 14433 9456 14467
rect 9404 14424 9456 14433
rect 9588 14467 9640 14476
rect 9588 14433 9597 14467
rect 9597 14433 9631 14467
rect 9631 14433 9640 14467
rect 9588 14424 9640 14433
rect 9680 14467 9732 14476
rect 9680 14433 9689 14467
rect 9689 14433 9723 14467
rect 9723 14433 9732 14467
rect 9680 14424 9732 14433
rect 10048 14424 10100 14476
rect 10600 14492 10652 14544
rect 12808 14560 12860 14612
rect 13176 14560 13228 14612
rect 13636 14560 13688 14612
rect 17316 14560 17368 14612
rect 17684 14603 17736 14612
rect 17684 14569 17693 14603
rect 17693 14569 17727 14603
rect 17727 14569 17736 14603
rect 17684 14560 17736 14569
rect 19248 14560 19300 14612
rect 21272 14560 21324 14612
rect 12716 14492 12768 14544
rect 14740 14492 14792 14544
rect 18696 14492 18748 14544
rect 21364 14535 21416 14544
rect 21364 14501 21373 14535
rect 21373 14501 21407 14535
rect 21407 14501 21416 14535
rect 21364 14492 21416 14501
rect 10968 14424 11020 14476
rect 11704 14424 11756 14476
rect 11796 14467 11848 14476
rect 11796 14433 11805 14467
rect 11805 14433 11839 14467
rect 11839 14433 11848 14467
rect 11796 14424 11848 14433
rect 12348 14424 12400 14476
rect 12624 14424 12676 14476
rect 12808 14467 12860 14476
rect 12808 14433 12817 14467
rect 12817 14433 12851 14467
rect 12851 14433 12860 14467
rect 12808 14424 12860 14433
rect 2412 14399 2464 14408
rect 2412 14365 2421 14399
rect 2421 14365 2455 14399
rect 2455 14365 2464 14399
rect 2412 14356 2464 14365
rect 2872 14399 2924 14408
rect 2872 14365 2881 14399
rect 2881 14365 2915 14399
rect 2915 14365 2924 14399
rect 2872 14356 2924 14365
rect 3516 14288 3568 14340
rect 9956 14356 10008 14408
rect 10416 14356 10468 14408
rect 11612 14356 11664 14408
rect 12072 14399 12124 14408
rect 12072 14365 12081 14399
rect 12081 14365 12115 14399
rect 12115 14365 12124 14399
rect 12072 14356 12124 14365
rect 12440 14356 12492 14408
rect 13268 14424 13320 14476
rect 14004 14467 14056 14476
rect 14004 14433 14013 14467
rect 14013 14433 14047 14467
rect 14047 14433 14056 14467
rect 14004 14424 14056 14433
rect 14188 14424 14240 14476
rect 15016 14424 15068 14476
rect 13176 14356 13228 14408
rect 10140 14288 10192 14340
rect 10324 14288 10376 14340
rect 14372 14399 14424 14408
rect 14372 14365 14381 14399
rect 14381 14365 14415 14399
rect 14415 14365 14424 14399
rect 14372 14356 14424 14365
rect 14924 14356 14976 14408
rect 1860 14263 1912 14272
rect 1860 14229 1869 14263
rect 1869 14229 1903 14263
rect 1903 14229 1912 14263
rect 1860 14220 1912 14229
rect 3148 14220 3200 14272
rect 5540 14263 5592 14272
rect 5540 14229 5549 14263
rect 5549 14229 5583 14263
rect 5583 14229 5592 14263
rect 5540 14220 5592 14229
rect 7012 14220 7064 14272
rect 8392 14220 8444 14272
rect 9772 14220 9824 14272
rect 9956 14220 10008 14272
rect 10508 14220 10560 14272
rect 10784 14220 10836 14272
rect 11060 14220 11112 14272
rect 11336 14220 11388 14272
rect 12624 14263 12676 14272
rect 12624 14229 12633 14263
rect 12633 14229 12667 14263
rect 12667 14229 12676 14263
rect 12624 14220 12676 14229
rect 16764 14288 16816 14340
rect 17132 14288 17184 14340
rect 17684 14467 17736 14476
rect 17684 14433 17693 14467
rect 17693 14433 17727 14467
rect 17727 14433 17736 14467
rect 17684 14424 17736 14433
rect 18420 14424 18472 14476
rect 18972 14424 19024 14476
rect 18696 14356 18748 14408
rect 19984 14424 20036 14476
rect 19340 14399 19392 14408
rect 19340 14365 19349 14399
rect 19349 14365 19383 14399
rect 19383 14365 19392 14399
rect 19340 14356 19392 14365
rect 19892 14356 19944 14408
rect 20352 14467 20404 14476
rect 20352 14433 20361 14467
rect 20361 14433 20395 14467
rect 20395 14433 20404 14467
rect 20352 14424 20404 14433
rect 20444 14467 20496 14476
rect 20444 14433 20453 14467
rect 20453 14433 20487 14467
rect 20487 14433 20496 14467
rect 20444 14424 20496 14433
rect 21180 14424 21232 14476
rect 21916 14424 21968 14476
rect 22008 14467 22060 14476
rect 22008 14433 22017 14467
rect 22017 14433 22051 14467
rect 22051 14433 22060 14467
rect 22008 14424 22060 14433
rect 22284 14467 22336 14476
rect 22284 14433 22293 14467
rect 22293 14433 22327 14467
rect 22327 14433 22336 14467
rect 22284 14424 22336 14433
rect 19248 14288 19300 14340
rect 14556 14220 14608 14272
rect 14832 14220 14884 14272
rect 15108 14220 15160 14272
rect 15844 14220 15896 14272
rect 19524 14220 19576 14272
rect 20444 14220 20496 14272
rect 21640 14220 21692 14272
rect 22468 14220 22520 14272
rect 1366 14118 1418 14170
rect 1430 14118 1482 14170
rect 1494 14118 1546 14170
rect 1558 14118 1610 14170
rect 1622 14118 1674 14170
rect 1686 14118 1738 14170
rect 7366 14118 7418 14170
rect 7430 14118 7482 14170
rect 7494 14118 7546 14170
rect 7558 14118 7610 14170
rect 7622 14118 7674 14170
rect 7686 14118 7738 14170
rect 13366 14118 13418 14170
rect 13430 14118 13482 14170
rect 13494 14118 13546 14170
rect 13558 14118 13610 14170
rect 13622 14118 13674 14170
rect 13686 14118 13738 14170
rect 19366 14118 19418 14170
rect 19430 14118 19482 14170
rect 19494 14118 19546 14170
rect 19558 14118 19610 14170
rect 19622 14118 19674 14170
rect 19686 14118 19738 14170
rect 2964 14059 3016 14068
rect 2964 14025 2973 14059
rect 2973 14025 3007 14059
rect 3007 14025 3016 14059
rect 2964 14016 3016 14025
rect 4068 14016 4120 14068
rect 6828 14016 6880 14068
rect 9772 14016 9824 14068
rect 10416 14016 10468 14068
rect 12348 14016 12400 14068
rect 12808 14016 12860 14068
rect 13360 14016 13412 14068
rect 14372 14016 14424 14068
rect 15476 14016 15528 14068
rect 2688 13948 2740 14000
rect 4528 13948 4580 14000
rect 5080 13948 5132 14000
rect 8116 13991 8168 14000
rect 8116 13957 8125 13991
rect 8125 13957 8159 13991
rect 8159 13957 8168 13991
rect 8116 13948 8168 13957
rect 10692 13948 10744 14000
rect 11244 13948 11296 14000
rect 11796 13948 11848 14000
rect 3056 13923 3108 13932
rect 3056 13889 3065 13923
rect 3065 13889 3099 13923
rect 3099 13889 3108 13923
rect 3056 13880 3108 13889
rect 848 13855 900 13864
rect 848 13821 857 13855
rect 857 13821 891 13855
rect 891 13821 900 13855
rect 848 13812 900 13821
rect 1124 13812 1176 13864
rect 1216 13812 1268 13864
rect 1860 13812 1912 13864
rect 1032 13787 1084 13796
rect 1032 13753 1041 13787
rect 1041 13753 1075 13787
rect 1075 13753 1084 13787
rect 1032 13744 1084 13753
rect 2412 13744 2464 13796
rect 3608 13812 3660 13864
rect 3976 13812 4028 13864
rect 5080 13812 5132 13864
rect 7380 13812 7432 13864
rect 7656 13812 7708 13864
rect 8760 13880 8812 13932
rect 8944 13855 8996 13864
rect 8944 13821 8953 13855
rect 8953 13821 8987 13855
rect 8987 13821 8996 13855
rect 8944 13812 8996 13821
rect 9404 13812 9456 13864
rect 7564 13787 7616 13796
rect 7564 13753 7573 13787
rect 7573 13753 7607 13787
rect 7607 13753 7616 13787
rect 7564 13744 7616 13753
rect 9312 13787 9364 13796
rect 9312 13753 9321 13787
rect 9321 13753 9355 13787
rect 9355 13753 9364 13787
rect 9312 13744 9364 13753
rect 9772 13744 9824 13796
rect 10232 13812 10284 13864
rect 10600 13744 10652 13796
rect 11336 13744 11388 13796
rect 11704 13812 11756 13864
rect 12992 13880 13044 13932
rect 12808 13812 12860 13864
rect 13268 13812 13320 13864
rect 13820 13855 13872 13864
rect 13820 13821 13829 13855
rect 13829 13821 13863 13855
rect 13863 13821 13872 13855
rect 13820 13812 13872 13821
rect 13912 13812 13964 13864
rect 14740 13812 14792 13864
rect 15108 13812 15160 13864
rect 16120 13880 16172 13932
rect 16396 13880 16448 13932
rect 15292 13855 15344 13864
rect 15292 13821 15301 13855
rect 15301 13821 15335 13855
rect 15335 13821 15344 13855
rect 15292 13812 15344 13821
rect 15476 13855 15528 13864
rect 15476 13821 15485 13855
rect 15485 13821 15519 13855
rect 15519 13821 15528 13855
rect 15476 13812 15528 13821
rect 15936 13812 15988 13864
rect 12072 13744 12124 13796
rect 1308 13676 1360 13728
rect 2596 13676 2648 13728
rect 3884 13676 3936 13728
rect 7472 13676 7524 13728
rect 8300 13676 8352 13728
rect 8668 13676 8720 13728
rect 9220 13676 9272 13728
rect 10048 13676 10100 13728
rect 10232 13676 10284 13728
rect 10324 13719 10376 13728
rect 10324 13685 10333 13719
rect 10333 13685 10367 13719
rect 10367 13685 10376 13719
rect 10324 13676 10376 13685
rect 10508 13676 10560 13728
rect 11704 13676 11756 13728
rect 12256 13676 12308 13728
rect 16212 13855 16264 13864
rect 16212 13821 16221 13855
rect 16221 13821 16255 13855
rect 16255 13821 16264 13855
rect 16212 13812 16264 13821
rect 16948 13948 17000 14000
rect 16856 13812 16908 13864
rect 17132 13880 17184 13932
rect 19340 14016 19392 14068
rect 21640 14016 21692 14068
rect 17776 13880 17828 13932
rect 19616 13948 19668 14000
rect 18236 13855 18288 13864
rect 18236 13821 18245 13855
rect 18245 13821 18279 13855
rect 18279 13821 18288 13855
rect 18236 13812 18288 13821
rect 18420 13787 18472 13796
rect 18420 13753 18429 13787
rect 18429 13753 18463 13787
rect 18463 13753 18472 13787
rect 18420 13744 18472 13753
rect 18788 13812 18840 13864
rect 19340 13855 19392 13864
rect 19340 13821 19349 13855
rect 19349 13821 19383 13855
rect 19383 13821 19392 13855
rect 19340 13812 19392 13821
rect 19708 13880 19760 13932
rect 19984 13880 20036 13932
rect 20352 13948 20404 14000
rect 20260 13923 20312 13932
rect 20260 13889 20269 13923
rect 20269 13889 20303 13923
rect 20303 13889 20312 13923
rect 20812 13948 20864 14000
rect 20260 13880 20312 13889
rect 20536 13812 20588 13864
rect 21640 13855 21692 13864
rect 21640 13821 21649 13855
rect 21649 13821 21683 13855
rect 21683 13821 21692 13855
rect 21640 13812 21692 13821
rect 22468 13855 22520 13864
rect 22468 13821 22477 13855
rect 22477 13821 22511 13855
rect 22511 13821 22520 13855
rect 22468 13812 22520 13821
rect 14556 13676 14608 13728
rect 15108 13719 15160 13728
rect 15108 13685 15117 13719
rect 15117 13685 15151 13719
rect 15151 13685 15160 13719
rect 15108 13676 15160 13685
rect 16212 13719 16264 13728
rect 16212 13685 16221 13719
rect 16221 13685 16255 13719
rect 16255 13685 16264 13719
rect 16212 13676 16264 13685
rect 16396 13676 16448 13728
rect 16764 13676 16816 13728
rect 17684 13676 17736 13728
rect 18696 13719 18748 13728
rect 18696 13685 18705 13719
rect 18705 13685 18739 13719
rect 18739 13685 18748 13719
rect 18696 13676 18748 13685
rect 19800 13676 19852 13728
rect 19984 13719 20036 13728
rect 19984 13685 19993 13719
rect 19993 13685 20027 13719
rect 20027 13685 20036 13719
rect 19984 13676 20036 13685
rect 20536 13676 20588 13728
rect 21180 13676 21232 13728
rect 4366 13574 4418 13626
rect 4430 13574 4482 13626
rect 4494 13574 4546 13626
rect 4558 13574 4610 13626
rect 4622 13574 4674 13626
rect 4686 13574 4738 13626
rect 10366 13574 10418 13626
rect 10430 13574 10482 13626
rect 10494 13574 10546 13626
rect 10558 13574 10610 13626
rect 10622 13574 10674 13626
rect 10686 13574 10738 13626
rect 16366 13574 16418 13626
rect 16430 13574 16482 13626
rect 16494 13574 16546 13626
rect 16558 13574 16610 13626
rect 16622 13574 16674 13626
rect 16686 13574 16738 13626
rect 22366 13574 22418 13626
rect 22430 13574 22482 13626
rect 22494 13574 22546 13626
rect 22558 13574 22610 13626
rect 22622 13574 22674 13626
rect 22686 13574 22738 13626
rect 1308 13472 1360 13524
rect 2044 13515 2096 13524
rect 2044 13481 2053 13515
rect 2053 13481 2087 13515
rect 2087 13481 2096 13515
rect 2044 13472 2096 13481
rect 2596 13472 2648 13524
rect 1124 13404 1176 13456
rect 3056 13404 3108 13456
rect 848 13379 900 13388
rect 848 13345 857 13379
rect 857 13345 891 13379
rect 891 13345 900 13379
rect 848 13336 900 13345
rect 1768 13336 1820 13388
rect 2412 13336 2464 13388
rect 6184 13472 6236 13524
rect 7564 13472 7616 13524
rect 7840 13472 7892 13524
rect 8024 13472 8076 13524
rect 8668 13515 8720 13524
rect 8668 13481 8677 13515
rect 8677 13481 8711 13515
rect 8711 13481 8720 13515
rect 8668 13472 8720 13481
rect 9680 13472 9732 13524
rect 10232 13472 10284 13524
rect 4620 13404 4672 13456
rect 5356 13404 5408 13456
rect 5540 13404 5592 13456
rect 6920 13404 6972 13456
rect 7104 13404 7156 13456
rect 7472 13404 7524 13456
rect 9312 13404 9364 13456
rect 2504 13268 2556 13320
rect 3608 13379 3660 13388
rect 3608 13345 3617 13379
rect 3617 13345 3651 13379
rect 3651 13345 3660 13379
rect 3608 13336 3660 13345
rect 4252 13379 4304 13388
rect 4252 13345 4261 13379
rect 4261 13345 4295 13379
rect 4295 13345 4304 13379
rect 4252 13336 4304 13345
rect 4988 13336 5040 13388
rect 2688 13311 2740 13320
rect 2688 13277 2697 13311
rect 2697 13277 2731 13311
rect 2731 13277 2740 13311
rect 2688 13268 2740 13277
rect 1768 13132 1820 13184
rect 2136 13132 2188 13184
rect 4160 13311 4212 13320
rect 4160 13277 4169 13311
rect 4169 13277 4203 13311
rect 4203 13277 4212 13311
rect 4160 13268 4212 13277
rect 7656 13268 7708 13320
rect 8300 13336 8352 13388
rect 9220 13379 9272 13388
rect 9220 13345 9229 13379
rect 9229 13345 9263 13379
rect 9263 13345 9272 13379
rect 9220 13336 9272 13345
rect 9036 13268 9088 13320
rect 9496 13379 9548 13388
rect 9496 13345 9505 13379
rect 9505 13345 9539 13379
rect 9539 13345 9548 13379
rect 9496 13336 9548 13345
rect 10140 13404 10192 13456
rect 9680 13336 9732 13388
rect 11336 13472 11388 13524
rect 10508 13379 10560 13388
rect 10508 13345 10517 13379
rect 10517 13345 10551 13379
rect 10551 13345 10560 13379
rect 10508 13336 10560 13345
rect 11704 13404 11756 13456
rect 11796 13447 11848 13456
rect 11796 13413 11805 13447
rect 11805 13413 11839 13447
rect 11839 13413 11848 13447
rect 11796 13404 11848 13413
rect 12348 13404 12400 13456
rect 11060 13336 11112 13388
rect 11244 13379 11296 13388
rect 11244 13345 11253 13379
rect 11253 13345 11287 13379
rect 11287 13345 11296 13379
rect 11244 13336 11296 13345
rect 5356 13200 5408 13252
rect 6184 13200 6236 13252
rect 9772 13200 9824 13252
rect 10968 13268 11020 13320
rect 12256 13336 12308 13388
rect 12716 13336 12768 13388
rect 14096 13404 14148 13456
rect 15292 13404 15344 13456
rect 15108 13379 15160 13388
rect 15108 13345 15117 13379
rect 15117 13345 15151 13379
rect 15151 13345 15160 13379
rect 15108 13336 15160 13345
rect 16580 13472 16632 13524
rect 17040 13472 17092 13524
rect 19708 13472 19760 13524
rect 18604 13404 18656 13456
rect 19892 13404 19944 13456
rect 17040 13336 17092 13388
rect 17500 13379 17552 13388
rect 17500 13345 17509 13379
rect 17509 13345 17543 13379
rect 17543 13345 17552 13379
rect 17500 13336 17552 13345
rect 17684 13379 17736 13388
rect 17684 13345 17693 13379
rect 17693 13345 17727 13379
rect 17727 13345 17736 13379
rect 17684 13336 17736 13345
rect 17776 13336 17828 13388
rect 19616 13379 19668 13388
rect 19616 13345 19625 13379
rect 19625 13345 19659 13379
rect 19659 13345 19668 13379
rect 19616 13336 19668 13345
rect 20536 13336 20588 13388
rect 12808 13311 12860 13320
rect 12808 13277 12817 13311
rect 12817 13277 12851 13311
rect 12851 13277 12860 13311
rect 12808 13268 12860 13277
rect 13360 13268 13412 13320
rect 14740 13268 14792 13320
rect 15200 13268 15252 13320
rect 16672 13268 16724 13320
rect 12256 13200 12308 13252
rect 3976 13132 4028 13184
rect 5448 13132 5500 13184
rect 10140 13175 10192 13184
rect 10140 13141 10149 13175
rect 10149 13141 10183 13175
rect 10183 13141 10192 13175
rect 10140 13132 10192 13141
rect 11612 13132 11664 13184
rect 13728 13200 13780 13252
rect 15108 13200 15160 13252
rect 18604 13268 18656 13320
rect 18420 13200 18472 13252
rect 20812 13200 20864 13252
rect 12992 13132 13044 13184
rect 14188 13175 14240 13184
rect 14188 13141 14197 13175
rect 14197 13141 14231 13175
rect 14231 13141 14240 13175
rect 14188 13132 14240 13141
rect 14924 13132 14976 13184
rect 15200 13132 15252 13184
rect 17132 13132 17184 13184
rect 17592 13132 17644 13184
rect 18880 13132 18932 13184
rect 20076 13132 20128 13184
rect 20260 13132 20312 13184
rect 20720 13132 20772 13184
rect 21088 13132 21140 13184
rect 1366 13030 1418 13082
rect 1430 13030 1482 13082
rect 1494 13030 1546 13082
rect 1558 13030 1610 13082
rect 1622 13030 1674 13082
rect 1686 13030 1738 13082
rect 7366 13030 7418 13082
rect 7430 13030 7482 13082
rect 7494 13030 7546 13082
rect 7558 13030 7610 13082
rect 7622 13030 7674 13082
rect 7686 13030 7738 13082
rect 13366 13030 13418 13082
rect 13430 13030 13482 13082
rect 13494 13030 13546 13082
rect 13558 13030 13610 13082
rect 13622 13030 13674 13082
rect 13686 13030 13738 13082
rect 19366 13030 19418 13082
rect 19430 13030 19482 13082
rect 19494 13030 19546 13082
rect 19558 13030 19610 13082
rect 19622 13030 19674 13082
rect 19686 13030 19738 13082
rect 848 12928 900 12980
rect 756 12860 808 12912
rect 1676 12903 1728 12912
rect 1676 12869 1685 12903
rect 1685 12869 1719 12903
rect 1719 12869 1728 12903
rect 1676 12860 1728 12869
rect 2320 12860 2372 12912
rect 664 12792 716 12844
rect 5080 12928 5132 12980
rect 7196 12928 7248 12980
rect 6276 12860 6328 12912
rect 8760 12928 8812 12980
rect 9220 12928 9272 12980
rect 10968 12971 11020 12980
rect 10968 12937 10977 12971
rect 10977 12937 11011 12971
rect 11011 12937 11020 12971
rect 10968 12928 11020 12937
rect 7840 12860 7892 12912
rect 10048 12860 10100 12912
rect 10508 12860 10560 12912
rect 6828 12792 6880 12844
rect 6920 12792 6972 12844
rect 11980 12928 12032 12980
rect 1032 12724 1084 12776
rect 2044 12724 2096 12776
rect 2964 12724 3016 12776
rect 1492 12656 1544 12708
rect 2228 12656 2280 12708
rect 2320 12699 2372 12708
rect 2320 12665 2329 12699
rect 2329 12665 2363 12699
rect 2363 12665 2372 12699
rect 2320 12656 2372 12665
rect 3332 12656 3384 12708
rect 3884 12767 3936 12776
rect 3884 12733 3893 12767
rect 3893 12733 3927 12767
rect 3927 12733 3936 12767
rect 3884 12724 3936 12733
rect 4160 12767 4212 12776
rect 4160 12733 4169 12767
rect 4169 12733 4203 12767
rect 4203 12733 4212 12767
rect 4160 12724 4212 12733
rect 4620 12767 4672 12776
rect 4620 12733 4629 12767
rect 4629 12733 4663 12767
rect 4663 12733 4672 12767
rect 4620 12724 4672 12733
rect 4988 12724 5040 12776
rect 7196 12724 7248 12776
rect 7472 12724 7524 12776
rect 3976 12656 4028 12708
rect 4252 12656 4304 12708
rect 1952 12631 2004 12640
rect 1952 12597 1961 12631
rect 1961 12597 1995 12631
rect 1995 12597 2004 12631
rect 1952 12588 2004 12597
rect 2412 12631 2464 12640
rect 2412 12597 2421 12631
rect 2421 12597 2455 12631
rect 2455 12597 2464 12631
rect 2412 12588 2464 12597
rect 3608 12588 3660 12640
rect 4160 12588 4212 12640
rect 4896 12656 4948 12708
rect 4988 12588 5040 12640
rect 5080 12631 5132 12640
rect 5080 12597 5089 12631
rect 5089 12597 5123 12631
rect 5123 12597 5132 12631
rect 5080 12588 5132 12597
rect 5172 12588 5224 12640
rect 5540 12656 5592 12708
rect 6184 12699 6236 12708
rect 6184 12665 6193 12699
rect 6193 12665 6227 12699
rect 6227 12665 6236 12699
rect 6184 12656 6236 12665
rect 8668 12724 8720 12776
rect 6460 12588 6512 12640
rect 6736 12588 6788 12640
rect 8392 12656 8444 12708
rect 9680 12767 9732 12776
rect 9680 12733 9689 12767
rect 9689 12733 9723 12767
rect 9723 12733 9732 12767
rect 9680 12724 9732 12733
rect 10232 12724 10284 12776
rect 10508 12724 10560 12776
rect 11336 12792 11388 12844
rect 12624 12860 12676 12912
rect 14464 12860 14516 12912
rect 8300 12588 8352 12640
rect 8852 12588 8904 12640
rect 9772 12588 9824 12640
rect 12072 12767 12124 12776
rect 12072 12733 12081 12767
rect 12081 12733 12115 12767
rect 12115 12733 12124 12767
rect 12072 12724 12124 12733
rect 12348 12767 12400 12776
rect 12348 12733 12357 12767
rect 12357 12733 12391 12767
rect 12391 12733 12400 12767
rect 12348 12724 12400 12733
rect 15108 12860 15160 12912
rect 11428 12588 11480 12640
rect 12440 12588 12492 12640
rect 12808 12724 12860 12776
rect 15016 12792 15068 12844
rect 14188 12767 14240 12776
rect 14188 12733 14197 12767
rect 14197 12733 14231 12767
rect 14231 12733 14240 12767
rect 19892 12928 19944 12980
rect 17224 12860 17276 12912
rect 18512 12860 18564 12912
rect 14188 12724 14240 12733
rect 15384 12767 15436 12776
rect 15384 12733 15393 12767
rect 15393 12733 15427 12767
rect 15427 12733 15436 12767
rect 15384 12724 15436 12733
rect 15476 12724 15528 12776
rect 16856 12724 16908 12776
rect 16948 12767 17000 12776
rect 16948 12733 16957 12767
rect 16957 12733 16991 12767
rect 16991 12733 17000 12767
rect 16948 12724 17000 12733
rect 15200 12656 15252 12708
rect 15292 12699 15344 12708
rect 15292 12665 15301 12699
rect 15301 12665 15335 12699
rect 15335 12665 15344 12699
rect 15292 12656 15344 12665
rect 18788 12835 18840 12844
rect 18788 12801 18797 12835
rect 18797 12801 18831 12835
rect 18831 12801 18840 12835
rect 18788 12792 18840 12801
rect 19432 12792 19484 12844
rect 20444 12792 20496 12844
rect 20996 12792 21048 12844
rect 18880 12767 18932 12776
rect 18880 12733 18889 12767
rect 18889 12733 18923 12767
rect 18923 12733 18932 12767
rect 18880 12724 18932 12733
rect 19524 12767 19576 12776
rect 19524 12733 19526 12767
rect 19526 12733 19560 12767
rect 19560 12733 19576 12767
rect 19524 12724 19576 12733
rect 19892 12767 19944 12776
rect 19892 12733 19901 12767
rect 19901 12733 19935 12767
rect 19935 12733 19944 12767
rect 19892 12724 19944 12733
rect 20076 12767 20128 12776
rect 20076 12733 20085 12767
rect 20085 12733 20119 12767
rect 20119 12733 20128 12767
rect 20076 12724 20128 12733
rect 20812 12767 20864 12776
rect 20812 12733 20821 12767
rect 20821 12733 20855 12767
rect 20855 12733 20864 12767
rect 20812 12724 20864 12733
rect 14372 12588 14424 12640
rect 14464 12588 14516 12640
rect 16028 12588 16080 12640
rect 17132 12588 17184 12640
rect 17592 12631 17644 12640
rect 17592 12597 17601 12631
rect 17601 12597 17635 12631
rect 17635 12597 17644 12631
rect 17592 12588 17644 12597
rect 18788 12588 18840 12640
rect 19294 12588 19346 12640
rect 21272 12588 21324 12640
rect 21456 12656 21508 12708
rect 21732 12656 21784 12708
rect 21824 12588 21876 12640
rect 22100 12588 22152 12640
rect 4366 12486 4418 12538
rect 4430 12486 4482 12538
rect 4494 12486 4546 12538
rect 4558 12486 4610 12538
rect 4622 12486 4674 12538
rect 4686 12486 4738 12538
rect 10366 12486 10418 12538
rect 10430 12486 10482 12538
rect 10494 12486 10546 12538
rect 10558 12486 10610 12538
rect 10622 12486 10674 12538
rect 10686 12486 10738 12538
rect 16366 12486 16418 12538
rect 16430 12486 16482 12538
rect 16494 12486 16546 12538
rect 16558 12486 16610 12538
rect 16622 12486 16674 12538
rect 16686 12486 16738 12538
rect 22366 12486 22418 12538
rect 22430 12486 22482 12538
rect 22494 12486 22546 12538
rect 22558 12486 22610 12538
rect 22622 12486 22674 12538
rect 22686 12486 22738 12538
rect 1032 12384 1084 12436
rect 1952 12384 2004 12436
rect 2228 12384 2280 12436
rect 3700 12384 3752 12436
rect 1676 12316 1728 12368
rect 1216 12248 1268 12300
rect 2412 12316 2464 12368
rect 4068 12316 4120 12368
rect 3424 12248 3476 12300
rect 3608 12248 3660 12300
rect 3884 12248 3936 12300
rect 4160 12248 4212 12300
rect 4896 12384 4948 12436
rect 6276 12384 6328 12436
rect 7472 12384 7524 12436
rect 9680 12384 9732 12436
rect 11428 12384 11480 12436
rect 15200 12384 15252 12436
rect 15384 12384 15436 12436
rect 15752 12384 15804 12436
rect 16304 12384 16356 12436
rect 4344 12291 4396 12300
rect 4344 12257 4353 12291
rect 4353 12257 4387 12291
rect 4387 12257 4396 12291
rect 4344 12248 4396 12257
rect 848 12112 900 12164
rect 1032 12112 1084 12164
rect 2044 12112 2096 12164
rect 2228 12044 2280 12096
rect 2780 12044 2832 12096
rect 4160 12112 4212 12164
rect 4252 12112 4304 12164
rect 5080 12248 5132 12300
rect 5264 12112 5316 12164
rect 5908 12223 5960 12232
rect 5908 12189 5917 12223
rect 5917 12189 5951 12223
rect 5951 12189 5960 12223
rect 5908 12180 5960 12189
rect 6736 12291 6788 12300
rect 6736 12257 6745 12291
rect 6745 12257 6779 12291
rect 6779 12257 6788 12291
rect 6736 12248 6788 12257
rect 7012 12291 7064 12300
rect 7012 12257 7021 12291
rect 7021 12257 7055 12291
rect 7055 12257 7064 12291
rect 7012 12248 7064 12257
rect 5816 12112 5868 12164
rect 3792 12044 3844 12096
rect 3976 12087 4028 12096
rect 3976 12053 3985 12087
rect 3985 12053 4019 12087
rect 4019 12053 4028 12087
rect 3976 12044 4028 12053
rect 4068 12087 4120 12096
rect 4068 12053 4077 12087
rect 4077 12053 4111 12087
rect 4111 12053 4120 12087
rect 4068 12044 4120 12053
rect 7472 12291 7524 12300
rect 7472 12257 7481 12291
rect 7481 12257 7515 12291
rect 7515 12257 7524 12291
rect 7472 12248 7524 12257
rect 8484 12316 8536 12368
rect 8392 12291 8444 12300
rect 8392 12257 8401 12291
rect 8401 12257 8435 12291
rect 8435 12257 8444 12291
rect 8392 12248 8444 12257
rect 8576 12248 8628 12300
rect 7012 12112 7064 12164
rect 8852 12291 8904 12300
rect 8852 12257 8861 12291
rect 8861 12257 8895 12291
rect 8895 12257 8904 12291
rect 8852 12248 8904 12257
rect 11060 12316 11112 12368
rect 11612 12248 11664 12300
rect 12072 12316 12124 12368
rect 11796 12291 11848 12300
rect 11796 12257 11805 12291
rect 11805 12257 11839 12291
rect 11839 12257 11848 12291
rect 11796 12248 11848 12257
rect 9220 12180 9272 12232
rect 12256 12223 12308 12232
rect 12256 12189 12265 12223
rect 12265 12189 12299 12223
rect 12299 12189 12308 12223
rect 12256 12180 12308 12189
rect 12716 12316 12768 12368
rect 14096 12316 14148 12368
rect 14832 12316 14884 12368
rect 14464 12248 14516 12300
rect 15016 12248 15068 12300
rect 15292 12248 15344 12300
rect 15936 12316 15988 12368
rect 16488 12359 16540 12368
rect 16488 12325 16497 12359
rect 16497 12325 16531 12359
rect 16531 12325 16540 12359
rect 16488 12316 16540 12325
rect 13268 12223 13320 12232
rect 13268 12189 13277 12223
rect 13277 12189 13311 12223
rect 13311 12189 13320 12223
rect 13268 12180 13320 12189
rect 14096 12180 14148 12232
rect 14280 12180 14332 12232
rect 16304 12291 16356 12300
rect 16304 12257 16313 12291
rect 16313 12257 16347 12291
rect 16347 12257 16356 12291
rect 16304 12248 16356 12257
rect 16396 12291 16448 12300
rect 16396 12257 16405 12291
rect 16405 12257 16439 12291
rect 16439 12257 16448 12291
rect 16396 12248 16448 12257
rect 9036 12112 9088 12164
rect 10784 12112 10836 12164
rect 10876 12112 10928 12164
rect 12072 12112 12124 12164
rect 12624 12112 12676 12164
rect 6644 12044 6696 12096
rect 7104 12044 7156 12096
rect 8576 12087 8628 12096
rect 8576 12053 8585 12087
rect 8585 12053 8619 12087
rect 8619 12053 8628 12087
rect 8576 12044 8628 12053
rect 8760 12044 8812 12096
rect 8852 12044 8904 12096
rect 9772 12044 9824 12096
rect 11428 12044 11480 12096
rect 13820 12044 13872 12096
rect 14740 12044 14792 12096
rect 15016 12044 15068 12096
rect 15660 12112 15712 12164
rect 16856 12291 16908 12300
rect 16856 12257 16865 12291
rect 16865 12257 16899 12291
rect 16899 12257 16908 12291
rect 16856 12248 16908 12257
rect 17592 12384 17644 12436
rect 17776 12384 17828 12436
rect 18696 12384 18748 12436
rect 19892 12427 19944 12436
rect 19892 12393 19901 12427
rect 19901 12393 19935 12427
rect 19935 12393 19944 12427
rect 19892 12384 19944 12393
rect 20352 12384 20404 12436
rect 21456 12427 21508 12436
rect 21456 12393 21465 12427
rect 21465 12393 21499 12427
rect 21499 12393 21508 12427
rect 21456 12384 21508 12393
rect 17132 12291 17184 12300
rect 17132 12257 17141 12291
rect 17141 12257 17175 12291
rect 17175 12257 17184 12291
rect 17132 12248 17184 12257
rect 18052 12291 18104 12300
rect 18052 12257 18061 12291
rect 18061 12257 18095 12291
rect 18095 12257 18104 12291
rect 18052 12248 18104 12257
rect 18328 12291 18380 12300
rect 18328 12257 18337 12291
rect 18337 12257 18371 12291
rect 18371 12257 18380 12291
rect 18328 12248 18380 12257
rect 18696 12248 18748 12300
rect 19432 12291 19484 12300
rect 19432 12257 19441 12291
rect 19441 12257 19475 12291
rect 19475 12257 19484 12291
rect 19432 12248 19484 12257
rect 19524 12291 19576 12300
rect 19524 12257 19533 12291
rect 19533 12257 19567 12291
rect 19567 12257 19576 12291
rect 19524 12248 19576 12257
rect 19984 12248 20036 12300
rect 20168 12180 20220 12232
rect 20260 12223 20312 12232
rect 20260 12189 20269 12223
rect 20269 12189 20303 12223
rect 20303 12189 20312 12223
rect 21640 12316 21692 12368
rect 20812 12248 20864 12300
rect 21272 12291 21324 12300
rect 21272 12257 21281 12291
rect 21281 12257 21315 12291
rect 21315 12257 21324 12291
rect 21272 12248 21324 12257
rect 21732 12248 21784 12300
rect 20260 12180 20312 12189
rect 20444 12180 20496 12232
rect 19524 12112 19576 12164
rect 20628 12223 20680 12232
rect 20628 12189 20637 12223
rect 20637 12189 20671 12223
rect 20671 12189 20680 12223
rect 20628 12180 20680 12189
rect 21824 12112 21876 12164
rect 15476 12044 15528 12096
rect 16028 12044 16080 12096
rect 16396 12044 16448 12096
rect 17316 12044 17368 12096
rect 17776 12044 17828 12096
rect 18144 12044 18196 12096
rect 18788 12087 18840 12096
rect 18788 12053 18797 12087
rect 18797 12053 18831 12087
rect 18831 12053 18840 12087
rect 18788 12044 18840 12053
rect 18880 12044 18932 12096
rect 21456 12044 21508 12096
rect 21548 12044 21600 12096
rect 1366 11942 1418 11994
rect 1430 11942 1482 11994
rect 1494 11942 1546 11994
rect 1558 11942 1610 11994
rect 1622 11942 1674 11994
rect 1686 11942 1738 11994
rect 7366 11942 7418 11994
rect 7430 11942 7482 11994
rect 7494 11942 7546 11994
rect 7558 11942 7610 11994
rect 7622 11942 7674 11994
rect 7686 11942 7738 11994
rect 13366 11942 13418 11994
rect 13430 11942 13482 11994
rect 13494 11942 13546 11994
rect 13558 11942 13610 11994
rect 13622 11942 13674 11994
rect 13686 11942 13738 11994
rect 19366 11942 19418 11994
rect 19430 11942 19482 11994
rect 19494 11942 19546 11994
rect 19558 11942 19610 11994
rect 19622 11942 19674 11994
rect 19686 11942 19738 11994
rect 940 11772 992 11824
rect 1308 11772 1360 11824
rect 1124 11704 1176 11756
rect 1584 11747 1636 11756
rect 1584 11713 1593 11747
rect 1593 11713 1627 11747
rect 1627 11713 1636 11747
rect 1584 11704 1636 11713
rect 1676 11747 1728 11756
rect 1676 11713 1685 11747
rect 1685 11713 1719 11747
rect 1719 11713 1728 11747
rect 1676 11704 1728 11713
rect 756 11636 808 11688
rect 1952 11704 2004 11756
rect 848 11568 900 11620
rect 1124 11611 1176 11620
rect 940 11543 992 11552
rect 940 11509 949 11543
rect 949 11509 983 11543
rect 983 11509 992 11543
rect 940 11500 992 11509
rect 1124 11577 1151 11611
rect 1151 11577 1176 11611
rect 1124 11568 1176 11577
rect 1308 11611 1360 11620
rect 1308 11577 1317 11611
rect 1317 11577 1351 11611
rect 1351 11577 1360 11611
rect 1308 11568 1360 11577
rect 1768 11568 1820 11620
rect 2780 11679 2832 11688
rect 2780 11645 2789 11679
rect 2789 11645 2823 11679
rect 2823 11645 2832 11679
rect 2780 11636 2832 11645
rect 3424 11679 3476 11688
rect 3424 11645 3433 11679
rect 3433 11645 3467 11679
rect 3467 11645 3476 11679
rect 3424 11636 3476 11645
rect 1952 11500 2004 11552
rect 2688 11500 2740 11552
rect 5080 11883 5132 11892
rect 5080 11849 5089 11883
rect 5089 11849 5123 11883
rect 5123 11849 5132 11883
rect 5080 11840 5132 11849
rect 5356 11840 5408 11892
rect 9772 11840 9824 11892
rect 9864 11840 9916 11892
rect 8760 11772 8812 11824
rect 12164 11840 12216 11892
rect 14280 11840 14332 11892
rect 16304 11840 16356 11892
rect 16856 11883 16908 11892
rect 16856 11849 16865 11883
rect 16865 11849 16899 11883
rect 16899 11849 16908 11883
rect 16856 11840 16908 11849
rect 16948 11883 17000 11892
rect 16948 11849 16957 11883
rect 16957 11849 16991 11883
rect 16991 11849 17000 11883
rect 16948 11840 17000 11849
rect 17592 11883 17644 11892
rect 17592 11849 17601 11883
rect 17601 11849 17635 11883
rect 17635 11849 17644 11883
rect 17592 11840 17644 11849
rect 18788 11883 18840 11892
rect 18788 11849 18797 11883
rect 18797 11849 18831 11883
rect 18831 11849 18840 11883
rect 18788 11840 18840 11849
rect 19892 11840 19944 11892
rect 19984 11840 20036 11892
rect 20076 11883 20128 11892
rect 20076 11849 20085 11883
rect 20085 11849 20119 11883
rect 20119 11849 20128 11883
rect 20076 11840 20128 11849
rect 21732 11840 21784 11892
rect 3792 11704 3844 11756
rect 4252 11747 4304 11756
rect 4252 11713 4261 11747
rect 4261 11713 4295 11747
rect 4295 11713 4304 11747
rect 4252 11704 4304 11713
rect 4344 11704 4396 11756
rect 4988 11704 5040 11756
rect 3608 11568 3660 11620
rect 4896 11636 4948 11688
rect 6092 11636 6144 11688
rect 7288 11636 7340 11688
rect 5356 11568 5408 11620
rect 8852 11704 8904 11756
rect 8484 11636 8536 11688
rect 8760 11636 8812 11688
rect 11428 11747 11480 11756
rect 11428 11713 11437 11747
rect 11437 11713 11471 11747
rect 11471 11713 11480 11747
rect 11428 11704 11480 11713
rect 11520 11747 11572 11756
rect 11520 11713 11529 11747
rect 11529 11713 11563 11747
rect 11563 11713 11572 11747
rect 11520 11704 11572 11713
rect 12440 11772 12492 11824
rect 12900 11772 12952 11824
rect 13728 11772 13780 11824
rect 9864 11679 9916 11688
rect 9864 11645 9873 11679
rect 9873 11645 9907 11679
rect 9907 11645 9916 11679
rect 9864 11636 9916 11645
rect 7656 11568 7708 11620
rect 11152 11636 11204 11688
rect 11336 11636 11388 11688
rect 11796 11679 11848 11688
rect 11796 11645 11805 11679
rect 11805 11645 11839 11679
rect 11839 11645 11848 11679
rect 11796 11636 11848 11645
rect 12348 11568 12400 11620
rect 13084 11704 13136 11756
rect 12992 11679 13044 11688
rect 12992 11645 13001 11679
rect 13001 11645 13035 11679
rect 13035 11645 13044 11679
rect 12992 11636 13044 11645
rect 13268 11679 13320 11688
rect 13268 11645 13277 11679
rect 13277 11645 13311 11679
rect 13311 11645 13320 11679
rect 13268 11636 13320 11645
rect 13084 11568 13136 11620
rect 13820 11679 13872 11688
rect 13820 11645 13829 11679
rect 13829 11645 13863 11679
rect 13863 11645 13872 11679
rect 13820 11636 13872 11645
rect 14188 11636 14240 11688
rect 14372 11704 14424 11756
rect 15016 11704 15068 11756
rect 14832 11636 14884 11688
rect 15200 11704 15252 11756
rect 15476 11747 15528 11756
rect 15476 11713 15485 11747
rect 15485 11713 15519 11747
rect 15519 11713 15528 11747
rect 15476 11704 15528 11713
rect 15568 11747 15620 11756
rect 15568 11713 15577 11747
rect 15577 11713 15611 11747
rect 15611 11713 15620 11747
rect 15568 11704 15620 11713
rect 15936 11772 15988 11824
rect 15752 11636 15804 11688
rect 16580 11679 16632 11688
rect 16580 11645 16589 11679
rect 16589 11645 16623 11679
rect 16623 11645 16632 11679
rect 16580 11636 16632 11645
rect 16672 11679 16724 11688
rect 16672 11645 16681 11679
rect 16681 11645 16715 11679
rect 16715 11645 16724 11679
rect 16672 11636 16724 11645
rect 17132 11679 17184 11688
rect 17132 11645 17141 11679
rect 17141 11645 17175 11679
rect 17175 11645 17184 11679
rect 17132 11636 17184 11645
rect 17500 11704 17552 11756
rect 17776 11704 17828 11756
rect 18144 11704 18196 11756
rect 15476 11568 15528 11620
rect 16948 11568 17000 11620
rect 3976 11500 4028 11552
rect 4252 11500 4304 11552
rect 4988 11500 5040 11552
rect 5080 11500 5132 11552
rect 5540 11500 5592 11552
rect 5816 11500 5868 11552
rect 9588 11500 9640 11552
rect 10968 11543 11020 11552
rect 10968 11509 10977 11543
rect 10977 11509 11011 11543
rect 11011 11509 11020 11543
rect 10968 11500 11020 11509
rect 11060 11543 11112 11552
rect 11060 11509 11069 11543
rect 11069 11509 11103 11543
rect 11103 11509 11112 11543
rect 11060 11500 11112 11509
rect 12808 11543 12860 11552
rect 12808 11509 12817 11543
rect 12817 11509 12851 11543
rect 12851 11509 12860 11543
rect 12808 11500 12860 11509
rect 14096 11500 14148 11552
rect 14188 11543 14240 11552
rect 14188 11509 14197 11543
rect 14197 11509 14231 11543
rect 14231 11509 14240 11543
rect 14188 11500 14240 11509
rect 14464 11500 14516 11552
rect 14832 11500 14884 11552
rect 15568 11500 15620 11552
rect 17408 11500 17460 11552
rect 18052 11568 18104 11620
rect 18880 11704 18932 11756
rect 19340 11747 19392 11756
rect 19340 11713 19349 11747
rect 19349 11713 19383 11747
rect 19383 11713 19392 11747
rect 19340 11704 19392 11713
rect 19432 11704 19484 11756
rect 19892 11704 19944 11756
rect 21088 11772 21140 11824
rect 18696 11568 18748 11620
rect 19064 11636 19116 11688
rect 19248 11636 19300 11688
rect 20168 11636 20220 11688
rect 20260 11679 20312 11688
rect 20260 11645 20269 11679
rect 20269 11645 20303 11679
rect 20303 11645 20312 11679
rect 20260 11636 20312 11645
rect 19984 11568 20036 11620
rect 19064 11500 19116 11552
rect 20260 11500 20312 11552
rect 20628 11704 20680 11756
rect 20904 11679 20956 11688
rect 20904 11645 20913 11679
rect 20913 11645 20947 11679
rect 20947 11645 20956 11679
rect 20904 11636 20956 11645
rect 21548 11704 21600 11756
rect 21456 11679 21508 11688
rect 21456 11645 21465 11679
rect 21465 11645 21499 11679
rect 21499 11645 21508 11679
rect 21456 11636 21508 11645
rect 22100 11636 22152 11688
rect 22284 11636 22336 11688
rect 20628 11568 20680 11620
rect 21548 11568 21600 11620
rect 20720 11543 20772 11552
rect 20720 11509 20729 11543
rect 20729 11509 20763 11543
rect 20763 11509 20772 11543
rect 20720 11500 20772 11509
rect 21732 11543 21784 11552
rect 21732 11509 21741 11543
rect 21741 11509 21775 11543
rect 21775 11509 21784 11543
rect 21732 11500 21784 11509
rect 22192 11500 22244 11552
rect 4366 11398 4418 11450
rect 4430 11398 4482 11450
rect 4494 11398 4546 11450
rect 4558 11398 4610 11450
rect 4622 11398 4674 11450
rect 4686 11398 4738 11450
rect 10366 11398 10418 11450
rect 10430 11398 10482 11450
rect 10494 11398 10546 11450
rect 10558 11398 10610 11450
rect 10622 11398 10674 11450
rect 10686 11398 10738 11450
rect 16366 11398 16418 11450
rect 16430 11398 16482 11450
rect 16494 11398 16546 11450
rect 16558 11398 16610 11450
rect 16622 11398 16674 11450
rect 16686 11398 16738 11450
rect 22366 11398 22418 11450
rect 22430 11398 22482 11450
rect 22494 11398 22546 11450
rect 22558 11398 22610 11450
rect 22622 11398 22674 11450
rect 22686 11398 22738 11450
rect 1676 11296 1728 11348
rect 2320 11296 2372 11348
rect 2964 11296 3016 11348
rect 3700 11296 3752 11348
rect 848 11092 900 11144
rect 1124 11160 1176 11212
rect 1308 11203 1360 11212
rect 1308 11169 1342 11203
rect 1342 11169 1360 11203
rect 1308 11160 1360 11169
rect 2780 11160 2832 11212
rect 3424 11228 3476 11280
rect 3148 11092 3200 11144
rect 2412 10999 2464 11008
rect 2412 10965 2421 10999
rect 2421 10965 2455 10999
rect 2455 10965 2464 10999
rect 2412 10956 2464 10965
rect 3148 10956 3200 11008
rect 3332 11203 3384 11212
rect 3332 11169 3341 11203
rect 3341 11169 3375 11203
rect 3375 11169 3384 11203
rect 3332 11160 3384 11169
rect 3700 11160 3752 11212
rect 4160 11160 4212 11212
rect 4896 11296 4948 11348
rect 4988 11160 5040 11212
rect 5448 11203 5500 11212
rect 5448 11169 5457 11203
rect 5457 11169 5491 11203
rect 5491 11169 5500 11203
rect 5448 11160 5500 11169
rect 5908 11160 5960 11212
rect 7012 11296 7064 11348
rect 7288 11296 7340 11348
rect 8760 11339 8812 11348
rect 8760 11305 8769 11339
rect 8769 11305 8803 11339
rect 8803 11305 8812 11339
rect 8760 11296 8812 11305
rect 9312 11296 9364 11348
rect 10140 11296 10192 11348
rect 12072 11296 12124 11348
rect 6092 11135 6144 11144
rect 6092 11101 6101 11135
rect 6101 11101 6135 11135
rect 6135 11101 6144 11135
rect 6092 11092 6144 11101
rect 6828 11160 6880 11212
rect 6552 11024 6604 11076
rect 7288 11160 7340 11212
rect 11428 11228 11480 11280
rect 8576 11203 8628 11212
rect 8576 11169 8585 11203
rect 8585 11169 8619 11203
rect 8619 11169 8628 11203
rect 8576 11160 8628 11169
rect 8668 11160 8720 11212
rect 9680 11160 9732 11212
rect 11060 11203 11112 11212
rect 11060 11169 11069 11203
rect 11069 11169 11103 11203
rect 11103 11169 11112 11203
rect 11060 11160 11112 11169
rect 11152 11160 11204 11212
rect 7104 11135 7156 11144
rect 7104 11101 7113 11135
rect 7113 11101 7147 11135
rect 7147 11101 7156 11135
rect 7104 11092 7156 11101
rect 7564 11135 7616 11144
rect 7564 11101 7573 11135
rect 7573 11101 7607 11135
rect 7607 11101 7616 11135
rect 7564 11092 7616 11101
rect 7656 11135 7708 11144
rect 7656 11101 7665 11135
rect 7665 11101 7699 11135
rect 7699 11101 7708 11135
rect 7656 11092 7708 11101
rect 8392 11092 8444 11144
rect 11520 11160 11572 11212
rect 12348 11228 12400 11280
rect 12072 11160 12124 11212
rect 13084 11228 13136 11280
rect 14004 11339 14056 11348
rect 14004 11305 14013 11339
rect 14013 11305 14047 11339
rect 14047 11305 14056 11339
rect 14004 11296 14056 11305
rect 16856 11296 16908 11348
rect 17316 11296 17368 11348
rect 17776 11296 17828 11348
rect 18604 11296 18656 11348
rect 20168 11296 20220 11348
rect 13544 11228 13596 11280
rect 8668 11024 8720 11076
rect 11520 11067 11572 11076
rect 11520 11033 11529 11067
rect 11529 11033 11563 11067
rect 11563 11033 11572 11067
rect 11520 11024 11572 11033
rect 12164 11024 12216 11076
rect 7564 10956 7616 11008
rect 8484 10956 8536 11008
rect 10784 10956 10836 11008
rect 12624 10956 12676 11008
rect 12808 10956 12860 11008
rect 13176 11160 13228 11212
rect 13360 11203 13412 11212
rect 13360 11169 13369 11203
rect 13369 11169 13403 11203
rect 13403 11169 13412 11203
rect 13360 11160 13412 11169
rect 15752 11228 15804 11280
rect 17132 11228 17184 11280
rect 14188 11160 14240 11212
rect 14464 11203 14516 11212
rect 14464 11169 14473 11203
rect 14473 11169 14507 11203
rect 14507 11169 14516 11203
rect 14464 11160 14516 11169
rect 14648 11160 14700 11212
rect 13176 11024 13228 11076
rect 14280 11092 14332 11144
rect 14924 11203 14976 11212
rect 14924 11169 14933 11203
rect 14933 11169 14967 11203
rect 14967 11169 14976 11203
rect 14924 11160 14976 11169
rect 15384 11160 15436 11212
rect 15660 11160 15712 11212
rect 16304 11203 16356 11212
rect 16304 11169 16313 11203
rect 16313 11169 16347 11203
rect 16347 11169 16356 11203
rect 16304 11160 16356 11169
rect 15200 11092 15252 11144
rect 15752 11092 15804 11144
rect 17316 11160 17368 11212
rect 17868 11160 17920 11212
rect 15292 10956 15344 11008
rect 17776 11135 17828 11144
rect 17776 11101 17785 11135
rect 17785 11101 17819 11135
rect 17819 11101 17828 11135
rect 17776 11092 17828 11101
rect 17960 11092 18012 11144
rect 18696 11203 18748 11212
rect 18696 11169 18705 11203
rect 18705 11169 18739 11203
rect 18739 11169 18748 11203
rect 18696 11160 18748 11169
rect 19064 11160 19116 11212
rect 18328 11024 18380 11076
rect 18696 11024 18748 11076
rect 19340 11092 19392 11144
rect 20076 11203 20128 11212
rect 20076 11169 20085 11203
rect 20085 11169 20119 11203
rect 20119 11169 20128 11203
rect 20076 11160 20128 11169
rect 20168 11203 20220 11212
rect 20168 11169 20177 11203
rect 20177 11169 20211 11203
rect 20211 11169 20220 11203
rect 20168 11160 20220 11169
rect 21272 11228 21324 11280
rect 21732 11228 21784 11280
rect 22192 11228 22244 11280
rect 20628 11160 20680 11212
rect 20904 11160 20956 11212
rect 21088 11203 21140 11212
rect 21088 11169 21097 11203
rect 21097 11169 21131 11203
rect 21131 11169 21140 11203
rect 21088 11160 21140 11169
rect 21548 11160 21600 11212
rect 21640 11203 21692 11212
rect 21640 11169 21649 11203
rect 21649 11169 21683 11203
rect 21683 11169 21692 11203
rect 21640 11160 21692 11169
rect 19340 10956 19392 11008
rect 19524 10956 19576 11008
rect 20260 11024 20312 11076
rect 23020 10999 23072 11008
rect 23020 10965 23029 10999
rect 23029 10965 23063 10999
rect 23063 10965 23072 10999
rect 23020 10956 23072 10965
rect 1366 10854 1418 10906
rect 1430 10854 1482 10906
rect 1494 10854 1546 10906
rect 1558 10854 1610 10906
rect 1622 10854 1674 10906
rect 1686 10854 1738 10906
rect 7366 10854 7418 10906
rect 7430 10854 7482 10906
rect 7494 10854 7546 10906
rect 7558 10854 7610 10906
rect 7622 10854 7674 10906
rect 7686 10854 7738 10906
rect 13366 10854 13418 10906
rect 13430 10854 13482 10906
rect 13494 10854 13546 10906
rect 13558 10854 13610 10906
rect 13622 10854 13674 10906
rect 13686 10854 13738 10906
rect 19366 10854 19418 10906
rect 19430 10854 19482 10906
rect 19494 10854 19546 10906
rect 19558 10854 19610 10906
rect 19622 10854 19674 10906
rect 19686 10854 19738 10906
rect 1216 10795 1268 10804
rect 1216 10761 1225 10795
rect 1225 10761 1259 10795
rect 1259 10761 1268 10795
rect 1216 10752 1268 10761
rect 1768 10752 1820 10804
rect 5448 10752 5500 10804
rect 6552 10752 6604 10804
rect 6920 10795 6972 10804
rect 6920 10761 6929 10795
rect 6929 10761 6963 10795
rect 6963 10761 6972 10795
rect 6920 10752 6972 10761
rect 7288 10752 7340 10804
rect 7748 10752 7800 10804
rect 8024 10752 8076 10804
rect 10232 10752 10284 10804
rect 1032 10684 1084 10736
rect 940 10548 992 10600
rect 2412 10616 2464 10668
rect 3332 10616 3384 10668
rect 6092 10684 6144 10736
rect 8300 10684 8352 10736
rect 5908 10659 5960 10668
rect 5908 10625 5917 10659
rect 5917 10625 5951 10659
rect 5951 10625 5960 10659
rect 5908 10616 5960 10625
rect 6000 10659 6052 10668
rect 6000 10625 6009 10659
rect 6009 10625 6043 10659
rect 6043 10625 6052 10659
rect 6000 10616 6052 10625
rect 10140 10684 10192 10736
rect 2228 10548 2280 10600
rect 3608 10548 3660 10600
rect 4344 10591 4396 10600
rect 4344 10557 4353 10591
rect 4353 10557 4387 10591
rect 4387 10557 4396 10591
rect 4344 10548 4396 10557
rect 5264 10591 5316 10600
rect 5264 10557 5273 10591
rect 5273 10557 5307 10591
rect 5307 10557 5316 10591
rect 5264 10548 5316 10557
rect 6184 10548 6236 10600
rect 6552 10591 6604 10600
rect 6552 10557 6561 10591
rect 6561 10557 6595 10591
rect 6595 10557 6604 10591
rect 6552 10548 6604 10557
rect 6828 10548 6880 10600
rect 8668 10591 8720 10600
rect 8668 10557 8677 10591
rect 8677 10557 8711 10591
rect 8711 10557 8720 10591
rect 8668 10548 8720 10557
rect 9404 10548 9456 10600
rect 1952 10480 2004 10532
rect 6460 10412 6512 10464
rect 7012 10523 7064 10532
rect 7012 10489 7021 10523
rect 7021 10489 7055 10523
rect 7055 10489 7064 10523
rect 7012 10480 7064 10489
rect 10232 10591 10284 10600
rect 10232 10557 10241 10591
rect 10241 10557 10275 10591
rect 10275 10557 10284 10591
rect 10232 10548 10284 10557
rect 10324 10591 10376 10600
rect 10324 10557 10333 10591
rect 10333 10557 10367 10591
rect 10367 10557 10376 10591
rect 10324 10548 10376 10557
rect 10876 10684 10928 10736
rect 11980 10684 12032 10736
rect 13820 10684 13872 10736
rect 14004 10752 14056 10804
rect 15200 10752 15252 10804
rect 15844 10752 15896 10804
rect 16764 10752 16816 10804
rect 16948 10752 17000 10804
rect 17592 10752 17644 10804
rect 20168 10752 20220 10804
rect 22100 10752 22152 10804
rect 22284 10752 22336 10804
rect 14372 10684 14424 10736
rect 11612 10659 11664 10668
rect 11612 10625 11621 10659
rect 11621 10625 11655 10659
rect 11655 10625 11664 10659
rect 11612 10616 11664 10625
rect 12072 10616 12124 10668
rect 12532 10616 12584 10668
rect 12900 10659 12952 10668
rect 12900 10625 12909 10659
rect 12909 10625 12943 10659
rect 12943 10625 12952 10659
rect 12900 10616 12952 10625
rect 10876 10591 10928 10600
rect 10876 10557 10885 10591
rect 10885 10557 10919 10591
rect 10919 10557 10928 10591
rect 10876 10548 10928 10557
rect 11336 10548 11388 10600
rect 11428 10591 11480 10600
rect 11428 10557 11437 10591
rect 11437 10557 11471 10591
rect 11471 10557 11480 10591
rect 11428 10548 11480 10557
rect 11980 10591 12032 10600
rect 11980 10557 11989 10591
rect 11989 10557 12023 10591
rect 12023 10557 12032 10591
rect 11980 10548 12032 10557
rect 12256 10548 12308 10600
rect 12624 10591 12676 10600
rect 12624 10557 12633 10591
rect 12633 10557 12667 10591
rect 12667 10557 12676 10591
rect 12624 10548 12676 10557
rect 8208 10412 8260 10464
rect 9956 10412 10008 10464
rect 11152 10523 11204 10532
rect 11152 10489 11161 10523
rect 11161 10489 11195 10523
rect 11195 10489 11204 10523
rect 11152 10480 11204 10489
rect 10876 10412 10928 10464
rect 12992 10548 13044 10600
rect 13360 10548 13412 10600
rect 13912 10548 13964 10600
rect 14740 10616 14792 10668
rect 15108 10659 15160 10668
rect 15108 10625 15117 10659
rect 15117 10625 15151 10659
rect 15151 10625 15160 10659
rect 15108 10616 15160 10625
rect 15292 10659 15344 10668
rect 15292 10625 15301 10659
rect 15301 10625 15335 10659
rect 15335 10625 15344 10659
rect 15292 10616 15344 10625
rect 15752 10616 15804 10668
rect 15108 10480 15160 10532
rect 15660 10548 15712 10600
rect 16212 10616 16264 10668
rect 16672 10616 16724 10668
rect 17776 10616 17828 10668
rect 18696 10659 18748 10668
rect 18696 10625 18705 10659
rect 18705 10625 18739 10659
rect 18739 10625 18748 10659
rect 18696 10616 18748 10625
rect 15292 10480 15344 10532
rect 15752 10480 15804 10532
rect 16212 10523 16264 10532
rect 16212 10489 16221 10523
rect 16221 10489 16255 10523
rect 16255 10489 16264 10523
rect 16212 10480 16264 10489
rect 16948 10591 17000 10600
rect 16948 10557 16957 10591
rect 16957 10557 16991 10591
rect 16991 10557 17000 10591
rect 16948 10548 17000 10557
rect 17316 10591 17368 10600
rect 17316 10557 17325 10591
rect 17325 10557 17359 10591
rect 17359 10557 17368 10591
rect 17316 10548 17368 10557
rect 17500 10548 17552 10600
rect 17592 10591 17644 10600
rect 17592 10557 17601 10591
rect 17601 10557 17635 10591
rect 17635 10557 17644 10591
rect 17592 10548 17644 10557
rect 17684 10548 17736 10600
rect 18420 10548 18472 10600
rect 18604 10548 18656 10600
rect 20076 10548 20128 10600
rect 21824 10659 21876 10668
rect 21824 10625 21833 10659
rect 21833 10625 21867 10659
rect 21867 10625 21876 10659
rect 21824 10616 21876 10625
rect 20536 10591 20588 10600
rect 20536 10557 20545 10591
rect 20545 10557 20579 10591
rect 20579 10557 20588 10591
rect 20536 10548 20588 10557
rect 20720 10548 20772 10600
rect 12072 10412 12124 10464
rect 12440 10455 12492 10464
rect 12440 10421 12449 10455
rect 12449 10421 12483 10455
rect 12483 10421 12492 10455
rect 12440 10412 12492 10421
rect 12716 10412 12768 10464
rect 13268 10455 13320 10464
rect 13268 10421 13277 10455
rect 13277 10421 13311 10455
rect 13311 10421 13320 10455
rect 13268 10412 13320 10421
rect 13912 10412 13964 10464
rect 14280 10412 14332 10464
rect 14464 10455 14516 10464
rect 14464 10421 14473 10455
rect 14473 10421 14507 10455
rect 14507 10421 14516 10455
rect 14464 10412 14516 10421
rect 19064 10480 19116 10532
rect 16396 10412 16448 10464
rect 17040 10412 17092 10464
rect 17316 10412 17368 10464
rect 17960 10412 18012 10464
rect 18328 10412 18380 10464
rect 19432 10412 19484 10464
rect 20168 10480 20220 10532
rect 21088 10548 21140 10600
rect 23388 10616 23440 10668
rect 23020 10591 23072 10600
rect 23020 10557 23029 10591
rect 23029 10557 23063 10591
rect 23063 10557 23072 10591
rect 23020 10548 23072 10557
rect 20076 10412 20128 10464
rect 20904 10412 20956 10464
rect 22836 10412 22888 10464
rect 22928 10455 22980 10464
rect 22928 10421 22937 10455
rect 22937 10421 22971 10455
rect 22971 10421 22980 10455
rect 22928 10412 22980 10421
rect 4366 10310 4418 10362
rect 4430 10310 4482 10362
rect 4494 10310 4546 10362
rect 4558 10310 4610 10362
rect 4622 10310 4674 10362
rect 4686 10310 4738 10362
rect 10366 10310 10418 10362
rect 10430 10310 10482 10362
rect 10494 10310 10546 10362
rect 10558 10310 10610 10362
rect 10622 10310 10674 10362
rect 10686 10310 10738 10362
rect 16366 10310 16418 10362
rect 16430 10310 16482 10362
rect 16494 10310 16546 10362
rect 16558 10310 16610 10362
rect 16622 10310 16674 10362
rect 16686 10310 16738 10362
rect 22366 10310 22418 10362
rect 22430 10310 22482 10362
rect 22494 10310 22546 10362
rect 22558 10310 22610 10362
rect 22622 10310 22674 10362
rect 22686 10310 22738 10362
rect 3608 10251 3660 10260
rect 3608 10217 3617 10251
rect 3617 10217 3651 10251
rect 3651 10217 3660 10251
rect 3608 10208 3660 10217
rect 5264 10208 5316 10260
rect 5448 10208 5500 10260
rect 4068 10140 4120 10192
rect 848 10115 900 10124
rect 848 10081 857 10115
rect 857 10081 891 10115
rect 891 10081 900 10115
rect 848 10072 900 10081
rect 1124 10115 1176 10124
rect 1124 10081 1158 10115
rect 1158 10081 1176 10115
rect 1124 10072 1176 10081
rect 1952 10072 2004 10124
rect 2596 10115 2648 10124
rect 2596 10081 2605 10115
rect 2605 10081 2639 10115
rect 2639 10081 2648 10115
rect 2596 10072 2648 10081
rect 3148 10115 3200 10124
rect 3148 10081 3157 10115
rect 3157 10081 3191 10115
rect 3191 10081 3200 10115
rect 3148 10072 3200 10081
rect 3976 10115 4028 10124
rect 3976 10081 3985 10115
rect 3985 10081 4019 10115
rect 4019 10081 4028 10115
rect 3976 10072 4028 10081
rect 5816 10140 5868 10192
rect 6184 10183 6236 10192
rect 6184 10149 6193 10183
rect 6193 10149 6227 10183
rect 6227 10149 6236 10183
rect 6184 10140 6236 10149
rect 8484 10208 8536 10260
rect 11152 10208 11204 10260
rect 11888 10208 11940 10260
rect 12624 10208 12676 10260
rect 12900 10208 12952 10260
rect 13084 10208 13136 10260
rect 6552 10072 6604 10124
rect 7104 10072 7156 10124
rect 7288 10072 7340 10124
rect 7012 10004 7064 10056
rect 8392 10140 8444 10192
rect 8208 10115 8260 10124
rect 8208 10081 8217 10115
rect 8217 10081 8251 10115
rect 8251 10081 8260 10115
rect 8208 10072 8260 10081
rect 8760 10115 8812 10124
rect 8760 10081 8769 10115
rect 8769 10081 8803 10115
rect 8803 10081 8812 10115
rect 8760 10072 8812 10081
rect 9036 10072 9088 10124
rect 9220 10115 9272 10124
rect 9220 10081 9229 10115
rect 9229 10081 9263 10115
rect 9263 10081 9272 10115
rect 9220 10072 9272 10081
rect 9404 10072 9456 10124
rect 10968 10140 11020 10192
rect 11428 10140 11480 10192
rect 12348 10140 12400 10192
rect 9956 10115 10008 10124
rect 9956 10081 9965 10115
rect 9965 10081 9999 10115
rect 9999 10081 10008 10115
rect 9956 10072 10008 10081
rect 3608 9936 3660 9988
rect 5540 9936 5592 9988
rect 10140 10072 10192 10124
rect 10508 10115 10560 10124
rect 10508 10081 10517 10115
rect 10517 10081 10551 10115
rect 10551 10081 10560 10115
rect 10508 10072 10560 10081
rect 11704 10072 11756 10124
rect 11888 10072 11940 10124
rect 2136 9868 2188 9920
rect 2964 9911 3016 9920
rect 2964 9877 2973 9911
rect 2973 9877 3007 9911
rect 3007 9877 3016 9911
rect 2964 9868 3016 9877
rect 3424 9911 3476 9920
rect 3424 9877 3433 9911
rect 3433 9877 3467 9911
rect 3467 9877 3476 9911
rect 3424 9868 3476 9877
rect 4252 9868 4304 9920
rect 5632 9868 5684 9920
rect 7196 9911 7248 9920
rect 7196 9877 7205 9911
rect 7205 9877 7239 9911
rect 7239 9877 7248 9911
rect 7196 9868 7248 9877
rect 8024 9868 8076 9920
rect 10140 9936 10192 9988
rect 11980 9936 12032 9988
rect 12900 10004 12952 10056
rect 13360 10115 13412 10124
rect 13360 10081 13369 10115
rect 13369 10081 13403 10115
rect 13403 10081 13412 10115
rect 13360 10072 13412 10081
rect 13636 10115 13688 10124
rect 13636 10081 13645 10115
rect 13645 10081 13679 10115
rect 13679 10081 13688 10115
rect 15476 10140 15528 10192
rect 13636 10072 13688 10081
rect 14556 10072 14608 10124
rect 15292 10072 15344 10124
rect 15844 10208 15896 10260
rect 15752 10183 15804 10192
rect 15752 10149 15761 10183
rect 15761 10149 15795 10183
rect 15795 10149 15804 10183
rect 17960 10208 18012 10260
rect 18420 10208 18472 10260
rect 15752 10140 15804 10149
rect 13452 10004 13504 10056
rect 13820 10004 13872 10056
rect 14832 10004 14884 10056
rect 14924 10004 14976 10056
rect 16120 10115 16172 10124
rect 16120 10081 16129 10115
rect 16129 10081 16163 10115
rect 16163 10081 16172 10115
rect 16120 10072 16172 10081
rect 16304 10115 16356 10124
rect 16304 10081 16313 10115
rect 16313 10081 16347 10115
rect 16347 10081 16356 10115
rect 16304 10072 16356 10081
rect 18236 10072 18288 10124
rect 18328 10115 18380 10124
rect 18328 10081 18337 10115
rect 18337 10081 18371 10115
rect 18371 10081 18380 10115
rect 18328 10072 18380 10081
rect 19248 10140 19300 10192
rect 19892 10208 19944 10260
rect 21272 10208 21324 10260
rect 21456 10251 21508 10260
rect 21456 10217 21465 10251
rect 21465 10217 21499 10251
rect 21499 10217 21508 10251
rect 21456 10208 21508 10217
rect 20076 10140 20128 10192
rect 21548 10140 21600 10192
rect 19616 10115 19668 10124
rect 19616 10081 19625 10115
rect 19625 10081 19659 10115
rect 19659 10081 19668 10115
rect 19616 10072 19668 10081
rect 19984 10072 20036 10124
rect 20536 10072 20588 10124
rect 20720 10072 20772 10124
rect 22652 10140 22704 10192
rect 22928 10140 22980 10192
rect 23204 10072 23256 10124
rect 8576 9868 8628 9920
rect 9128 9911 9180 9920
rect 9128 9877 9137 9911
rect 9137 9877 9171 9911
rect 9171 9877 9180 9911
rect 9128 9868 9180 9877
rect 9404 9911 9456 9920
rect 9404 9877 9413 9911
rect 9413 9877 9447 9911
rect 9447 9877 9456 9911
rect 9404 9868 9456 9877
rect 9588 9868 9640 9920
rect 10508 9868 10560 9920
rect 11704 9868 11756 9920
rect 12072 9911 12124 9920
rect 12072 9877 12081 9911
rect 12081 9877 12115 9911
rect 12115 9877 12124 9911
rect 12072 9868 12124 9877
rect 12532 9868 12584 9920
rect 12808 9868 12860 9920
rect 15016 9979 15068 9988
rect 15016 9945 15025 9979
rect 15025 9945 15059 9979
rect 15059 9945 15068 9979
rect 15016 9936 15068 9945
rect 15292 9936 15344 9988
rect 16396 9936 16448 9988
rect 17500 9936 17552 9988
rect 18144 9936 18196 9988
rect 20260 10004 20312 10056
rect 21272 10047 21324 10056
rect 21272 10013 21281 10047
rect 21281 10013 21315 10047
rect 21315 10013 21324 10047
rect 21272 10004 21324 10013
rect 20168 9936 20220 9988
rect 19064 9868 19116 9920
rect 19432 9868 19484 9920
rect 19984 9868 20036 9920
rect 20904 9936 20956 9988
rect 21456 9936 21508 9988
rect 20352 9868 20404 9920
rect 21548 9868 21600 9920
rect 22468 9936 22520 9988
rect 22744 9868 22796 9920
rect 1366 9766 1418 9818
rect 1430 9766 1482 9818
rect 1494 9766 1546 9818
rect 1558 9766 1610 9818
rect 1622 9766 1674 9818
rect 1686 9766 1738 9818
rect 7366 9766 7418 9818
rect 7430 9766 7482 9818
rect 7494 9766 7546 9818
rect 7558 9766 7610 9818
rect 7622 9766 7674 9818
rect 7686 9766 7738 9818
rect 13366 9766 13418 9818
rect 13430 9766 13482 9818
rect 13494 9766 13546 9818
rect 13558 9766 13610 9818
rect 13622 9766 13674 9818
rect 13686 9766 13738 9818
rect 19366 9766 19418 9818
rect 19430 9766 19482 9818
rect 19494 9766 19546 9818
rect 19558 9766 19610 9818
rect 19622 9766 19674 9818
rect 19686 9766 19738 9818
rect 1952 9664 2004 9716
rect 1676 9596 1728 9648
rect 3424 9528 3476 9580
rect 4068 9596 4120 9648
rect 4804 9664 4856 9716
rect 4252 9596 4304 9648
rect 572 9460 624 9512
rect 1400 9503 1452 9512
rect 1400 9469 1409 9503
rect 1409 9469 1443 9503
rect 1443 9469 1452 9503
rect 1400 9460 1452 9469
rect 2596 9460 2648 9512
rect 3608 9503 3660 9512
rect 3608 9469 3617 9503
rect 3617 9469 3651 9503
rect 3651 9469 3660 9503
rect 3608 9460 3660 9469
rect 2044 9367 2096 9376
rect 2044 9333 2053 9367
rect 2053 9333 2087 9367
rect 2087 9333 2096 9367
rect 2044 9324 2096 9333
rect 3056 9324 3108 9376
rect 3332 9324 3384 9376
rect 4344 9571 4396 9580
rect 4344 9537 4353 9571
rect 4353 9537 4387 9571
rect 4387 9537 4396 9571
rect 4344 9528 4396 9537
rect 3976 9503 4028 9512
rect 3976 9469 3985 9503
rect 3985 9469 4019 9503
rect 4019 9469 4028 9503
rect 3976 9460 4028 9469
rect 4160 9503 4212 9512
rect 4160 9469 4169 9503
rect 4169 9469 4203 9503
rect 4203 9469 4212 9503
rect 4160 9460 4212 9469
rect 7288 9664 7340 9716
rect 7564 9664 7616 9716
rect 8300 9664 8352 9716
rect 8760 9664 8812 9716
rect 8852 9664 8904 9716
rect 9404 9664 9456 9716
rect 8392 9596 8444 9648
rect 12072 9664 12124 9716
rect 6092 9571 6144 9580
rect 4068 9435 4120 9444
rect 4068 9401 4077 9435
rect 4077 9401 4111 9435
rect 4111 9401 4120 9435
rect 5540 9460 5592 9512
rect 5632 9503 5684 9512
rect 5632 9469 5641 9503
rect 5641 9469 5675 9503
rect 5675 9469 5684 9503
rect 5632 9460 5684 9469
rect 6092 9537 6101 9571
rect 6101 9537 6135 9571
rect 6135 9537 6144 9571
rect 6092 9528 6144 9537
rect 6276 9460 6328 9512
rect 6368 9460 6420 9512
rect 6552 9460 6604 9512
rect 7196 9528 7248 9580
rect 7564 9460 7616 9512
rect 8208 9528 8260 9580
rect 8484 9528 8536 9580
rect 8668 9528 8720 9580
rect 8944 9571 8996 9580
rect 8944 9537 8953 9571
rect 8953 9537 8987 9571
rect 8987 9537 8996 9571
rect 8944 9528 8996 9537
rect 9404 9528 9456 9580
rect 10784 9596 10836 9648
rect 12716 9664 12768 9716
rect 8024 9460 8076 9512
rect 8576 9503 8628 9512
rect 8576 9469 8585 9503
rect 8585 9469 8619 9503
rect 8619 9469 8628 9503
rect 8576 9460 8628 9469
rect 4068 9392 4120 9401
rect 3976 9324 4028 9376
rect 7104 9392 7156 9444
rect 7288 9392 7340 9444
rect 8668 9392 8720 9444
rect 9036 9392 9088 9444
rect 9680 9503 9732 9512
rect 9680 9469 9689 9503
rect 9689 9469 9723 9503
rect 9723 9469 9732 9503
rect 9680 9460 9732 9469
rect 11612 9571 11664 9580
rect 11612 9537 11621 9571
rect 11621 9537 11655 9571
rect 11655 9537 11664 9571
rect 11612 9528 11664 9537
rect 10692 9503 10744 9512
rect 10692 9469 10701 9503
rect 10701 9469 10735 9503
rect 10735 9469 10744 9503
rect 10692 9460 10744 9469
rect 10876 9460 10928 9512
rect 11060 9460 11112 9512
rect 11152 9503 11204 9512
rect 11152 9469 11161 9503
rect 11161 9469 11195 9503
rect 11195 9469 11204 9503
rect 11152 9460 11204 9469
rect 11336 9460 11388 9512
rect 11428 9503 11480 9512
rect 11428 9469 11437 9503
rect 11437 9469 11471 9503
rect 11471 9469 11480 9503
rect 11428 9460 11480 9469
rect 12256 9528 12308 9580
rect 13084 9596 13136 9648
rect 13268 9596 13320 9648
rect 12900 9571 12952 9580
rect 12900 9537 12909 9571
rect 12909 9537 12943 9571
rect 12943 9537 12952 9571
rect 12900 9528 12952 9537
rect 5264 9367 5316 9376
rect 5264 9333 5273 9367
rect 5273 9333 5307 9367
rect 5307 9333 5316 9367
rect 5264 9324 5316 9333
rect 8208 9324 8260 9376
rect 8760 9324 8812 9376
rect 10048 9392 10100 9444
rect 10324 9435 10376 9444
rect 10324 9401 10333 9435
rect 10333 9401 10367 9435
rect 10367 9401 10376 9435
rect 10324 9392 10376 9401
rect 12716 9503 12768 9512
rect 12716 9469 12725 9503
rect 12725 9469 12759 9503
rect 12759 9469 12768 9503
rect 12716 9460 12768 9469
rect 14648 9664 14700 9716
rect 19892 9664 19944 9716
rect 20076 9664 20128 9716
rect 20628 9664 20680 9716
rect 21732 9707 21784 9716
rect 21732 9673 21741 9707
rect 21741 9673 21775 9707
rect 21775 9673 21784 9707
rect 21732 9664 21784 9673
rect 14096 9596 14148 9648
rect 14740 9596 14792 9648
rect 15016 9596 15068 9648
rect 15844 9528 15896 9580
rect 16304 9528 16356 9580
rect 16396 9571 16448 9580
rect 16396 9537 16405 9571
rect 16405 9537 16439 9571
rect 16439 9537 16448 9571
rect 16396 9528 16448 9537
rect 11060 9324 11112 9376
rect 11704 9324 11756 9376
rect 12808 9392 12860 9444
rect 13820 9503 13872 9512
rect 13820 9469 13829 9503
rect 13829 9469 13863 9503
rect 13863 9469 13872 9503
rect 13820 9460 13872 9469
rect 14280 9503 14332 9512
rect 14280 9469 14289 9503
rect 14289 9469 14323 9503
rect 14323 9469 14332 9503
rect 14280 9460 14332 9469
rect 14740 9460 14792 9512
rect 16672 9503 16724 9512
rect 16672 9469 16681 9503
rect 16681 9469 16715 9503
rect 16715 9469 16724 9503
rect 16672 9460 16724 9469
rect 14648 9392 14700 9444
rect 15660 9392 15712 9444
rect 17316 9503 17368 9512
rect 17316 9469 17325 9503
rect 17325 9469 17359 9503
rect 17359 9469 17368 9503
rect 17316 9460 17368 9469
rect 17592 9503 17644 9512
rect 17592 9469 17601 9503
rect 17601 9469 17635 9503
rect 17635 9469 17644 9503
rect 17592 9460 17644 9469
rect 19064 9596 19116 9648
rect 19892 9528 19944 9580
rect 20996 9596 21048 9648
rect 21088 9596 21140 9648
rect 21548 9596 21600 9648
rect 17868 9503 17920 9512
rect 17868 9469 17877 9503
rect 17877 9469 17911 9503
rect 17911 9469 17920 9503
rect 17868 9460 17920 9469
rect 18236 9392 18288 9444
rect 19432 9503 19484 9512
rect 19432 9469 19441 9503
rect 19441 9469 19475 9503
rect 19475 9469 19484 9503
rect 19432 9460 19484 9469
rect 20076 9460 20128 9512
rect 20352 9460 20404 9512
rect 21272 9460 21324 9512
rect 22468 9503 22520 9512
rect 22468 9469 22477 9503
rect 22477 9469 22511 9503
rect 22511 9469 22520 9503
rect 22468 9460 22520 9469
rect 22652 9503 22704 9512
rect 22652 9469 22661 9503
rect 22661 9469 22695 9503
rect 22695 9469 22704 9503
rect 22652 9460 22704 9469
rect 13268 9367 13320 9376
rect 13268 9333 13277 9367
rect 13277 9333 13311 9367
rect 13311 9333 13320 9367
rect 13268 9324 13320 9333
rect 14004 9367 14056 9376
rect 14004 9333 14013 9367
rect 14013 9333 14047 9367
rect 14047 9333 14056 9367
rect 14004 9324 14056 9333
rect 14280 9324 14332 9376
rect 17040 9367 17092 9376
rect 17040 9333 17049 9367
rect 17049 9333 17083 9367
rect 17083 9333 17092 9367
rect 17040 9324 17092 9333
rect 17684 9324 17736 9376
rect 18144 9324 18196 9376
rect 22928 9503 22980 9512
rect 22928 9469 22937 9503
rect 22937 9469 22971 9503
rect 22971 9469 22980 9503
rect 22928 9460 22980 9469
rect 22836 9392 22888 9444
rect 19248 9324 19300 9376
rect 20076 9324 20128 9376
rect 20444 9367 20496 9376
rect 20444 9333 20453 9367
rect 20453 9333 20487 9367
rect 20487 9333 20496 9367
rect 20444 9324 20496 9333
rect 21272 9324 21324 9376
rect 21824 9324 21876 9376
rect 4366 9222 4418 9274
rect 4430 9222 4482 9274
rect 4494 9222 4546 9274
rect 4558 9222 4610 9274
rect 4622 9222 4674 9274
rect 4686 9222 4738 9274
rect 10366 9222 10418 9274
rect 10430 9222 10482 9274
rect 10494 9222 10546 9274
rect 10558 9222 10610 9274
rect 10622 9222 10674 9274
rect 10686 9222 10738 9274
rect 16366 9222 16418 9274
rect 16430 9222 16482 9274
rect 16494 9222 16546 9274
rect 16558 9222 16610 9274
rect 16622 9222 16674 9274
rect 16686 9222 16738 9274
rect 22366 9222 22418 9274
rect 22430 9222 22482 9274
rect 22494 9222 22546 9274
rect 22558 9222 22610 9274
rect 22622 9222 22674 9274
rect 22686 9222 22738 9274
rect 1124 9163 1176 9172
rect 1124 9129 1133 9163
rect 1133 9129 1167 9163
rect 1167 9129 1176 9163
rect 1124 9120 1176 9129
rect 1584 9163 1636 9172
rect 1124 8984 1176 9036
rect 1584 9129 1593 9163
rect 1593 9129 1627 9163
rect 1627 9129 1636 9163
rect 1584 9120 1636 9129
rect 1860 9052 1912 9104
rect 2596 9120 2648 9172
rect 3332 9120 3384 9172
rect 3792 9120 3844 9172
rect 4252 9120 4304 9172
rect 6276 9163 6328 9172
rect 6276 9129 6285 9163
rect 6285 9129 6319 9163
rect 6319 9129 6328 9163
rect 6276 9120 6328 9129
rect 7840 9120 7892 9172
rect 8116 9120 8168 9172
rect 8300 9120 8352 9172
rect 2872 9052 2924 9104
rect 4160 9052 4212 9104
rect 4988 9052 5040 9104
rect 6184 9052 6236 9104
rect 11152 9095 11204 9104
rect 1768 9027 1820 9036
rect 1768 8993 1777 9027
rect 1777 8993 1811 9027
rect 1811 8993 1820 9027
rect 1768 8984 1820 8993
rect 1032 8916 1084 8968
rect 1676 8916 1728 8968
rect 2780 9027 2832 9036
rect 2780 8993 2789 9027
rect 2789 8993 2823 9027
rect 2823 8993 2832 9027
rect 2780 8984 2832 8993
rect 2964 9027 3016 9036
rect 2964 8993 2973 9027
rect 2973 8993 3007 9027
rect 3007 8993 3016 9027
rect 2964 8984 3016 8993
rect 3056 9027 3108 9036
rect 3056 8993 3065 9027
rect 3065 8993 3099 9027
rect 3099 8993 3108 9027
rect 3056 8984 3108 8993
rect 3516 8984 3568 9036
rect 4068 8984 4120 9036
rect 4804 8984 4856 9036
rect 5632 8984 5684 9036
rect 5908 8984 5960 9036
rect 6920 8984 6972 9036
rect 7104 8984 7156 9036
rect 7288 8984 7340 9036
rect 8300 8984 8352 9036
rect 11152 9061 11161 9095
rect 11161 9061 11195 9095
rect 11195 9061 11204 9095
rect 11152 9052 11204 9061
rect 11336 9163 11388 9172
rect 11336 9129 11345 9163
rect 11345 9129 11379 9163
rect 11379 9129 11388 9163
rect 11336 9120 11388 9129
rect 11428 9120 11480 9172
rect 12532 9120 12584 9172
rect 9772 8984 9824 9036
rect 3792 8916 3844 8968
rect 5356 8916 5408 8968
rect 6368 8916 6420 8968
rect 2044 8780 2096 8832
rect 7196 8848 7248 8900
rect 7748 8916 7800 8968
rect 8116 8959 8168 8968
rect 8116 8925 8125 8959
rect 8125 8925 8159 8959
rect 8159 8925 8168 8959
rect 8116 8916 8168 8925
rect 11060 8984 11112 9036
rect 13820 9052 13872 9104
rect 12164 8984 12216 9036
rect 14096 9027 14148 9036
rect 14096 8993 14105 9027
rect 14105 8993 14139 9027
rect 14139 8993 14148 9027
rect 14096 8984 14148 8993
rect 10416 8916 10468 8968
rect 14740 9027 14792 9036
rect 14740 8993 14749 9027
rect 14749 8993 14783 9027
rect 14783 8993 14792 9027
rect 14740 8984 14792 8993
rect 15016 8984 15068 9036
rect 15108 9027 15160 9036
rect 15108 8993 15117 9027
rect 15117 8993 15151 9027
rect 15151 8993 15160 9027
rect 15108 8984 15160 8993
rect 17776 9120 17828 9172
rect 17132 9052 17184 9104
rect 17592 9052 17644 9104
rect 18144 9120 18196 9172
rect 19248 9120 19300 9172
rect 21916 9120 21968 9172
rect 22652 9120 22704 9172
rect 22928 9120 22980 9172
rect 15844 8984 15896 9036
rect 8944 8848 8996 8900
rect 10876 8848 10928 8900
rect 11336 8848 11388 8900
rect 15752 8916 15804 8968
rect 16304 8916 16356 8968
rect 16580 8916 16632 8968
rect 17224 8916 17276 8968
rect 18236 9027 18288 9036
rect 18236 8993 18265 9027
rect 18265 8993 18288 9027
rect 18236 8984 18288 8993
rect 18512 9027 18564 9036
rect 18512 8993 18521 9027
rect 18521 8993 18555 9027
rect 18555 8993 18564 9027
rect 18512 8984 18564 8993
rect 21732 9052 21784 9104
rect 22284 9052 22336 9104
rect 19064 9027 19116 9036
rect 19064 8993 19073 9027
rect 19073 8993 19107 9027
rect 19107 8993 19116 9027
rect 19064 8984 19116 8993
rect 19708 8984 19760 9036
rect 19892 8984 19944 9036
rect 21456 9027 21508 9036
rect 21456 8993 21465 9027
rect 21465 8993 21499 9027
rect 21499 8993 21508 9027
rect 21456 8984 21508 8993
rect 22100 8984 22152 9036
rect 22652 9027 22704 9036
rect 22652 8993 22661 9027
rect 22661 8993 22695 9027
rect 22695 8993 22704 9027
rect 22652 8984 22704 8993
rect 3516 8780 3568 8832
rect 4160 8823 4212 8832
rect 4160 8789 4169 8823
rect 4169 8789 4203 8823
rect 4203 8789 4212 8823
rect 4160 8780 4212 8789
rect 5540 8780 5592 8832
rect 6920 8780 6972 8832
rect 7104 8780 7156 8832
rect 7748 8780 7800 8832
rect 8576 8780 8628 8832
rect 9680 8780 9732 8832
rect 11704 8780 11756 8832
rect 11980 8780 12032 8832
rect 12256 8780 12308 8832
rect 12348 8780 12400 8832
rect 12900 8780 12952 8832
rect 13820 8780 13872 8832
rect 14556 8823 14608 8832
rect 14556 8789 14565 8823
rect 14565 8789 14599 8823
rect 14599 8789 14608 8823
rect 14556 8780 14608 8789
rect 14648 8780 14700 8832
rect 15108 8780 15160 8832
rect 16672 8848 16724 8900
rect 18512 8848 18564 8900
rect 19892 8891 19944 8900
rect 19892 8857 19901 8891
rect 19901 8857 19935 8891
rect 19935 8857 19944 8891
rect 19892 8848 19944 8857
rect 20352 8848 20404 8900
rect 20720 8848 20772 8900
rect 16028 8780 16080 8832
rect 16856 8780 16908 8832
rect 18420 8780 18472 8832
rect 18880 8780 18932 8832
rect 19800 8780 19852 8832
rect 20628 8780 20680 8832
rect 21088 8780 21140 8832
rect 1366 8678 1418 8730
rect 1430 8678 1482 8730
rect 1494 8678 1546 8730
rect 1558 8678 1610 8730
rect 1622 8678 1674 8730
rect 1686 8678 1738 8730
rect 7366 8678 7418 8730
rect 7430 8678 7482 8730
rect 7494 8678 7546 8730
rect 7558 8678 7610 8730
rect 7622 8678 7674 8730
rect 7686 8678 7738 8730
rect 13366 8678 13418 8730
rect 13430 8678 13482 8730
rect 13494 8678 13546 8730
rect 13558 8678 13610 8730
rect 13622 8678 13674 8730
rect 13686 8678 13738 8730
rect 19366 8678 19418 8730
rect 19430 8678 19482 8730
rect 19494 8678 19546 8730
rect 19558 8678 19610 8730
rect 19622 8678 19674 8730
rect 19686 8678 19738 8730
rect 1952 8576 2004 8628
rect 2504 8576 2556 8628
rect 3516 8619 3568 8628
rect 3516 8585 3525 8619
rect 3525 8585 3559 8619
rect 3559 8585 3568 8619
rect 3516 8576 3568 8585
rect 4804 8576 4856 8628
rect 2044 8372 2096 8424
rect 2228 8415 2280 8424
rect 2228 8381 2237 8415
rect 2237 8381 2271 8415
rect 2271 8381 2280 8415
rect 2228 8372 2280 8381
rect 5172 8508 5224 8560
rect 5724 8619 5776 8628
rect 5724 8585 5733 8619
rect 5733 8585 5767 8619
rect 5767 8585 5776 8619
rect 5724 8576 5776 8585
rect 6552 8576 6604 8628
rect 8944 8576 8996 8628
rect 9496 8576 9548 8628
rect 9588 8576 9640 8628
rect 9404 8508 9456 8560
rect 4804 8483 4856 8492
rect 4804 8449 4813 8483
rect 4813 8449 4847 8483
rect 4847 8449 4856 8483
rect 4804 8440 4856 8449
rect 5356 8440 5408 8492
rect 3148 8372 3200 8424
rect 3516 8372 3568 8424
rect 3516 8236 3568 8288
rect 3792 8236 3844 8288
rect 4068 8347 4120 8356
rect 4068 8313 4077 8347
rect 4077 8313 4111 8347
rect 4111 8313 4120 8347
rect 4068 8304 4120 8313
rect 4896 8372 4948 8424
rect 6092 8372 6144 8424
rect 6368 8440 6420 8492
rect 6736 8440 6788 8492
rect 7104 8440 7156 8492
rect 8392 8483 8444 8492
rect 8392 8449 8401 8483
rect 8401 8449 8435 8483
rect 8435 8449 8444 8483
rect 8392 8440 8444 8449
rect 8944 8440 8996 8492
rect 9864 8508 9916 8560
rect 10048 8508 10100 8560
rect 6276 8415 6328 8424
rect 6276 8381 6285 8415
rect 6285 8381 6319 8415
rect 6319 8381 6328 8415
rect 6276 8372 6328 8381
rect 7748 8372 7800 8424
rect 8300 8372 8352 8424
rect 8576 8372 8628 8424
rect 4896 8236 4948 8288
rect 9220 8304 9272 8356
rect 6092 8279 6144 8288
rect 6092 8245 6101 8279
rect 6101 8245 6135 8279
rect 6135 8245 6144 8279
rect 6092 8236 6144 8245
rect 8944 8236 8996 8288
rect 9588 8415 9640 8424
rect 9588 8381 9597 8415
rect 9597 8381 9631 8415
rect 9631 8381 9640 8415
rect 9588 8372 9640 8381
rect 9680 8415 9732 8424
rect 9680 8381 9689 8415
rect 9689 8381 9723 8415
rect 9723 8381 9732 8415
rect 9680 8372 9732 8381
rect 10324 8415 10376 8424
rect 10324 8381 10333 8415
rect 10333 8381 10367 8415
rect 10367 8381 10376 8415
rect 10324 8372 10376 8381
rect 10416 8415 10468 8424
rect 10416 8381 10425 8415
rect 10425 8381 10459 8415
rect 10459 8381 10468 8415
rect 10416 8372 10468 8381
rect 11152 8576 11204 8628
rect 12164 8576 12216 8628
rect 11060 8508 11112 8560
rect 12348 8508 12400 8560
rect 12624 8508 12676 8560
rect 11336 8440 11388 8492
rect 10876 8372 10928 8424
rect 11704 8415 11756 8424
rect 11704 8381 11713 8415
rect 11713 8381 11747 8415
rect 11747 8381 11756 8415
rect 11704 8372 11756 8381
rect 11796 8415 11848 8424
rect 11796 8381 11805 8415
rect 11805 8381 11839 8415
rect 11839 8381 11848 8415
rect 11796 8372 11848 8381
rect 11888 8372 11940 8424
rect 12440 8415 12492 8424
rect 12440 8381 12449 8415
rect 12449 8381 12483 8415
rect 12483 8381 12492 8415
rect 12440 8372 12492 8381
rect 15476 8508 15528 8560
rect 15752 8508 15804 8560
rect 16764 8508 16816 8560
rect 17132 8508 17184 8560
rect 12808 8415 12860 8424
rect 12808 8381 12817 8415
rect 12817 8381 12851 8415
rect 12851 8381 12860 8415
rect 12808 8372 12860 8381
rect 13820 8483 13872 8492
rect 13820 8449 13829 8483
rect 13829 8449 13863 8483
rect 13863 8449 13872 8483
rect 13820 8440 13872 8449
rect 15844 8440 15896 8492
rect 12992 8415 13044 8424
rect 12992 8381 13001 8415
rect 13001 8381 13035 8415
rect 13035 8381 13044 8415
rect 12992 8372 13044 8381
rect 13084 8372 13136 8424
rect 13544 8415 13596 8424
rect 13544 8381 13553 8415
rect 13553 8381 13587 8415
rect 13587 8381 13596 8415
rect 13544 8372 13596 8381
rect 14096 8415 14148 8424
rect 14096 8381 14105 8415
rect 14105 8381 14139 8415
rect 14139 8381 14148 8415
rect 14096 8372 14148 8381
rect 15108 8372 15160 8424
rect 16028 8415 16080 8424
rect 16028 8381 16037 8415
rect 16037 8381 16071 8415
rect 16071 8381 16080 8415
rect 16028 8372 16080 8381
rect 9496 8236 9548 8288
rect 9864 8236 9916 8288
rect 11520 8279 11572 8288
rect 11520 8245 11529 8279
rect 11529 8245 11563 8279
rect 11563 8245 11572 8279
rect 11520 8236 11572 8245
rect 11796 8236 11848 8288
rect 15016 8304 15068 8356
rect 15292 8304 15344 8356
rect 16304 8415 16356 8424
rect 16304 8381 16313 8415
rect 16313 8381 16347 8415
rect 16347 8381 16356 8415
rect 16304 8372 16356 8381
rect 16580 8415 16632 8424
rect 16580 8381 16589 8415
rect 16589 8381 16623 8415
rect 16623 8381 16632 8415
rect 16580 8372 16632 8381
rect 16856 8415 16908 8424
rect 16856 8381 16865 8415
rect 16865 8381 16899 8415
rect 16899 8381 16908 8415
rect 16856 8372 16908 8381
rect 13084 8236 13136 8288
rect 14464 8236 14516 8288
rect 14556 8236 14608 8288
rect 14832 8236 14884 8288
rect 16764 8347 16816 8356
rect 16764 8313 16773 8347
rect 16773 8313 16807 8347
rect 16807 8313 16816 8347
rect 16764 8304 16816 8313
rect 17132 8415 17184 8424
rect 17132 8381 17141 8415
rect 17141 8381 17175 8415
rect 17175 8381 17184 8415
rect 17132 8372 17184 8381
rect 17868 8508 17920 8560
rect 17592 8440 17644 8492
rect 18144 8551 18196 8560
rect 18144 8517 18153 8551
rect 18153 8517 18187 8551
rect 18187 8517 18196 8551
rect 18144 8508 18196 8517
rect 18972 8576 19024 8628
rect 20352 8576 20404 8628
rect 21088 8576 21140 8628
rect 21180 8619 21232 8628
rect 21180 8585 21189 8619
rect 21189 8585 21223 8619
rect 21223 8585 21232 8619
rect 21180 8576 21232 8585
rect 18420 8508 18472 8560
rect 22008 8508 22060 8560
rect 20352 8440 20404 8492
rect 17592 8347 17644 8356
rect 17592 8313 17601 8347
rect 17601 8313 17635 8347
rect 17635 8313 17644 8347
rect 17592 8304 17644 8313
rect 18420 8372 18472 8424
rect 20720 8372 20772 8424
rect 21272 8372 21324 8424
rect 21456 8415 21508 8424
rect 21456 8381 21465 8415
rect 21465 8381 21499 8415
rect 21499 8381 21508 8415
rect 21456 8372 21508 8381
rect 21916 8415 21968 8424
rect 21916 8381 21925 8415
rect 21925 8381 21959 8415
rect 21959 8381 21968 8415
rect 21916 8372 21968 8381
rect 22192 8415 22244 8424
rect 22192 8381 22201 8415
rect 22201 8381 22235 8415
rect 22235 8381 22244 8415
rect 22192 8372 22244 8381
rect 17684 8279 17736 8288
rect 17684 8245 17693 8279
rect 17693 8245 17727 8279
rect 17727 8245 17736 8279
rect 17684 8236 17736 8245
rect 17868 8236 17920 8288
rect 19892 8236 19944 8288
rect 20076 8279 20128 8288
rect 20076 8245 20085 8279
rect 20085 8245 20119 8279
rect 20119 8245 20128 8279
rect 20076 8236 20128 8245
rect 20352 8236 20404 8288
rect 20536 8236 20588 8288
rect 20720 8236 20772 8288
rect 21088 8236 21140 8288
rect 21640 8279 21692 8288
rect 21640 8245 21649 8279
rect 21649 8245 21683 8279
rect 21683 8245 21692 8279
rect 21640 8236 21692 8245
rect 21916 8236 21968 8288
rect 4366 8134 4418 8186
rect 4430 8134 4482 8186
rect 4494 8134 4546 8186
rect 4558 8134 4610 8186
rect 4622 8134 4674 8186
rect 4686 8134 4738 8186
rect 10366 8134 10418 8186
rect 10430 8134 10482 8186
rect 10494 8134 10546 8186
rect 10558 8134 10610 8186
rect 10622 8134 10674 8186
rect 10686 8134 10738 8186
rect 16366 8134 16418 8186
rect 16430 8134 16482 8186
rect 16494 8134 16546 8186
rect 16558 8134 16610 8186
rect 16622 8134 16674 8186
rect 16686 8134 16738 8186
rect 22366 8134 22418 8186
rect 22430 8134 22482 8186
rect 22494 8134 22546 8186
rect 22558 8134 22610 8186
rect 22622 8134 22674 8186
rect 22686 8134 22738 8186
rect 1768 8032 1820 8084
rect 2228 8032 2280 8084
rect 1124 7896 1176 7948
rect 1860 7939 1912 7948
rect 1860 7905 1869 7939
rect 1869 7905 1903 7939
rect 1903 7905 1912 7939
rect 1860 7896 1912 7905
rect 2136 7939 2188 7948
rect 2136 7905 2145 7939
rect 2145 7905 2179 7939
rect 2179 7905 2188 7939
rect 2136 7896 2188 7905
rect 1308 7871 1360 7880
rect 1308 7837 1317 7871
rect 1317 7837 1351 7871
rect 1351 7837 1360 7871
rect 1308 7828 1360 7837
rect 2136 7760 2188 7812
rect 848 7735 900 7744
rect 848 7701 857 7735
rect 857 7701 891 7735
rect 891 7701 900 7735
rect 848 7692 900 7701
rect 1032 7692 1084 7744
rect 2504 7939 2556 7948
rect 2504 7905 2513 7939
rect 2513 7905 2547 7939
rect 2547 7905 2556 7939
rect 2504 7896 2556 7905
rect 2688 7939 2740 7948
rect 2688 7905 2697 7939
rect 2697 7905 2731 7939
rect 2731 7905 2740 7939
rect 2688 7896 2740 7905
rect 2780 7939 2832 7948
rect 2780 7905 2789 7939
rect 2789 7905 2823 7939
rect 2823 7905 2832 7939
rect 2780 7896 2832 7905
rect 2872 7939 2924 7948
rect 2872 7905 2881 7939
rect 2881 7905 2915 7939
rect 2915 7905 2924 7939
rect 2872 7896 2924 7905
rect 3424 7964 3476 8016
rect 3976 7964 4028 8016
rect 3148 7939 3200 7948
rect 3148 7905 3157 7939
rect 3157 7905 3191 7939
rect 3191 7905 3200 7939
rect 3148 7896 3200 7905
rect 3332 7896 3384 7948
rect 3608 7939 3660 7948
rect 3608 7905 3617 7939
rect 3617 7905 3651 7939
rect 3651 7905 3660 7939
rect 3608 7896 3660 7905
rect 4896 7964 4948 8016
rect 5816 7896 5868 7948
rect 6276 7896 6328 7948
rect 6368 7939 6420 7948
rect 6368 7905 6377 7939
rect 6377 7905 6411 7939
rect 6411 7905 6420 7939
rect 6368 7896 6420 7905
rect 6552 7964 6604 8016
rect 8852 8032 8904 8084
rect 9036 8032 9088 8084
rect 9220 8032 9272 8084
rect 6828 7964 6880 8016
rect 6920 7939 6972 7948
rect 6920 7905 6929 7939
rect 6929 7905 6963 7939
rect 6963 7905 6972 7939
rect 6920 7896 6972 7905
rect 7196 7896 7248 7948
rect 2964 7828 3016 7880
rect 4804 7828 4856 7880
rect 7564 7939 7616 7948
rect 7564 7905 7573 7939
rect 7573 7905 7607 7939
rect 7607 7905 7616 7939
rect 7564 7896 7616 7905
rect 7840 7939 7892 7948
rect 7840 7905 7849 7939
rect 7849 7905 7883 7939
rect 7883 7905 7892 7939
rect 7840 7896 7892 7905
rect 3056 7760 3108 7812
rect 5080 7760 5132 7812
rect 3424 7692 3476 7744
rect 7196 7760 7248 7812
rect 7932 7760 7984 7812
rect 8944 7828 8996 7880
rect 9220 7939 9272 7948
rect 9220 7905 9229 7939
rect 9229 7905 9263 7939
rect 9263 7905 9272 7939
rect 9220 7896 9272 7905
rect 9404 7896 9456 7948
rect 9496 7871 9548 7880
rect 9496 7837 9505 7871
rect 9505 7837 9539 7871
rect 9539 7837 9548 7871
rect 9496 7828 9548 7837
rect 10508 8032 10560 8084
rect 11704 8032 11756 8084
rect 9772 7896 9824 7948
rect 11796 7964 11848 8016
rect 12440 8032 12492 8084
rect 12808 8032 12860 8084
rect 12164 8007 12216 8016
rect 12164 7973 12173 8007
rect 12173 7973 12207 8007
rect 12207 7973 12216 8007
rect 12164 7964 12216 7973
rect 15292 8032 15344 8084
rect 17868 7964 17920 8016
rect 10324 7939 10376 7948
rect 10324 7905 10333 7939
rect 10333 7905 10367 7939
rect 10367 7905 10376 7939
rect 10324 7896 10376 7905
rect 10508 7939 10560 7948
rect 10508 7905 10517 7939
rect 10517 7905 10551 7939
rect 10551 7905 10560 7939
rect 10508 7896 10560 7905
rect 10876 7828 10928 7880
rect 11060 7828 11112 7880
rect 6276 7735 6328 7744
rect 6276 7701 6285 7735
rect 6285 7701 6319 7735
rect 6319 7701 6328 7735
rect 6276 7692 6328 7701
rect 7472 7735 7524 7744
rect 7472 7701 7481 7735
rect 7481 7701 7515 7735
rect 7515 7701 7524 7735
rect 7472 7692 7524 7701
rect 7564 7692 7616 7744
rect 9128 7760 9180 7812
rect 9588 7760 9640 7812
rect 11336 7871 11388 7880
rect 11336 7837 11345 7871
rect 11345 7837 11379 7871
rect 11379 7837 11388 7871
rect 11336 7828 11388 7837
rect 11888 7896 11940 7948
rect 13544 7896 13596 7948
rect 15660 7939 15712 7948
rect 15660 7905 15669 7939
rect 15669 7905 15703 7939
rect 15703 7905 15712 7939
rect 15660 7896 15712 7905
rect 16028 7896 16080 7948
rect 17224 7896 17276 7948
rect 17960 7896 18012 7948
rect 11704 7828 11756 7880
rect 14832 7828 14884 7880
rect 17040 7828 17092 7880
rect 11152 7760 11204 7812
rect 14096 7760 14148 7812
rect 15108 7760 15160 7812
rect 15660 7760 15712 7812
rect 19156 8007 19208 8016
rect 19156 7973 19165 8007
rect 19165 7973 19199 8007
rect 19199 7973 19208 8007
rect 19156 7964 19208 7973
rect 20168 8032 20220 8084
rect 20536 8032 20588 8084
rect 20720 7964 20772 8016
rect 21180 7964 21232 8016
rect 18696 7939 18748 7948
rect 18696 7905 18705 7939
rect 18705 7905 18739 7939
rect 18739 7905 18748 7939
rect 18696 7896 18748 7905
rect 18880 7896 18932 7948
rect 18420 7871 18472 7880
rect 18420 7837 18429 7871
rect 18429 7837 18463 7871
rect 18463 7837 18472 7871
rect 18420 7828 18472 7837
rect 19616 7896 19668 7948
rect 19708 7939 19760 7948
rect 19708 7905 19717 7939
rect 19717 7905 19751 7939
rect 19751 7905 19760 7939
rect 19708 7896 19760 7905
rect 21916 7896 21968 7948
rect 20076 7760 20128 7812
rect 8208 7692 8260 7744
rect 9404 7735 9456 7744
rect 9404 7701 9413 7735
rect 9413 7701 9447 7735
rect 9447 7701 9456 7735
rect 9404 7692 9456 7701
rect 9680 7735 9732 7744
rect 9680 7701 9689 7735
rect 9689 7701 9723 7735
rect 9723 7701 9732 7735
rect 9680 7692 9732 7701
rect 11060 7692 11112 7744
rect 11796 7692 11848 7744
rect 14556 7692 14608 7744
rect 14740 7735 14792 7744
rect 14740 7701 14749 7735
rect 14749 7701 14783 7735
rect 14783 7701 14792 7735
rect 14740 7692 14792 7701
rect 14832 7735 14884 7744
rect 14832 7701 14841 7735
rect 14841 7701 14875 7735
rect 14875 7701 14884 7735
rect 14832 7692 14884 7701
rect 15292 7692 15344 7744
rect 15752 7692 15804 7744
rect 15844 7692 15896 7744
rect 17960 7735 18012 7744
rect 17960 7701 17969 7735
rect 17969 7701 18003 7735
rect 18003 7701 18012 7735
rect 17960 7692 18012 7701
rect 18788 7735 18840 7744
rect 18788 7701 18797 7735
rect 18797 7701 18831 7735
rect 18831 7701 18840 7735
rect 18788 7692 18840 7701
rect 18880 7692 18932 7744
rect 19892 7692 19944 7744
rect 20168 7692 20220 7744
rect 20996 7692 21048 7744
rect 22284 7692 22336 7744
rect 1366 7590 1418 7642
rect 1430 7590 1482 7642
rect 1494 7590 1546 7642
rect 1558 7590 1610 7642
rect 1622 7590 1674 7642
rect 1686 7590 1738 7642
rect 7366 7590 7418 7642
rect 7430 7590 7482 7642
rect 7494 7590 7546 7642
rect 7558 7590 7610 7642
rect 7622 7590 7674 7642
rect 7686 7590 7738 7642
rect 13366 7590 13418 7642
rect 13430 7590 13482 7642
rect 13494 7590 13546 7642
rect 13558 7590 13610 7642
rect 13622 7590 13674 7642
rect 13686 7590 13738 7642
rect 19366 7590 19418 7642
rect 19430 7590 19482 7642
rect 19494 7590 19546 7642
rect 19558 7590 19610 7642
rect 19622 7590 19674 7642
rect 19686 7590 19738 7642
rect 1952 7488 2004 7540
rect 2504 7488 2556 7540
rect 6736 7488 6788 7540
rect 7196 7531 7248 7540
rect 7196 7497 7205 7531
rect 7205 7497 7239 7531
rect 7239 7497 7248 7531
rect 7196 7488 7248 7497
rect 8392 7488 8444 7540
rect 10508 7488 10560 7540
rect 10876 7488 10928 7540
rect 11612 7488 11664 7540
rect 3332 7420 3384 7472
rect 5172 7420 5224 7472
rect 6920 7463 6972 7472
rect 6920 7429 6929 7463
rect 6929 7429 6963 7463
rect 6963 7429 6972 7463
rect 6920 7420 6972 7429
rect 9128 7420 9180 7472
rect 15844 7488 15896 7540
rect 16672 7488 16724 7540
rect 17132 7488 17184 7540
rect 19800 7488 19852 7540
rect 1768 7395 1820 7404
rect 1768 7361 1777 7395
rect 1777 7361 1811 7395
rect 1811 7361 1820 7395
rect 1768 7352 1820 7361
rect 2964 7352 3016 7404
rect 3148 7352 3200 7404
rect 1124 7284 1176 7336
rect 1492 7327 1544 7336
rect 1492 7293 1501 7327
rect 1501 7293 1535 7327
rect 1535 7293 1544 7327
rect 1492 7284 1544 7293
rect 3424 7352 3476 7404
rect 3608 7395 3660 7404
rect 3608 7361 3617 7395
rect 3617 7361 3651 7395
rect 3651 7361 3660 7395
rect 3608 7352 3660 7361
rect 3884 7352 3936 7404
rect 6092 7352 6144 7404
rect 2136 7216 2188 7268
rect 1860 7148 1912 7200
rect 4252 7284 4304 7336
rect 4896 7284 4948 7336
rect 5356 7284 5408 7336
rect 5816 7284 5868 7336
rect 6000 7327 6052 7336
rect 6000 7293 6009 7327
rect 6009 7293 6043 7327
rect 6043 7293 6052 7327
rect 6000 7284 6052 7293
rect 7196 7352 7248 7404
rect 7748 7395 7800 7404
rect 7748 7361 7757 7395
rect 7757 7361 7791 7395
rect 7791 7361 7800 7395
rect 7748 7352 7800 7361
rect 6736 7327 6788 7336
rect 6736 7293 6745 7327
rect 6745 7293 6779 7327
rect 6779 7293 6788 7327
rect 6736 7284 6788 7293
rect 4804 7148 4856 7200
rect 5172 7148 5224 7200
rect 5724 7191 5776 7200
rect 5724 7157 5733 7191
rect 5733 7157 5767 7191
rect 5767 7157 5776 7191
rect 5724 7148 5776 7157
rect 6828 7216 6880 7268
rect 7288 7327 7340 7336
rect 7288 7293 7297 7327
rect 7297 7293 7331 7327
rect 7331 7293 7340 7327
rect 7288 7284 7340 7293
rect 7104 7216 7156 7268
rect 7656 7284 7708 7336
rect 8392 7327 8444 7336
rect 8392 7293 8401 7327
rect 8401 7293 8435 7327
rect 8435 7293 8444 7327
rect 8392 7284 8444 7293
rect 9680 7352 9732 7404
rect 9772 7352 9824 7404
rect 10968 7352 11020 7404
rect 8116 7216 8168 7268
rect 6552 7191 6604 7200
rect 6552 7157 6561 7191
rect 6561 7157 6595 7191
rect 6595 7157 6604 7191
rect 6552 7148 6604 7157
rect 7196 7148 7248 7200
rect 7472 7148 7524 7200
rect 9220 7284 9272 7336
rect 10048 7284 10100 7336
rect 11520 7395 11572 7404
rect 11520 7361 11529 7395
rect 11529 7361 11563 7395
rect 11563 7361 11572 7395
rect 11520 7352 11572 7361
rect 11612 7352 11664 7404
rect 14740 7420 14792 7472
rect 18696 7420 18748 7472
rect 21456 7488 21508 7540
rect 21548 7488 21600 7540
rect 12992 7352 13044 7404
rect 14464 7352 14516 7404
rect 10140 7216 10192 7268
rect 11796 7284 11848 7336
rect 9128 7148 9180 7200
rect 11704 7216 11756 7268
rect 13636 7327 13688 7336
rect 13636 7293 13645 7327
rect 13645 7293 13679 7327
rect 13679 7293 13688 7327
rect 13636 7284 13688 7293
rect 11796 7148 11848 7200
rect 11888 7148 11940 7200
rect 14188 7284 14240 7336
rect 17684 7352 17736 7404
rect 20168 7420 20220 7472
rect 21732 7420 21784 7472
rect 14924 7284 14976 7336
rect 15476 7327 15528 7336
rect 15476 7293 15485 7327
rect 15485 7293 15519 7327
rect 15519 7293 15528 7327
rect 15476 7284 15528 7293
rect 16672 7284 16724 7336
rect 19616 7327 19668 7336
rect 19616 7293 19625 7327
rect 19625 7293 19659 7327
rect 19659 7293 19668 7327
rect 19616 7284 19668 7293
rect 20076 7352 20128 7404
rect 22284 7395 22336 7404
rect 22284 7361 22293 7395
rect 22293 7361 22327 7395
rect 22327 7361 22336 7395
rect 22284 7352 22336 7361
rect 14096 7191 14148 7200
rect 14096 7157 14105 7191
rect 14105 7157 14139 7191
rect 14139 7157 14148 7191
rect 14096 7148 14148 7157
rect 14188 7191 14240 7200
rect 14188 7157 14197 7191
rect 14197 7157 14231 7191
rect 14231 7157 14240 7191
rect 14188 7148 14240 7157
rect 14648 7148 14700 7200
rect 15016 7148 15068 7200
rect 19800 7216 19852 7268
rect 21824 7284 21876 7336
rect 21916 7327 21968 7336
rect 21916 7293 21925 7327
rect 21925 7293 21959 7327
rect 21959 7293 21968 7327
rect 21916 7284 21968 7293
rect 21456 7259 21508 7268
rect 21456 7225 21465 7259
rect 21465 7225 21499 7259
rect 21499 7225 21508 7259
rect 21456 7216 21508 7225
rect 21640 7259 21692 7268
rect 21640 7225 21665 7259
rect 21665 7225 21692 7259
rect 21640 7216 21692 7225
rect 22100 7216 22152 7268
rect 16856 7148 16908 7200
rect 20168 7148 20220 7200
rect 21548 7148 21600 7200
rect 4366 7046 4418 7098
rect 4430 7046 4482 7098
rect 4494 7046 4546 7098
rect 4558 7046 4610 7098
rect 4622 7046 4674 7098
rect 4686 7046 4738 7098
rect 10366 7046 10418 7098
rect 10430 7046 10482 7098
rect 10494 7046 10546 7098
rect 10558 7046 10610 7098
rect 10622 7046 10674 7098
rect 10686 7046 10738 7098
rect 16366 7046 16418 7098
rect 16430 7046 16482 7098
rect 16494 7046 16546 7098
rect 16558 7046 16610 7098
rect 16622 7046 16674 7098
rect 16686 7046 16738 7098
rect 22366 7046 22418 7098
rect 22430 7046 22482 7098
rect 22494 7046 22546 7098
rect 22558 7046 22610 7098
rect 22622 7046 22674 7098
rect 22686 7046 22738 7098
rect 1492 6944 1544 6996
rect 1768 6944 1820 6996
rect 1124 6783 1176 6792
rect 1124 6749 1133 6783
rect 1133 6749 1167 6783
rect 1167 6749 1176 6783
rect 1124 6740 1176 6749
rect 1768 6808 1820 6860
rect 1860 6851 1912 6860
rect 1860 6817 1869 6851
rect 1869 6817 1903 6851
rect 1903 6817 1912 6851
rect 1860 6808 1912 6817
rect 2136 6851 2188 6860
rect 2136 6817 2145 6851
rect 2145 6817 2179 6851
rect 2179 6817 2188 6851
rect 2136 6808 2188 6817
rect 4068 6944 4120 6996
rect 4436 6944 4488 6996
rect 5816 6944 5868 6996
rect 6000 6944 6052 6996
rect 6276 6987 6328 6996
rect 6276 6953 6285 6987
rect 6285 6953 6319 6987
rect 6319 6953 6328 6987
rect 6276 6944 6328 6953
rect 7748 6944 7800 6996
rect 2504 6851 2556 6860
rect 2504 6817 2513 6851
rect 2513 6817 2547 6851
rect 2547 6817 2556 6851
rect 2964 6876 3016 6928
rect 2504 6808 2556 6817
rect 2688 6808 2740 6860
rect 3516 6851 3568 6860
rect 3516 6817 3525 6851
rect 3525 6817 3559 6851
rect 3559 6817 3568 6851
rect 3516 6808 3568 6817
rect 3700 6851 3752 6860
rect 3700 6817 3709 6851
rect 3709 6817 3743 6851
rect 3743 6817 3752 6851
rect 3700 6808 3752 6817
rect 4252 6851 4304 6860
rect 4252 6817 4261 6851
rect 4261 6817 4295 6851
rect 4295 6817 4304 6851
rect 4252 6808 4304 6817
rect 3056 6740 3108 6792
rect 2780 6672 2832 6724
rect 4896 6876 4948 6928
rect 7472 6876 7524 6928
rect 4436 6851 4488 6860
rect 4436 6817 4445 6851
rect 4445 6817 4479 6851
rect 4479 6817 4488 6851
rect 4436 6808 4488 6817
rect 4804 6851 4856 6860
rect 4804 6817 4813 6851
rect 4813 6817 4847 6851
rect 4847 6817 4856 6851
rect 4804 6808 4856 6817
rect 5540 6851 5592 6860
rect 5540 6817 5549 6851
rect 5549 6817 5583 6851
rect 5583 6817 5592 6851
rect 5540 6808 5592 6817
rect 6184 6808 6236 6860
rect 7196 6808 7248 6860
rect 6920 6740 6972 6792
rect 8116 6808 8168 6860
rect 8852 6876 8904 6928
rect 9864 6944 9916 6996
rect 10232 6944 10284 6996
rect 11612 6944 11664 6996
rect 11704 6944 11756 6996
rect 11888 6876 11940 6928
rect 9036 6808 9088 6860
rect 9312 6808 9364 6860
rect 9588 6851 9640 6860
rect 9588 6817 9597 6851
rect 9597 6817 9631 6851
rect 9631 6817 9640 6851
rect 9588 6808 9640 6817
rect 9772 6851 9824 6860
rect 9772 6817 9781 6851
rect 9781 6817 9815 6851
rect 9815 6817 9824 6851
rect 9772 6808 9824 6817
rect 6368 6672 6420 6724
rect 6460 6715 6512 6724
rect 6460 6681 6469 6715
rect 6469 6681 6503 6715
rect 6503 6681 6512 6715
rect 6460 6672 6512 6681
rect 6552 6672 6604 6724
rect 8760 6783 8812 6792
rect 8760 6749 8769 6783
rect 8769 6749 8803 6783
rect 8803 6749 8812 6783
rect 8760 6740 8812 6749
rect 10324 6808 10376 6860
rect 10416 6851 10468 6860
rect 10416 6817 10425 6851
rect 10425 6817 10459 6851
rect 10459 6817 10468 6851
rect 10416 6808 10468 6817
rect 10692 6808 10744 6860
rect 11152 6851 11204 6860
rect 11152 6817 11161 6851
rect 11161 6817 11195 6851
rect 11195 6817 11204 6851
rect 11152 6808 11204 6817
rect 11244 6851 11296 6860
rect 11244 6817 11253 6851
rect 11253 6817 11287 6851
rect 11287 6817 11296 6851
rect 11244 6808 11296 6817
rect 10508 6740 10560 6792
rect 11428 6740 11480 6792
rect 11612 6808 11664 6860
rect 12532 6944 12584 6996
rect 13084 6944 13136 6996
rect 14740 6944 14792 6996
rect 17224 6944 17276 6996
rect 19800 6944 19852 6996
rect 20260 6944 20312 6996
rect 21548 6944 21600 6996
rect 15660 6876 15712 6928
rect 11704 6740 11756 6792
rect 12808 6783 12860 6792
rect 12808 6749 12817 6783
rect 12817 6749 12851 6783
rect 12851 6749 12860 6783
rect 12808 6740 12860 6749
rect 4528 6604 4580 6656
rect 5448 6604 5500 6656
rect 5908 6647 5960 6656
rect 5908 6613 5917 6647
rect 5917 6613 5951 6647
rect 5951 6613 5960 6647
rect 5908 6604 5960 6613
rect 7196 6604 7248 6656
rect 7748 6604 7800 6656
rect 8392 6604 8444 6656
rect 8668 6604 8720 6656
rect 11520 6672 11572 6724
rect 13084 6808 13136 6860
rect 14096 6808 14148 6860
rect 14188 6851 14240 6860
rect 14188 6817 14197 6851
rect 14197 6817 14231 6851
rect 14231 6817 14240 6851
rect 14188 6808 14240 6817
rect 14372 6851 14424 6860
rect 14372 6817 14381 6851
rect 14381 6817 14415 6851
rect 14415 6817 14424 6851
rect 14372 6808 14424 6817
rect 14464 6808 14516 6860
rect 14648 6851 14700 6860
rect 14648 6817 14657 6851
rect 14657 6817 14691 6851
rect 14691 6817 14700 6851
rect 14648 6808 14700 6817
rect 13912 6783 13964 6792
rect 13912 6749 13921 6783
rect 13921 6749 13955 6783
rect 13955 6749 13964 6783
rect 13912 6740 13964 6749
rect 15016 6783 15068 6792
rect 15016 6749 15025 6783
rect 15025 6749 15059 6783
rect 15059 6749 15068 6783
rect 15016 6740 15068 6749
rect 15200 6851 15252 6860
rect 15200 6817 15209 6851
rect 15209 6817 15243 6851
rect 15243 6817 15252 6851
rect 15200 6808 15252 6817
rect 15292 6851 15344 6860
rect 15292 6817 15301 6851
rect 15301 6817 15335 6851
rect 15335 6817 15344 6851
rect 15292 6808 15344 6817
rect 15384 6851 15436 6860
rect 15384 6817 15393 6851
rect 15393 6817 15427 6851
rect 15427 6817 15436 6851
rect 15384 6808 15436 6817
rect 15476 6808 15528 6860
rect 17040 6851 17092 6860
rect 17040 6817 17049 6851
rect 17049 6817 17083 6851
rect 17083 6817 17092 6851
rect 17040 6808 17092 6817
rect 17316 6851 17368 6860
rect 17316 6817 17325 6851
rect 17325 6817 17359 6851
rect 17359 6817 17368 6851
rect 17316 6808 17368 6817
rect 17408 6851 17460 6860
rect 17408 6817 17417 6851
rect 17417 6817 17451 6851
rect 17451 6817 17460 6851
rect 17408 6808 17460 6817
rect 17500 6851 17552 6860
rect 17500 6817 17509 6851
rect 17509 6817 17543 6851
rect 17543 6817 17552 6851
rect 17500 6808 17552 6817
rect 18236 6851 18288 6860
rect 18236 6817 18245 6851
rect 18245 6817 18279 6851
rect 18279 6817 18288 6851
rect 18236 6808 18288 6817
rect 18328 6851 18380 6860
rect 18328 6817 18337 6851
rect 18337 6817 18371 6851
rect 18371 6817 18380 6851
rect 18328 6808 18380 6817
rect 16764 6783 16816 6792
rect 16764 6749 16773 6783
rect 16773 6749 16807 6783
rect 16807 6749 16816 6783
rect 16764 6740 16816 6749
rect 19708 6808 19760 6860
rect 19892 6876 19944 6928
rect 20260 6808 20312 6860
rect 9496 6604 9548 6656
rect 10232 6604 10284 6656
rect 11152 6604 11204 6656
rect 12808 6604 12860 6656
rect 14096 6604 14148 6656
rect 15292 6672 15344 6724
rect 14556 6647 14608 6656
rect 14556 6613 14565 6647
rect 14565 6613 14599 6647
rect 14599 6613 14608 6647
rect 14556 6604 14608 6613
rect 14924 6604 14976 6656
rect 15476 6604 15528 6656
rect 15752 6604 15804 6656
rect 16488 6672 16540 6724
rect 18512 6783 18564 6792
rect 18512 6749 18521 6783
rect 18521 6749 18555 6783
rect 18555 6749 18564 6783
rect 18512 6740 18564 6749
rect 18972 6740 19024 6792
rect 19800 6783 19852 6792
rect 19800 6749 19809 6783
rect 19809 6749 19843 6783
rect 19843 6749 19852 6783
rect 19800 6740 19852 6749
rect 20168 6783 20220 6792
rect 20168 6749 20177 6783
rect 20177 6749 20211 6783
rect 20211 6749 20220 6783
rect 20168 6740 20220 6749
rect 20536 6851 20588 6860
rect 20536 6817 20545 6851
rect 20545 6817 20579 6851
rect 20579 6817 20588 6851
rect 20536 6808 20588 6817
rect 20720 6876 20772 6928
rect 21640 6808 21692 6860
rect 22008 6808 22060 6860
rect 21916 6672 21968 6724
rect 18144 6604 18196 6656
rect 18420 6647 18472 6656
rect 18420 6613 18429 6647
rect 18429 6613 18463 6647
rect 18463 6613 18472 6647
rect 18420 6604 18472 6613
rect 18512 6604 18564 6656
rect 19892 6604 19944 6656
rect 20536 6604 20588 6656
rect 21456 6604 21508 6656
rect 21824 6604 21876 6656
rect 1366 6502 1418 6554
rect 1430 6502 1482 6554
rect 1494 6502 1546 6554
rect 1558 6502 1610 6554
rect 1622 6502 1674 6554
rect 1686 6502 1738 6554
rect 7366 6502 7418 6554
rect 7430 6502 7482 6554
rect 7494 6502 7546 6554
rect 7558 6502 7610 6554
rect 7622 6502 7674 6554
rect 7686 6502 7738 6554
rect 13366 6502 13418 6554
rect 13430 6502 13482 6554
rect 13494 6502 13546 6554
rect 13558 6502 13610 6554
rect 13622 6502 13674 6554
rect 13686 6502 13738 6554
rect 19366 6502 19418 6554
rect 19430 6502 19482 6554
rect 19494 6502 19546 6554
rect 19558 6502 19610 6554
rect 19622 6502 19674 6554
rect 19686 6502 19738 6554
rect 1768 6196 1820 6248
rect 2044 6239 2096 6248
rect 2044 6205 2053 6239
rect 2053 6205 2087 6239
rect 2087 6205 2096 6239
rect 2044 6196 2096 6205
rect 2136 6196 2188 6248
rect 2412 6196 2464 6248
rect 3700 6400 3752 6452
rect 5724 6400 5776 6452
rect 5816 6443 5868 6452
rect 5816 6409 5825 6443
rect 5825 6409 5859 6443
rect 5859 6409 5868 6443
rect 5816 6400 5868 6409
rect 5908 6400 5960 6452
rect 8852 6400 8904 6452
rect 9220 6400 9272 6452
rect 9588 6443 9640 6452
rect 9588 6409 9597 6443
rect 9597 6409 9631 6443
rect 9631 6409 9640 6443
rect 9588 6400 9640 6409
rect 10324 6400 10376 6452
rect 11244 6400 11296 6452
rect 12440 6400 12492 6452
rect 3516 6196 3568 6248
rect 4068 6307 4120 6316
rect 4068 6273 4077 6307
rect 4077 6273 4111 6307
rect 4111 6273 4120 6307
rect 4068 6264 4120 6273
rect 4528 6264 4580 6316
rect 7840 6332 7892 6384
rect 8300 6332 8352 6384
rect 1952 6103 2004 6112
rect 1952 6069 1961 6103
rect 1961 6069 1995 6103
rect 1995 6069 2004 6103
rect 1952 6060 2004 6069
rect 2228 6060 2280 6112
rect 2412 6060 2464 6112
rect 5448 6239 5500 6248
rect 5448 6205 5457 6239
rect 5457 6205 5491 6239
rect 5491 6205 5500 6239
rect 5448 6196 5500 6205
rect 6000 6239 6052 6248
rect 6000 6205 6009 6239
rect 6009 6205 6043 6239
rect 6043 6205 6052 6239
rect 6000 6196 6052 6205
rect 6092 6239 6144 6248
rect 6092 6205 6101 6239
rect 6101 6205 6135 6239
rect 6135 6205 6144 6239
rect 6092 6196 6144 6205
rect 6276 6239 6328 6248
rect 6276 6205 6285 6239
rect 6285 6205 6319 6239
rect 6319 6205 6328 6239
rect 6276 6196 6328 6205
rect 6828 6196 6880 6248
rect 7104 6196 7156 6248
rect 7196 6239 7248 6248
rect 7196 6205 7205 6239
rect 7205 6205 7239 6239
rect 7239 6205 7248 6239
rect 7196 6196 7248 6205
rect 7748 6196 7800 6248
rect 7840 6196 7892 6248
rect 8392 6196 8444 6248
rect 8576 6239 8628 6248
rect 8576 6205 8585 6239
rect 8585 6205 8619 6239
rect 8619 6205 8628 6239
rect 8576 6196 8628 6205
rect 8668 6239 8720 6248
rect 8668 6205 8677 6239
rect 8677 6205 8711 6239
rect 8711 6205 8720 6239
rect 8668 6196 8720 6205
rect 8852 6196 8904 6248
rect 9312 6264 9364 6316
rect 11336 6332 11388 6384
rect 14740 6332 14792 6384
rect 15016 6400 15068 6452
rect 19892 6400 19944 6452
rect 20536 6400 20588 6452
rect 9036 6239 9088 6248
rect 9036 6205 9045 6239
rect 9045 6205 9079 6239
rect 9079 6205 9088 6239
rect 9036 6196 9088 6205
rect 9220 6239 9272 6248
rect 9220 6205 9229 6239
rect 9229 6205 9263 6239
rect 9263 6205 9272 6239
rect 9220 6196 9272 6205
rect 7380 6128 7432 6180
rect 9588 6196 9640 6248
rect 12440 6264 12492 6316
rect 14924 6264 14976 6316
rect 6552 6060 6604 6112
rect 6736 6060 6788 6112
rect 8392 6103 8444 6112
rect 8392 6069 8401 6103
rect 8401 6069 8435 6103
rect 8435 6069 8444 6103
rect 8392 6060 8444 6069
rect 10416 6128 10468 6180
rect 11244 6128 11296 6180
rect 14004 6196 14056 6248
rect 14188 6239 14240 6248
rect 14188 6205 14197 6239
rect 14197 6205 14231 6239
rect 14231 6205 14240 6239
rect 14188 6196 14240 6205
rect 14372 6239 14424 6248
rect 14372 6205 14381 6239
rect 14381 6205 14415 6239
rect 14415 6205 14424 6239
rect 14372 6196 14424 6205
rect 11428 6060 11480 6112
rect 11520 6060 11572 6112
rect 13084 6128 13136 6180
rect 14648 6239 14700 6248
rect 14648 6205 14657 6239
rect 14657 6205 14691 6239
rect 14691 6205 14700 6239
rect 14648 6196 14700 6205
rect 15108 6264 15160 6316
rect 15200 6239 15252 6248
rect 15200 6205 15209 6239
rect 15209 6205 15243 6239
rect 15243 6205 15252 6239
rect 15200 6196 15252 6205
rect 15568 6239 15620 6248
rect 15568 6205 15577 6239
rect 15577 6205 15611 6239
rect 15611 6205 15620 6239
rect 15568 6196 15620 6205
rect 15936 6264 15988 6316
rect 16212 6307 16264 6316
rect 16212 6273 16221 6307
rect 16221 6273 16255 6307
rect 16255 6273 16264 6307
rect 16212 6264 16264 6273
rect 17960 6332 18012 6384
rect 18144 6332 18196 6384
rect 18328 6264 18380 6316
rect 18880 6264 18932 6316
rect 21180 6332 21232 6384
rect 15844 6239 15896 6248
rect 15844 6205 15853 6239
rect 15853 6205 15887 6239
rect 15887 6205 15896 6239
rect 15844 6196 15896 6205
rect 16304 6239 16356 6248
rect 16304 6205 16313 6239
rect 16313 6205 16347 6239
rect 16347 6205 16356 6239
rect 16304 6196 16356 6205
rect 16488 6196 16540 6248
rect 11980 6060 12032 6112
rect 14648 6060 14700 6112
rect 18788 6196 18840 6248
rect 20536 6264 20588 6316
rect 15936 6103 15988 6112
rect 15936 6069 15945 6103
rect 15945 6069 15979 6103
rect 15979 6069 15988 6103
rect 15936 6060 15988 6069
rect 17132 6103 17184 6112
rect 17132 6069 17141 6103
rect 17141 6069 17175 6103
rect 17175 6069 17184 6103
rect 17132 6060 17184 6069
rect 18512 6103 18564 6112
rect 18512 6069 18521 6103
rect 18521 6069 18555 6103
rect 18555 6069 18564 6103
rect 18512 6060 18564 6069
rect 18696 6103 18748 6112
rect 18696 6069 18705 6103
rect 18705 6069 18739 6103
rect 18739 6069 18748 6103
rect 18696 6060 18748 6069
rect 19064 6103 19116 6112
rect 19064 6069 19073 6103
rect 19073 6069 19107 6103
rect 19107 6069 19116 6103
rect 19064 6060 19116 6069
rect 19800 6060 19852 6112
rect 20168 6128 20220 6180
rect 20628 6128 20680 6180
rect 20904 6060 20956 6112
rect 21272 6060 21324 6112
rect 22192 6103 22244 6112
rect 22192 6069 22201 6103
rect 22201 6069 22235 6103
rect 22235 6069 22244 6103
rect 22192 6060 22244 6069
rect 22284 6103 22336 6112
rect 22284 6069 22293 6103
rect 22293 6069 22327 6103
rect 22327 6069 22336 6103
rect 22284 6060 22336 6069
rect 4366 5958 4418 6010
rect 4430 5958 4482 6010
rect 4494 5958 4546 6010
rect 4558 5958 4610 6010
rect 4622 5958 4674 6010
rect 4686 5958 4738 6010
rect 10366 5958 10418 6010
rect 10430 5958 10482 6010
rect 10494 5958 10546 6010
rect 10558 5958 10610 6010
rect 10622 5958 10674 6010
rect 10686 5958 10738 6010
rect 16366 5958 16418 6010
rect 16430 5958 16482 6010
rect 16494 5958 16546 6010
rect 16558 5958 16610 6010
rect 16622 5958 16674 6010
rect 16686 5958 16738 6010
rect 22366 5958 22418 6010
rect 22430 5958 22482 6010
rect 22494 5958 22546 6010
rect 22558 5958 22610 6010
rect 22622 5958 22674 6010
rect 22686 5958 22738 6010
rect 3976 5856 4028 5908
rect 4160 5856 4212 5908
rect 5172 5856 5224 5908
rect 6276 5856 6328 5908
rect 6736 5856 6788 5908
rect 7748 5856 7800 5908
rect 8852 5856 8904 5908
rect 5356 5788 5408 5840
rect 6092 5788 6144 5840
rect 7196 5788 7248 5840
rect 8116 5788 8168 5840
rect 1768 5720 1820 5772
rect 1952 5763 2004 5772
rect 1952 5729 1961 5763
rect 1961 5729 1995 5763
rect 1995 5729 2004 5763
rect 1952 5720 2004 5729
rect 2504 5720 2556 5772
rect 3792 5763 3844 5772
rect 3792 5729 3801 5763
rect 3801 5729 3835 5763
rect 3835 5729 3844 5763
rect 3792 5720 3844 5729
rect 3976 5720 4028 5772
rect 848 5652 900 5704
rect 2412 5695 2464 5704
rect 2412 5661 2421 5695
rect 2421 5661 2455 5695
rect 2455 5661 2464 5695
rect 2412 5652 2464 5661
rect 2872 5652 2924 5704
rect 4528 5720 4580 5772
rect 4620 5763 4672 5772
rect 4620 5729 4629 5763
rect 4629 5729 4663 5763
rect 4663 5729 4672 5763
rect 4620 5720 4672 5729
rect 4804 5720 4856 5772
rect 5540 5720 5592 5772
rect 5908 5720 5960 5772
rect 6460 5720 6512 5772
rect 8208 5763 8260 5772
rect 8208 5729 8217 5763
rect 8217 5729 8251 5763
rect 8251 5729 8260 5763
rect 8208 5720 8260 5729
rect 8484 5763 8536 5772
rect 8484 5729 8493 5763
rect 8493 5729 8527 5763
rect 8527 5729 8536 5763
rect 8484 5720 8536 5729
rect 12992 5856 13044 5908
rect 13084 5856 13136 5908
rect 9404 5763 9456 5772
rect 9404 5729 9413 5763
rect 9413 5729 9447 5763
rect 9447 5729 9456 5763
rect 9404 5720 9456 5729
rect 5080 5695 5132 5704
rect 5080 5661 5089 5695
rect 5089 5661 5123 5695
rect 5123 5661 5132 5695
rect 5080 5652 5132 5661
rect 1952 5584 2004 5636
rect 4344 5584 4396 5636
rect 6368 5652 6420 5704
rect 6644 5652 6696 5704
rect 7012 5652 7064 5704
rect 5540 5627 5592 5636
rect 5540 5593 5549 5627
rect 5549 5593 5583 5627
rect 5583 5593 5592 5627
rect 5540 5584 5592 5593
rect 6000 5627 6052 5636
rect 6000 5593 6009 5627
rect 6009 5593 6043 5627
rect 6043 5593 6052 5627
rect 6000 5584 6052 5593
rect 7380 5584 7432 5636
rect 3976 5559 4028 5568
rect 3976 5525 3985 5559
rect 3985 5525 4019 5559
rect 4019 5525 4028 5559
rect 3976 5516 4028 5525
rect 4252 5559 4304 5568
rect 4252 5525 4261 5559
rect 4261 5525 4295 5559
rect 4295 5525 4304 5559
rect 4252 5516 4304 5525
rect 4528 5516 4580 5568
rect 6368 5559 6420 5568
rect 6368 5525 6377 5559
rect 6377 5525 6411 5559
rect 6411 5525 6420 5559
rect 6368 5516 6420 5525
rect 6920 5516 6972 5568
rect 8116 5695 8168 5704
rect 8116 5661 8125 5695
rect 8125 5661 8159 5695
rect 8159 5661 8168 5695
rect 8116 5652 8168 5661
rect 8668 5652 8720 5704
rect 9956 5763 10008 5772
rect 9956 5729 9965 5763
rect 9965 5729 9999 5763
rect 9999 5729 10008 5763
rect 9956 5720 10008 5729
rect 10416 5763 10468 5772
rect 10416 5729 10425 5763
rect 10425 5729 10459 5763
rect 10459 5729 10468 5763
rect 10416 5720 10468 5729
rect 11336 5720 11388 5772
rect 11428 5763 11480 5772
rect 11428 5729 11437 5763
rect 11437 5729 11471 5763
rect 11471 5729 11480 5763
rect 11428 5720 11480 5729
rect 11520 5763 11572 5772
rect 11520 5729 11529 5763
rect 11529 5729 11563 5763
rect 11563 5729 11572 5763
rect 11520 5720 11572 5729
rect 11888 5720 11940 5772
rect 12072 5763 12124 5772
rect 12072 5729 12081 5763
rect 12081 5729 12115 5763
rect 12115 5729 12124 5763
rect 12072 5720 12124 5729
rect 12716 5720 12768 5772
rect 14648 5856 14700 5908
rect 15108 5856 15160 5908
rect 15844 5856 15896 5908
rect 19064 5856 19116 5908
rect 22284 5856 22336 5908
rect 14004 5720 14056 5772
rect 9772 5584 9824 5636
rect 10968 5584 11020 5636
rect 11244 5627 11296 5636
rect 11244 5593 11253 5627
rect 11253 5593 11287 5627
rect 11287 5593 11296 5627
rect 11244 5584 11296 5593
rect 11612 5584 11664 5636
rect 13268 5652 13320 5704
rect 14372 5763 14424 5772
rect 14372 5729 14381 5763
rect 14381 5729 14415 5763
rect 14415 5729 14424 5763
rect 14372 5720 14424 5729
rect 16580 5788 16632 5840
rect 16856 5831 16908 5840
rect 16856 5797 16865 5831
rect 16865 5797 16899 5831
rect 16899 5797 16908 5831
rect 16856 5788 16908 5797
rect 18696 5788 18748 5840
rect 14740 5652 14792 5704
rect 15568 5652 15620 5704
rect 18052 5763 18104 5772
rect 18052 5729 18061 5763
rect 18061 5729 18095 5763
rect 18095 5729 18104 5763
rect 18052 5720 18104 5729
rect 18420 5720 18472 5772
rect 18604 5763 18656 5772
rect 18604 5729 18613 5763
rect 18613 5729 18647 5763
rect 18647 5729 18656 5763
rect 18604 5720 18656 5729
rect 19156 5763 19208 5772
rect 19156 5729 19165 5763
rect 19165 5729 19199 5763
rect 19199 5729 19208 5763
rect 19156 5720 19208 5729
rect 19984 5788 20036 5840
rect 19432 5763 19484 5772
rect 19432 5729 19441 5763
rect 19441 5729 19475 5763
rect 19475 5729 19484 5763
rect 19432 5720 19484 5729
rect 19524 5763 19576 5772
rect 19524 5729 19533 5763
rect 19533 5729 19567 5763
rect 19567 5729 19576 5763
rect 19524 5720 19576 5729
rect 20168 5720 20220 5772
rect 21180 5788 21232 5840
rect 22192 5788 22244 5840
rect 20904 5763 20956 5772
rect 20904 5729 20913 5763
rect 20913 5729 20947 5763
rect 20947 5729 20956 5763
rect 20904 5720 20956 5729
rect 21456 5720 21508 5772
rect 21640 5720 21692 5772
rect 14372 5584 14424 5636
rect 17132 5584 17184 5636
rect 18604 5584 18656 5636
rect 20260 5652 20312 5704
rect 20720 5584 20772 5636
rect 8576 5559 8628 5568
rect 8576 5525 8585 5559
rect 8585 5525 8619 5559
rect 8619 5525 8628 5559
rect 8576 5516 8628 5525
rect 8852 5559 8904 5568
rect 8852 5525 8861 5559
rect 8861 5525 8895 5559
rect 8895 5525 8904 5559
rect 8852 5516 8904 5525
rect 8944 5516 8996 5568
rect 10140 5516 10192 5568
rect 10784 5559 10836 5568
rect 10784 5525 10793 5559
rect 10793 5525 10827 5559
rect 10827 5525 10836 5559
rect 10784 5516 10836 5525
rect 11704 5559 11756 5568
rect 11704 5525 11713 5559
rect 11713 5525 11747 5559
rect 11747 5525 11756 5559
rect 11704 5516 11756 5525
rect 13912 5516 13964 5568
rect 14464 5516 14516 5568
rect 15200 5516 15252 5568
rect 17224 5559 17276 5568
rect 17224 5525 17233 5559
rect 17233 5525 17267 5559
rect 17267 5525 17276 5559
rect 17224 5516 17276 5525
rect 17316 5516 17368 5568
rect 18512 5559 18564 5568
rect 18512 5525 18521 5559
rect 18521 5525 18555 5559
rect 18555 5525 18564 5559
rect 18512 5516 18564 5525
rect 18880 5559 18932 5568
rect 18880 5525 18889 5559
rect 18889 5525 18923 5559
rect 18923 5525 18932 5559
rect 18880 5516 18932 5525
rect 20352 5516 20404 5568
rect 21180 5516 21232 5568
rect 22008 5559 22060 5568
rect 22008 5525 22017 5559
rect 22017 5525 22051 5559
rect 22051 5525 22060 5559
rect 22008 5516 22060 5525
rect 1366 5414 1418 5466
rect 1430 5414 1482 5466
rect 1494 5414 1546 5466
rect 1558 5414 1610 5466
rect 1622 5414 1674 5466
rect 1686 5414 1738 5466
rect 7366 5414 7418 5466
rect 7430 5414 7482 5466
rect 7494 5414 7546 5466
rect 7558 5414 7610 5466
rect 7622 5414 7674 5466
rect 7686 5414 7738 5466
rect 13366 5414 13418 5466
rect 13430 5414 13482 5466
rect 13494 5414 13546 5466
rect 13558 5414 13610 5466
rect 13622 5414 13674 5466
rect 13686 5414 13738 5466
rect 19366 5414 19418 5466
rect 19430 5414 19482 5466
rect 19494 5414 19546 5466
rect 19558 5414 19610 5466
rect 19622 5414 19674 5466
rect 19686 5414 19738 5466
rect 1768 5312 1820 5364
rect 1860 5312 1912 5364
rect 2044 5312 2096 5364
rect 4620 5312 4672 5364
rect 8484 5312 8536 5364
rect 9956 5312 10008 5364
rect 10416 5355 10468 5364
rect 10416 5321 10425 5355
rect 10425 5321 10459 5355
rect 10459 5321 10468 5355
rect 10416 5312 10468 5321
rect 11520 5312 11572 5364
rect 11888 5355 11940 5364
rect 11888 5321 11897 5355
rect 11897 5321 11931 5355
rect 11931 5321 11940 5355
rect 11888 5312 11940 5321
rect 1676 5244 1728 5296
rect 3332 5244 3384 5296
rect 3608 5244 3660 5296
rect 1860 5176 1912 5228
rect 3792 5176 3844 5228
rect 6828 5244 6880 5296
rect 8944 5244 8996 5296
rect 1492 5151 1544 5160
rect 1492 5117 1501 5151
rect 1501 5117 1535 5151
rect 1535 5117 1544 5151
rect 1492 5108 1544 5117
rect 1676 5151 1728 5160
rect 1676 5117 1685 5151
rect 1685 5117 1719 5151
rect 1719 5117 1728 5151
rect 1676 5108 1728 5117
rect 2136 5151 2188 5160
rect 2136 5117 2145 5151
rect 2145 5117 2179 5151
rect 2179 5117 2188 5151
rect 2136 5108 2188 5117
rect 2872 5151 2924 5160
rect 2872 5117 2881 5151
rect 2881 5117 2915 5151
rect 2915 5117 2924 5151
rect 2872 5108 2924 5117
rect 2228 5040 2280 5092
rect 3976 5108 4028 5160
rect 4988 5151 5040 5160
rect 4988 5117 4997 5151
rect 4997 5117 5031 5151
rect 5031 5117 5040 5151
rect 4988 5108 5040 5117
rect 5264 5151 5316 5160
rect 5264 5117 5273 5151
rect 5273 5117 5307 5151
rect 5307 5117 5316 5151
rect 5264 5108 5316 5117
rect 5356 5108 5408 5160
rect 5448 5151 5500 5160
rect 5448 5117 5457 5151
rect 5457 5117 5491 5151
rect 5491 5117 5500 5151
rect 5448 5108 5500 5117
rect 5540 5108 5592 5160
rect 5908 5151 5960 5160
rect 5908 5117 5917 5151
rect 5917 5117 5951 5151
rect 5951 5117 5960 5151
rect 5908 5108 5960 5117
rect 1308 5015 1360 5024
rect 1308 4981 1317 5015
rect 1317 4981 1351 5015
rect 1351 4981 1360 5015
rect 1308 4972 1360 4981
rect 1676 4972 1728 5024
rect 3516 4972 3568 5024
rect 4896 4972 4948 5024
rect 5172 5015 5224 5024
rect 5172 4981 5181 5015
rect 5181 4981 5215 5015
rect 5215 4981 5224 5015
rect 5172 4972 5224 4981
rect 5356 5015 5408 5024
rect 5356 4981 5365 5015
rect 5365 4981 5399 5015
rect 5399 4981 5408 5015
rect 5356 4972 5408 4981
rect 5632 5040 5684 5092
rect 6460 5083 6512 5092
rect 6460 5049 6469 5083
rect 6469 5049 6503 5083
rect 6503 5049 6512 5083
rect 6460 5040 6512 5049
rect 5540 4972 5592 5024
rect 6184 4972 6236 5024
rect 6644 5151 6696 5160
rect 6644 5117 6653 5151
rect 6653 5117 6687 5151
rect 6687 5117 6696 5151
rect 6644 5108 6696 5117
rect 6920 5151 6972 5160
rect 6920 5117 6929 5151
rect 6929 5117 6963 5151
rect 6963 5117 6972 5151
rect 6920 5108 6972 5117
rect 7012 5151 7064 5160
rect 7012 5117 7021 5151
rect 7021 5117 7055 5151
rect 7055 5117 7064 5151
rect 7012 5108 7064 5117
rect 8576 5176 8628 5228
rect 10140 5244 10192 5296
rect 12716 5312 12768 5364
rect 12992 5312 13044 5364
rect 7656 5108 7708 5160
rect 7196 5040 7248 5092
rect 6920 4972 6972 5024
rect 8760 5108 8812 5160
rect 9128 5219 9180 5228
rect 9128 5185 9137 5219
rect 9137 5185 9171 5219
rect 9171 5185 9180 5219
rect 9128 5176 9180 5185
rect 10048 5176 10100 5228
rect 11060 5176 11112 5228
rect 12900 5244 12952 5296
rect 19064 5312 19116 5364
rect 19800 5312 19852 5364
rect 20168 5312 20220 5364
rect 20720 5312 20772 5364
rect 21456 5312 21508 5364
rect 22008 5312 22060 5364
rect 9220 5108 9272 5160
rect 11244 5151 11296 5160
rect 11244 5117 11253 5151
rect 11253 5117 11287 5151
rect 11287 5117 11296 5151
rect 11244 5108 11296 5117
rect 11336 5151 11388 5160
rect 11336 5117 11345 5151
rect 11345 5117 11379 5151
rect 11379 5117 11388 5151
rect 11336 5108 11388 5117
rect 11796 5108 11848 5160
rect 12164 5108 12216 5160
rect 12992 5176 13044 5228
rect 14096 5219 14148 5228
rect 14096 5185 14105 5219
rect 14105 5185 14139 5219
rect 14139 5185 14148 5219
rect 14096 5176 14148 5185
rect 14464 5176 14516 5228
rect 8116 5040 8168 5092
rect 9312 5040 9364 5092
rect 10140 5040 10192 5092
rect 13268 5108 13320 5160
rect 13820 5108 13872 5160
rect 14004 5151 14056 5160
rect 14004 5117 14013 5151
rect 14013 5117 14047 5151
rect 14047 5117 14056 5151
rect 14004 5108 14056 5117
rect 14188 5108 14240 5160
rect 14740 5108 14792 5160
rect 16580 5176 16632 5228
rect 16672 5219 16724 5228
rect 16672 5185 16681 5219
rect 16681 5185 16715 5219
rect 16715 5185 16724 5219
rect 16672 5176 16724 5185
rect 20260 5244 20312 5296
rect 17040 5176 17092 5228
rect 19064 5219 19116 5228
rect 19064 5185 19073 5219
rect 19073 5185 19107 5219
rect 19107 5185 19116 5219
rect 19064 5176 19116 5185
rect 7932 4972 7984 5024
rect 9772 4972 9824 5024
rect 12256 4972 12308 5024
rect 16028 5040 16080 5092
rect 17408 5151 17460 5160
rect 17408 5117 17417 5151
rect 17417 5117 17451 5151
rect 17451 5117 17460 5151
rect 17408 5108 17460 5117
rect 17592 5151 17644 5160
rect 17592 5117 17601 5151
rect 17601 5117 17635 5151
rect 17635 5117 17644 5151
rect 17592 5108 17644 5117
rect 18696 5108 18748 5160
rect 17868 5040 17920 5092
rect 12716 4972 12768 5024
rect 12992 4972 13044 5024
rect 14372 5015 14424 5024
rect 14372 4981 14381 5015
rect 14381 4981 14415 5015
rect 14415 4981 14424 5015
rect 14372 4972 14424 4981
rect 14648 5015 14700 5024
rect 14648 4981 14657 5015
rect 14657 4981 14691 5015
rect 14691 4981 14700 5015
rect 14648 4972 14700 4981
rect 16212 4972 16264 5024
rect 18236 4972 18288 5024
rect 18972 5151 19024 5160
rect 18972 5117 18981 5151
rect 18981 5117 19015 5151
rect 19015 5117 19024 5151
rect 18972 5108 19024 5117
rect 19984 5176 20036 5228
rect 22284 5176 22336 5228
rect 19064 5040 19116 5092
rect 19892 5108 19944 5160
rect 21088 5108 21140 5160
rect 21180 5151 21232 5160
rect 21180 5117 21189 5151
rect 21189 5117 21223 5151
rect 21223 5117 21232 5151
rect 21180 5108 21232 5117
rect 21548 5151 21600 5160
rect 21548 5117 21557 5151
rect 21557 5117 21591 5151
rect 21591 5117 21600 5151
rect 21548 5108 21600 5117
rect 19156 4972 19208 5024
rect 19708 4972 19760 5024
rect 19984 5015 20036 5024
rect 19984 4981 19993 5015
rect 19993 4981 20027 5015
rect 20027 4981 20036 5015
rect 19984 4972 20036 4981
rect 20628 4972 20680 5024
rect 21364 5040 21416 5092
rect 21732 5040 21784 5092
rect 4366 4870 4418 4922
rect 4430 4870 4482 4922
rect 4494 4870 4546 4922
rect 4558 4870 4610 4922
rect 4622 4870 4674 4922
rect 4686 4870 4738 4922
rect 10366 4870 10418 4922
rect 10430 4870 10482 4922
rect 10494 4870 10546 4922
rect 10558 4870 10610 4922
rect 10622 4870 10674 4922
rect 10686 4870 10738 4922
rect 16366 4870 16418 4922
rect 16430 4870 16482 4922
rect 16494 4870 16546 4922
rect 16558 4870 16610 4922
rect 16622 4870 16674 4922
rect 16686 4870 16738 4922
rect 22366 4870 22418 4922
rect 22430 4870 22482 4922
rect 22494 4870 22546 4922
rect 22558 4870 22610 4922
rect 22622 4870 22674 4922
rect 22686 4870 22738 4922
rect 1124 4811 1176 4820
rect 1124 4777 1133 4811
rect 1133 4777 1167 4811
rect 1167 4777 1176 4811
rect 1124 4768 1176 4777
rect 664 4632 716 4684
rect 1492 4700 1544 4752
rect 2320 4768 2372 4820
rect 2688 4768 2740 4820
rect 2780 4811 2832 4820
rect 2780 4777 2789 4811
rect 2789 4777 2823 4811
rect 2823 4777 2832 4811
rect 2780 4768 2832 4777
rect 3240 4768 3292 4820
rect 3516 4768 3568 4820
rect 3792 4768 3844 4820
rect 2228 4700 2280 4752
rect 4804 4768 4856 4820
rect 5264 4768 5316 4820
rect 5632 4811 5684 4820
rect 5632 4777 5641 4811
rect 5641 4777 5675 4811
rect 5675 4777 5684 4811
rect 5632 4768 5684 4777
rect 7012 4768 7064 4820
rect 9220 4811 9272 4820
rect 9220 4777 9229 4811
rect 9229 4777 9263 4811
rect 9263 4777 9272 4811
rect 9220 4768 9272 4777
rect 10140 4811 10192 4820
rect 10140 4777 10149 4811
rect 10149 4777 10183 4811
rect 10183 4777 10192 4811
rect 10140 4768 10192 4777
rect 4528 4700 4580 4752
rect 4896 4700 4948 4752
rect 1308 4675 1360 4684
rect 1308 4641 1317 4675
rect 1317 4641 1351 4675
rect 1351 4641 1360 4675
rect 1308 4632 1360 4641
rect 1124 4607 1176 4616
rect 1124 4573 1133 4607
rect 1133 4573 1167 4607
rect 1167 4573 1176 4607
rect 1124 4564 1176 4573
rect 1860 4675 1912 4684
rect 1860 4641 1869 4675
rect 1869 4641 1903 4675
rect 1903 4641 1912 4675
rect 1860 4632 1912 4641
rect 2044 4675 2096 4684
rect 2044 4641 2053 4675
rect 2053 4641 2087 4675
rect 2087 4641 2096 4675
rect 2044 4632 2096 4641
rect 2320 4675 2372 4684
rect 2320 4641 2329 4675
rect 2329 4641 2363 4675
rect 2363 4641 2372 4675
rect 2320 4632 2372 4641
rect 2964 4632 3016 4684
rect 3700 4675 3752 4684
rect 3700 4641 3709 4675
rect 3709 4641 3743 4675
rect 3743 4641 3752 4675
rect 3700 4632 3752 4641
rect 4068 4675 4120 4684
rect 4068 4641 4077 4675
rect 4077 4641 4111 4675
rect 4111 4641 4120 4675
rect 4068 4632 4120 4641
rect 4160 4675 4212 4684
rect 4160 4641 4169 4675
rect 4169 4641 4203 4675
rect 4203 4641 4212 4675
rect 4160 4632 4212 4641
rect 5724 4700 5776 4752
rect 7196 4700 7248 4752
rect 7656 4700 7708 4752
rect 9772 4700 9824 4752
rect 1768 4496 1820 4548
rect 2596 4496 2648 4548
rect 4252 4564 4304 4616
rect 4896 4564 4948 4616
rect 4988 4496 5040 4548
rect 6184 4632 6236 4684
rect 8392 4632 8444 4684
rect 8576 4675 8628 4684
rect 8576 4641 8585 4675
rect 8585 4641 8619 4675
rect 8619 4641 8628 4675
rect 12256 4768 12308 4820
rect 8576 4632 8628 4641
rect 11520 4632 11572 4684
rect 11888 4632 11940 4684
rect 12624 4700 12676 4752
rect 14004 4768 14056 4820
rect 14464 4811 14516 4820
rect 14464 4777 14473 4811
rect 14473 4777 14507 4811
rect 14507 4777 14516 4811
rect 14464 4768 14516 4777
rect 14648 4768 14700 4820
rect 17868 4768 17920 4820
rect 5356 4607 5408 4616
rect 5356 4573 5365 4607
rect 5365 4573 5399 4607
rect 5399 4573 5408 4607
rect 5356 4564 5408 4573
rect 2964 4471 3016 4480
rect 2964 4437 2973 4471
rect 2973 4437 3007 4471
rect 3007 4437 3016 4471
rect 2964 4428 3016 4437
rect 5264 4428 5316 4480
rect 6736 4564 6788 4616
rect 5908 4496 5960 4548
rect 7012 4607 7064 4616
rect 7012 4573 7021 4607
rect 7021 4573 7055 4607
rect 7055 4573 7064 4607
rect 7012 4564 7064 4573
rect 7840 4564 7892 4616
rect 8116 4564 8168 4616
rect 8300 4564 8352 4616
rect 8392 4496 8444 4548
rect 7840 4428 7892 4480
rect 9956 4564 10008 4616
rect 10232 4607 10284 4616
rect 10232 4573 10241 4607
rect 10241 4573 10275 4607
rect 10275 4573 10284 4607
rect 10232 4564 10284 4573
rect 11244 4564 11296 4616
rect 12164 4564 12216 4616
rect 12992 4675 13044 4684
rect 12992 4641 13001 4675
rect 13001 4641 13035 4675
rect 13035 4641 13044 4675
rect 12992 4632 13044 4641
rect 13176 4632 13228 4684
rect 15476 4700 15528 4752
rect 17592 4700 17644 4752
rect 18972 4768 19024 4820
rect 19708 4768 19760 4820
rect 19892 4768 19944 4820
rect 21824 4768 21876 4820
rect 21916 4768 21968 4820
rect 13912 4632 13964 4684
rect 12900 4564 12952 4616
rect 14832 4564 14884 4616
rect 16120 4675 16172 4684
rect 16120 4641 16129 4675
rect 16129 4641 16163 4675
rect 16163 4641 16172 4675
rect 16120 4632 16172 4641
rect 17224 4675 17276 4684
rect 17224 4641 17233 4675
rect 17233 4641 17267 4675
rect 17267 4641 17276 4675
rect 17224 4632 17276 4641
rect 17868 4675 17920 4684
rect 17868 4641 17877 4675
rect 17877 4641 17911 4675
rect 17911 4641 17920 4675
rect 17868 4632 17920 4641
rect 11152 4496 11204 4548
rect 8668 4428 8720 4480
rect 8944 4428 8996 4480
rect 9772 4428 9824 4480
rect 12348 4428 12400 4480
rect 13176 4496 13228 4548
rect 13268 4428 13320 4480
rect 15384 4496 15436 4548
rect 14004 4471 14056 4480
rect 14004 4437 14013 4471
rect 14013 4437 14047 4471
rect 14047 4437 14056 4471
rect 14004 4428 14056 4437
rect 14924 4471 14976 4480
rect 14924 4437 14933 4471
rect 14933 4437 14967 4471
rect 14967 4437 14976 4471
rect 14924 4428 14976 4437
rect 16212 4471 16264 4480
rect 16212 4437 16221 4471
rect 16221 4437 16255 4471
rect 16255 4437 16264 4471
rect 16212 4428 16264 4437
rect 18052 4564 18104 4616
rect 18420 4675 18472 4684
rect 18420 4641 18429 4675
rect 18429 4641 18463 4675
rect 18463 4641 18472 4675
rect 18420 4632 18472 4641
rect 18512 4675 18564 4684
rect 18512 4641 18521 4675
rect 18521 4641 18555 4675
rect 18555 4641 18564 4675
rect 18512 4632 18564 4641
rect 18880 4632 18932 4684
rect 18604 4564 18656 4616
rect 17040 4471 17092 4480
rect 17040 4437 17049 4471
rect 17049 4437 17083 4471
rect 17083 4437 17092 4471
rect 17040 4428 17092 4437
rect 18696 4496 18748 4548
rect 19800 4632 19852 4684
rect 18788 4471 18840 4480
rect 18788 4437 18797 4471
rect 18797 4437 18831 4471
rect 18831 4437 18840 4471
rect 18788 4428 18840 4437
rect 20628 4632 20680 4684
rect 21180 4700 21232 4752
rect 21088 4675 21140 4684
rect 21088 4641 21097 4675
rect 21097 4641 21131 4675
rect 21131 4641 21140 4675
rect 21088 4632 21140 4641
rect 21732 4700 21784 4752
rect 21548 4675 21600 4684
rect 21548 4641 21557 4675
rect 21557 4641 21591 4675
rect 21591 4641 21600 4675
rect 21548 4632 21600 4641
rect 21640 4675 21692 4684
rect 21640 4641 21649 4675
rect 21649 4641 21683 4675
rect 21683 4641 21692 4675
rect 21640 4632 21692 4641
rect 20444 4496 20496 4548
rect 22008 4607 22060 4616
rect 22008 4573 22017 4607
rect 22017 4573 22051 4607
rect 22051 4573 22060 4607
rect 22008 4564 22060 4573
rect 22284 4675 22336 4684
rect 22284 4641 22293 4675
rect 22293 4641 22327 4675
rect 22327 4641 22336 4675
rect 22284 4632 22336 4641
rect 23388 4564 23440 4616
rect 22284 4496 22336 4548
rect 21088 4428 21140 4480
rect 21640 4428 21692 4480
rect 22100 4428 22152 4480
rect 1366 4326 1418 4378
rect 1430 4326 1482 4378
rect 1494 4326 1546 4378
rect 1558 4326 1610 4378
rect 1622 4326 1674 4378
rect 1686 4326 1738 4378
rect 7366 4326 7418 4378
rect 7430 4326 7482 4378
rect 7494 4326 7546 4378
rect 7558 4326 7610 4378
rect 7622 4326 7674 4378
rect 7686 4326 7738 4378
rect 13366 4326 13418 4378
rect 13430 4326 13482 4378
rect 13494 4326 13546 4378
rect 13558 4326 13610 4378
rect 13622 4326 13674 4378
rect 13686 4326 13738 4378
rect 19366 4326 19418 4378
rect 19430 4326 19482 4378
rect 19494 4326 19546 4378
rect 19558 4326 19610 4378
rect 19622 4326 19674 4378
rect 19686 4326 19738 4378
rect 2320 4267 2372 4276
rect 2320 4233 2329 4267
rect 2329 4233 2363 4267
rect 2363 4233 2372 4267
rect 2320 4224 2372 4233
rect 4988 4267 5040 4276
rect 4988 4233 4997 4267
rect 4997 4233 5031 4267
rect 5031 4233 5040 4267
rect 4988 4224 5040 4233
rect 5356 4267 5408 4276
rect 5356 4233 5365 4267
rect 5365 4233 5399 4267
rect 5399 4233 5408 4267
rect 5356 4224 5408 4233
rect 7012 4224 7064 4276
rect 7656 4224 7708 4276
rect 7840 4224 7892 4276
rect 8024 4267 8076 4276
rect 8024 4233 8033 4267
rect 8033 4233 8067 4267
rect 8067 4233 8076 4267
rect 8024 4224 8076 4233
rect 8392 4267 8444 4276
rect 8392 4233 8401 4267
rect 8401 4233 8435 4267
rect 8435 4233 8444 4267
rect 8392 4224 8444 4233
rect 9680 4224 9732 4276
rect 12532 4267 12584 4276
rect 12532 4233 12541 4267
rect 12541 4233 12575 4267
rect 12575 4233 12584 4267
rect 12532 4224 12584 4233
rect 12716 4224 12768 4276
rect 3056 4156 3108 4208
rect 1676 4088 1728 4140
rect 4160 4088 4212 4140
rect 1768 4020 1820 4072
rect 2780 4020 2832 4072
rect 3424 4020 3476 4072
rect 4344 4063 4396 4072
rect 4344 4029 4353 4063
rect 4353 4029 4387 4063
rect 4387 4029 4396 4063
rect 4344 4020 4396 4029
rect 4528 4063 4580 4072
rect 4528 4029 4537 4063
rect 4537 4029 4571 4063
rect 4571 4029 4580 4063
rect 4528 4020 4580 4029
rect 4896 4063 4948 4072
rect 4896 4029 4905 4063
rect 4905 4029 4939 4063
rect 4939 4029 4948 4063
rect 4896 4020 4948 4029
rect 4988 4020 5040 4072
rect 2964 3952 3016 4004
rect 5264 4063 5316 4072
rect 5264 4029 5273 4063
rect 5273 4029 5307 4063
rect 5307 4029 5316 4063
rect 5264 4020 5316 4029
rect 5448 4020 5500 4072
rect 6092 4088 6144 4140
rect 6276 4020 6328 4072
rect 7104 4156 7156 4208
rect 9404 4156 9456 4208
rect 9588 4156 9640 4208
rect 9772 4156 9824 4208
rect 11060 4156 11112 4208
rect 11428 4156 11480 4208
rect 11796 4156 11848 4208
rect 5356 3952 5408 4004
rect 7104 4063 7156 4072
rect 7104 4029 7113 4063
rect 7113 4029 7147 4063
rect 7147 4029 7156 4063
rect 7104 4020 7156 4029
rect 8116 4088 8168 4140
rect 7656 4020 7708 4072
rect 8944 4088 8996 4140
rect 9128 4088 9180 4140
rect 8576 4063 8628 4072
rect 8576 4029 8585 4063
rect 8585 4029 8619 4063
rect 8619 4029 8628 4063
rect 8576 4020 8628 4029
rect 9312 4063 9364 4072
rect 9312 4029 9321 4063
rect 9321 4029 9355 4063
rect 9355 4029 9364 4063
rect 9312 4020 9364 4029
rect 8944 3952 8996 4004
rect 9680 4020 9732 4072
rect 10692 4063 10744 4072
rect 10692 4029 10701 4063
rect 10701 4029 10735 4063
rect 10735 4029 10744 4063
rect 10692 4020 10744 4029
rect 11336 4088 11388 4140
rect 14188 4224 14240 4276
rect 14924 4224 14976 4276
rect 21548 4224 21600 4276
rect 11244 4020 11296 4072
rect 11796 4020 11848 4072
rect 9588 3995 9640 4004
rect 9588 3961 9597 3995
rect 9597 3961 9631 3995
rect 9631 3961 9640 3995
rect 9588 3952 9640 3961
rect 10232 3995 10284 4004
rect 10232 3961 10241 3995
rect 10241 3961 10275 3995
rect 10275 3961 10284 3995
rect 10232 3952 10284 3961
rect 10784 3952 10836 4004
rect 3148 3884 3200 3936
rect 4344 3927 4396 3936
rect 4344 3893 4353 3927
rect 4353 3893 4387 3927
rect 4387 3893 4396 3927
rect 4344 3884 4396 3893
rect 6828 3884 6880 3936
rect 7472 3884 7524 3936
rect 7748 3884 7800 3936
rect 9220 3884 9272 3936
rect 9680 3884 9732 3936
rect 10140 3884 10192 3936
rect 11336 3884 11388 3936
rect 11796 3927 11848 3936
rect 11796 3893 11805 3927
rect 11805 3893 11839 3927
rect 11839 3893 11848 3927
rect 11796 3884 11848 3893
rect 11980 3884 12032 3936
rect 12440 4063 12492 4072
rect 12440 4029 12449 4063
rect 12449 4029 12483 4063
rect 12483 4029 12492 4063
rect 12440 4020 12492 4029
rect 12808 4063 12860 4072
rect 12808 4029 12817 4063
rect 12817 4029 12851 4063
rect 12851 4029 12860 4063
rect 12808 4020 12860 4029
rect 12900 4020 12952 4072
rect 13728 4020 13780 4072
rect 13820 4063 13872 4072
rect 13820 4029 13829 4063
rect 13829 4029 13863 4063
rect 13863 4029 13872 4063
rect 13820 4020 13872 4029
rect 14096 4156 14148 4208
rect 14464 4156 14516 4208
rect 14004 4088 14056 4140
rect 14740 4131 14792 4140
rect 14740 4097 14749 4131
rect 14749 4097 14783 4131
rect 14783 4097 14792 4131
rect 14740 4088 14792 4097
rect 15200 4131 15252 4140
rect 15200 4097 15209 4131
rect 15209 4097 15243 4131
rect 15243 4097 15252 4131
rect 15200 4088 15252 4097
rect 15292 4131 15344 4140
rect 15292 4097 15301 4131
rect 15301 4097 15335 4131
rect 15335 4097 15344 4131
rect 15292 4088 15344 4097
rect 15384 4131 15436 4140
rect 15384 4097 15393 4131
rect 15393 4097 15427 4131
rect 15427 4097 15436 4131
rect 15384 4088 15436 4097
rect 14188 4020 14240 4072
rect 14464 4063 14516 4072
rect 14464 4029 14473 4063
rect 14473 4029 14507 4063
rect 14507 4029 14516 4063
rect 14464 4020 14516 4029
rect 15660 4088 15712 4140
rect 16304 4131 16356 4140
rect 16304 4097 16313 4131
rect 16313 4097 16347 4131
rect 16347 4097 16356 4131
rect 16304 4088 16356 4097
rect 16396 4131 16448 4140
rect 16396 4097 16405 4131
rect 16405 4097 16439 4131
rect 16439 4097 16448 4131
rect 16396 4088 16448 4097
rect 15844 4063 15896 4072
rect 15844 4029 15853 4063
rect 15853 4029 15887 4063
rect 15887 4029 15896 4063
rect 15844 4020 15896 4029
rect 16120 4063 16172 4072
rect 16120 4029 16129 4063
rect 16129 4029 16163 4063
rect 16163 4029 16172 4063
rect 16120 4020 16172 4029
rect 12624 3952 12676 4004
rect 18052 4156 18104 4208
rect 16856 4088 16908 4140
rect 19892 4088 19944 4140
rect 19340 4063 19392 4072
rect 19340 4029 19349 4063
rect 19349 4029 19383 4063
rect 19383 4029 19392 4063
rect 19340 4020 19392 4029
rect 20260 4020 20312 4072
rect 20352 4063 20404 4072
rect 20352 4029 20361 4063
rect 20361 4029 20395 4063
rect 20395 4029 20404 4063
rect 20352 4020 20404 4029
rect 20444 4063 20496 4072
rect 20444 4029 20453 4063
rect 20453 4029 20487 4063
rect 20487 4029 20496 4063
rect 20444 4020 20496 4029
rect 20628 4063 20680 4072
rect 20628 4029 20637 4063
rect 20637 4029 20671 4063
rect 20671 4029 20680 4063
rect 20628 4020 20680 4029
rect 21088 4131 21140 4140
rect 21088 4097 21097 4131
rect 21097 4097 21131 4131
rect 21131 4097 21140 4131
rect 21088 4088 21140 4097
rect 21180 4063 21232 4072
rect 21180 4029 21189 4063
rect 21189 4029 21223 4063
rect 21223 4029 21232 4063
rect 21180 4020 21232 4029
rect 21364 4063 21416 4072
rect 21364 4029 21377 4063
rect 21377 4029 21416 4063
rect 21364 4020 21416 4029
rect 21456 4020 21508 4072
rect 21916 4020 21968 4072
rect 22008 4063 22060 4072
rect 22008 4029 22017 4063
rect 22017 4029 22051 4063
rect 22051 4029 22060 4063
rect 22008 4020 22060 4029
rect 22100 4063 22152 4072
rect 22100 4029 22109 4063
rect 22109 4029 22143 4063
rect 22143 4029 22152 4063
rect 22100 4020 22152 4029
rect 22928 4156 22980 4208
rect 12808 3884 12860 3936
rect 12992 3927 13044 3936
rect 12992 3893 13001 3927
rect 13001 3893 13035 3927
rect 13035 3893 13044 3927
rect 12992 3884 13044 3893
rect 13176 3884 13228 3936
rect 13820 3884 13872 3936
rect 14924 3927 14976 3936
rect 14924 3893 14933 3927
rect 14933 3893 14967 3927
rect 14967 3893 14976 3927
rect 14924 3884 14976 3893
rect 15108 3884 15160 3936
rect 15660 3927 15712 3936
rect 15660 3893 15669 3927
rect 15669 3893 15703 3927
rect 15703 3893 15712 3927
rect 15660 3884 15712 3893
rect 16764 3884 16816 3936
rect 19340 3884 19392 3936
rect 20076 3884 20128 3936
rect 20168 3927 20220 3936
rect 20168 3893 20177 3927
rect 20177 3893 20211 3927
rect 20211 3893 20220 3927
rect 20168 3884 20220 3893
rect 20352 3884 20404 3936
rect 20904 3927 20956 3936
rect 20904 3893 20913 3927
rect 20913 3893 20947 3927
rect 20947 3893 20956 3927
rect 20904 3884 20956 3893
rect 21180 3884 21232 3936
rect 22192 3952 22244 4004
rect 23112 4020 23164 4072
rect 23388 3952 23440 4004
rect 22836 3927 22888 3936
rect 22836 3893 22845 3927
rect 22845 3893 22879 3927
rect 22879 3893 22888 3927
rect 22836 3884 22888 3893
rect 4366 3782 4418 3834
rect 4430 3782 4482 3834
rect 4494 3782 4546 3834
rect 4558 3782 4610 3834
rect 4622 3782 4674 3834
rect 4686 3782 4738 3834
rect 10366 3782 10418 3834
rect 10430 3782 10482 3834
rect 10494 3782 10546 3834
rect 10558 3782 10610 3834
rect 10622 3782 10674 3834
rect 10686 3782 10738 3834
rect 16366 3782 16418 3834
rect 16430 3782 16482 3834
rect 16494 3782 16546 3834
rect 16558 3782 16610 3834
rect 16622 3782 16674 3834
rect 16686 3782 16738 3834
rect 22366 3782 22418 3834
rect 22430 3782 22482 3834
rect 22494 3782 22546 3834
rect 22558 3782 22610 3834
rect 22622 3782 22674 3834
rect 22686 3782 22738 3834
rect 1676 3723 1728 3732
rect 1676 3689 1685 3723
rect 1685 3689 1719 3723
rect 1719 3689 1728 3723
rect 1676 3680 1728 3689
rect 1216 3655 1268 3664
rect 1216 3621 1225 3655
rect 1225 3621 1259 3655
rect 1259 3621 1268 3655
rect 1216 3612 1268 3621
rect 6092 3655 6144 3664
rect 6092 3621 6101 3655
rect 6101 3621 6135 3655
rect 6135 3621 6144 3655
rect 6092 3612 6144 3621
rect 6184 3612 6236 3664
rect 3148 3587 3200 3596
rect 3148 3553 3157 3587
rect 3157 3553 3191 3587
rect 3191 3553 3200 3587
rect 3148 3544 3200 3553
rect 4252 3544 4304 3596
rect 5172 3544 5224 3596
rect 6276 3587 6328 3596
rect 6276 3553 6285 3587
rect 6285 3553 6319 3587
rect 6319 3553 6328 3587
rect 6276 3544 6328 3553
rect 7932 3680 7984 3732
rect 8852 3680 8904 3732
rect 7840 3612 7892 3664
rect 7288 3544 7340 3596
rect 8300 3544 8352 3596
rect 3056 3519 3108 3528
rect 3056 3485 3065 3519
rect 3065 3485 3099 3519
rect 3099 3485 3108 3519
rect 3056 3476 3108 3485
rect 8760 3544 8812 3596
rect 8944 3587 8996 3596
rect 8944 3553 8953 3587
rect 8953 3553 8987 3587
rect 8987 3553 8996 3587
rect 8944 3544 8996 3553
rect 9588 3680 9640 3732
rect 9312 3544 9364 3596
rect 9680 3612 9732 3664
rect 9772 3612 9824 3664
rect 9496 3544 9548 3596
rect 9772 3519 9824 3528
rect 9772 3485 9781 3519
rect 9781 3485 9815 3519
rect 9815 3485 9824 3519
rect 9772 3476 9824 3485
rect 10232 3680 10284 3732
rect 10140 3544 10192 3596
rect 10508 3587 10560 3596
rect 10508 3553 10517 3587
rect 10517 3553 10551 3587
rect 10551 3553 10560 3587
rect 10508 3544 10560 3553
rect 10968 3544 11020 3596
rect 11336 3587 11388 3596
rect 11336 3553 11345 3587
rect 11345 3553 11379 3587
rect 11379 3553 11388 3587
rect 11336 3544 11388 3553
rect 1124 3408 1176 3460
rect 9312 3408 9364 3460
rect 9496 3408 9548 3460
rect 10600 3519 10652 3528
rect 10600 3485 10609 3519
rect 10609 3485 10643 3519
rect 10643 3485 10652 3519
rect 10600 3476 10652 3485
rect 10692 3519 10744 3528
rect 10692 3485 10701 3519
rect 10701 3485 10735 3519
rect 10735 3485 10744 3519
rect 10692 3476 10744 3485
rect 10784 3476 10836 3528
rect 11428 3519 11480 3528
rect 11428 3485 11437 3519
rect 11437 3485 11471 3519
rect 11471 3485 11480 3519
rect 11428 3476 11480 3485
rect 12624 3612 12676 3664
rect 11888 3544 11940 3596
rect 12072 3587 12124 3596
rect 12072 3553 12081 3587
rect 12081 3553 12115 3587
rect 12115 3553 12124 3587
rect 12072 3544 12124 3553
rect 12348 3587 12400 3596
rect 12348 3553 12357 3587
rect 12357 3553 12391 3587
rect 12391 3553 12400 3587
rect 12348 3544 12400 3553
rect 12440 3476 12492 3528
rect 12900 3680 12952 3732
rect 14740 3680 14792 3732
rect 14832 3680 14884 3732
rect 16120 3680 16172 3732
rect 16672 3680 16724 3732
rect 15660 3612 15712 3664
rect 19800 3680 19852 3732
rect 12808 3408 12860 3460
rect 13820 3587 13872 3596
rect 13820 3553 13829 3587
rect 13829 3553 13863 3587
rect 13863 3553 13872 3587
rect 13820 3544 13872 3553
rect 14096 3587 14148 3596
rect 14096 3553 14105 3587
rect 14105 3553 14139 3587
rect 14139 3553 14148 3587
rect 14096 3544 14148 3553
rect 15936 3544 15988 3596
rect 13268 3476 13320 3528
rect 15384 3476 15436 3528
rect 15844 3476 15896 3528
rect 16672 3587 16724 3596
rect 16672 3553 16681 3587
rect 16681 3553 16715 3587
rect 16715 3553 16724 3587
rect 16672 3544 16724 3553
rect 17960 3612 18012 3664
rect 18880 3612 18932 3664
rect 20168 3612 20220 3664
rect 21364 3680 21416 3732
rect 19524 3587 19576 3596
rect 19524 3553 19533 3587
rect 19533 3553 19567 3587
rect 19567 3553 19576 3587
rect 19524 3544 19576 3553
rect 19800 3544 19852 3596
rect 19892 3587 19944 3596
rect 19892 3553 19901 3587
rect 19901 3553 19935 3587
rect 19935 3553 19944 3587
rect 19892 3544 19944 3553
rect 20904 3544 20956 3596
rect 18512 3476 18564 3528
rect 18880 3519 18932 3528
rect 18880 3485 18889 3519
rect 18889 3485 18923 3519
rect 18923 3485 18932 3519
rect 18880 3476 18932 3485
rect 19340 3519 19392 3528
rect 19340 3485 19349 3519
rect 19349 3485 19383 3519
rect 19383 3485 19392 3519
rect 19340 3476 19392 3485
rect 20076 3476 20128 3528
rect 21088 3519 21140 3528
rect 21088 3485 21097 3519
rect 21097 3485 21131 3519
rect 21131 3485 21140 3519
rect 21088 3476 21140 3485
rect 22284 3612 22336 3664
rect 21916 3544 21968 3596
rect 23020 3544 23072 3596
rect 23204 3476 23256 3528
rect 16764 3408 16816 3460
rect 17684 3408 17736 3460
rect 4620 3383 4672 3392
rect 4620 3349 4629 3383
rect 4629 3349 4663 3383
rect 4663 3349 4672 3383
rect 4620 3340 4672 3349
rect 8300 3383 8352 3392
rect 8300 3349 8309 3383
rect 8309 3349 8343 3383
rect 8343 3349 8352 3383
rect 8300 3340 8352 3349
rect 8760 3383 8812 3392
rect 8760 3349 8769 3383
rect 8769 3349 8803 3383
rect 8803 3349 8812 3383
rect 8760 3340 8812 3349
rect 8852 3340 8904 3392
rect 9956 3340 10008 3392
rect 10048 3340 10100 3392
rect 10324 3340 10376 3392
rect 11980 3340 12032 3392
rect 13820 3340 13872 3392
rect 14188 3340 14240 3392
rect 15200 3340 15252 3392
rect 15844 3340 15896 3392
rect 17408 3340 17460 3392
rect 18052 3408 18104 3460
rect 20260 3408 20312 3460
rect 20168 3340 20220 3392
rect 20536 3340 20588 3392
rect 21180 3340 21232 3392
rect 21732 3340 21784 3392
rect 22284 3383 22336 3392
rect 22284 3349 22293 3383
rect 22293 3349 22327 3383
rect 22327 3349 22336 3383
rect 22284 3340 22336 3349
rect 22744 3383 22796 3392
rect 22744 3349 22753 3383
rect 22753 3349 22787 3383
rect 22787 3349 22796 3383
rect 22744 3340 22796 3349
rect 1366 3238 1418 3290
rect 1430 3238 1482 3290
rect 1494 3238 1546 3290
rect 1558 3238 1610 3290
rect 1622 3238 1674 3290
rect 1686 3238 1738 3290
rect 7366 3238 7418 3290
rect 7430 3238 7482 3290
rect 7494 3238 7546 3290
rect 7558 3238 7610 3290
rect 7622 3238 7674 3290
rect 7686 3238 7738 3290
rect 13366 3238 13418 3290
rect 13430 3238 13482 3290
rect 13494 3238 13546 3290
rect 13558 3238 13610 3290
rect 13622 3238 13674 3290
rect 13686 3238 13738 3290
rect 19366 3238 19418 3290
rect 19430 3238 19482 3290
rect 19494 3238 19546 3290
rect 19558 3238 19610 3290
rect 19622 3238 19674 3290
rect 19686 3238 19738 3290
rect 1032 3000 1084 3052
rect 2044 3136 2096 3188
rect 6736 3136 6788 3188
rect 7196 3136 7248 3188
rect 8668 3136 8720 3188
rect 9404 3136 9456 3188
rect 10692 3136 10744 3188
rect 10784 3179 10836 3188
rect 10784 3145 10793 3179
rect 10793 3145 10827 3179
rect 10827 3145 10836 3179
rect 10784 3136 10836 3145
rect 11520 3136 11572 3188
rect 11888 3136 11940 3188
rect 1952 3068 2004 3120
rect 3884 3068 3936 3120
rect 4620 3043 4672 3052
rect 4620 3009 4629 3043
rect 4629 3009 4663 3043
rect 4663 3009 4672 3043
rect 4620 3000 4672 3009
rect 4988 3043 5040 3052
rect 4988 3009 4997 3043
rect 4997 3009 5031 3043
rect 5031 3009 5040 3043
rect 4988 3000 5040 3009
rect 3148 2932 3200 2984
rect 4252 2932 4304 2984
rect 5356 2975 5408 2984
rect 5356 2941 5365 2975
rect 5365 2941 5399 2975
rect 5399 2941 5408 2975
rect 5356 2932 5408 2941
rect 6000 3068 6052 3120
rect 6828 3000 6880 3052
rect 8300 3000 8352 3052
rect 9220 3068 9272 3120
rect 5724 2932 5776 2984
rect 7288 2932 7340 2984
rect 7472 2975 7524 2984
rect 7472 2941 7481 2975
rect 7481 2941 7515 2975
rect 7515 2941 7524 2975
rect 7472 2932 7524 2941
rect 9312 3043 9364 3052
rect 9312 3009 9321 3043
rect 9321 3009 9355 3043
rect 9355 3009 9364 3043
rect 9312 3000 9364 3009
rect 9588 3068 9640 3120
rect 12532 3068 12584 3120
rect 13452 3068 13504 3120
rect 15200 3068 15252 3120
rect 17132 3068 17184 3120
rect 17316 3111 17368 3120
rect 17316 3077 17325 3111
rect 17325 3077 17359 3111
rect 17359 3077 17368 3111
rect 17316 3068 17368 3077
rect 17408 3111 17460 3120
rect 17408 3077 17417 3111
rect 17417 3077 17451 3111
rect 17451 3077 17460 3111
rect 17408 3068 17460 3077
rect 17776 3111 17828 3120
rect 17776 3077 17785 3111
rect 17785 3077 17819 3111
rect 17819 3077 17828 3111
rect 17776 3068 17828 3077
rect 19892 3136 19944 3188
rect 20444 3136 20496 3188
rect 20536 3179 20588 3188
rect 20536 3145 20545 3179
rect 20545 3145 20579 3179
rect 20579 3145 20588 3179
rect 20536 3136 20588 3145
rect 9588 2975 9640 2984
rect 9588 2941 9597 2975
rect 9597 2941 9631 2975
rect 9631 2941 9640 2975
rect 9588 2932 9640 2941
rect 10232 3000 10284 3052
rect 10140 2975 10192 2984
rect 10140 2941 10149 2975
rect 10149 2941 10183 2975
rect 10183 2941 10192 2975
rect 10140 2932 10192 2941
rect 11796 3000 11848 3052
rect 12256 3000 12308 3052
rect 10784 2932 10836 2984
rect 11060 2932 11112 2984
rect 11244 2932 11296 2984
rect 11336 2975 11388 2984
rect 11336 2941 11345 2975
rect 11345 2941 11379 2975
rect 11379 2941 11388 2975
rect 11336 2932 11388 2941
rect 11520 2975 11572 2984
rect 11520 2941 11529 2975
rect 11529 2941 11563 2975
rect 11563 2941 11572 2975
rect 11520 2932 11572 2941
rect 11612 2975 11664 2984
rect 11612 2941 11621 2975
rect 11621 2941 11655 2975
rect 11655 2941 11664 2975
rect 11612 2932 11664 2941
rect 12900 2932 12952 2984
rect 13728 2975 13780 2984
rect 13728 2941 13737 2975
rect 13737 2941 13771 2975
rect 13771 2941 13780 2975
rect 13728 2932 13780 2941
rect 14096 2975 14148 2984
rect 14096 2941 14105 2975
rect 14105 2941 14139 2975
rect 14139 2941 14148 2975
rect 14096 2932 14148 2941
rect 14464 2932 14516 2984
rect 16672 2932 16724 2984
rect 17408 2932 17460 2984
rect 12348 2864 12400 2916
rect 4252 2796 4304 2848
rect 5816 2839 5868 2848
rect 5816 2805 5825 2839
rect 5825 2805 5859 2839
rect 5859 2805 5868 2839
rect 5816 2796 5868 2805
rect 7288 2796 7340 2848
rect 8484 2839 8536 2848
rect 8484 2805 8493 2839
rect 8493 2805 8527 2839
rect 8527 2805 8536 2839
rect 8484 2796 8536 2805
rect 9128 2839 9180 2848
rect 9128 2805 9137 2839
rect 9137 2805 9171 2839
rect 9171 2805 9180 2839
rect 9128 2796 9180 2805
rect 11520 2796 11572 2848
rect 12072 2796 12124 2848
rect 12624 2839 12676 2848
rect 12624 2805 12633 2839
rect 12633 2805 12667 2839
rect 12667 2805 12676 2839
rect 12624 2796 12676 2805
rect 13544 2907 13596 2916
rect 13544 2873 13553 2907
rect 13553 2873 13587 2907
rect 13587 2873 13596 2907
rect 13544 2864 13596 2873
rect 17592 2932 17644 2984
rect 18604 2932 18656 2984
rect 19800 3000 19852 3052
rect 19984 2975 20036 2984
rect 19984 2941 19993 2975
rect 19993 2941 20027 2975
rect 20027 2941 20036 2975
rect 19984 2932 20036 2941
rect 20628 3043 20680 3052
rect 20628 3009 20637 3043
rect 20637 3009 20671 3043
rect 20671 3009 20680 3043
rect 20628 3000 20680 3009
rect 20996 3000 21048 3052
rect 21916 3068 21968 3120
rect 23572 3068 23624 3120
rect 20904 2975 20956 2984
rect 20904 2941 20913 2975
rect 20913 2941 20947 2975
rect 20947 2941 20956 2975
rect 20904 2932 20956 2941
rect 21272 2975 21324 2984
rect 21272 2941 21281 2975
rect 21281 2941 21315 2975
rect 21315 2941 21324 2975
rect 21272 2932 21324 2941
rect 22008 3000 22060 3052
rect 21824 2975 21876 2984
rect 21824 2941 21833 2975
rect 21833 2941 21867 2975
rect 21867 2941 21876 2975
rect 21824 2932 21876 2941
rect 22836 3000 22888 3052
rect 22744 2975 22796 2984
rect 22744 2941 22753 2975
rect 22753 2941 22787 2975
rect 22787 2941 22796 2975
rect 22744 2932 22796 2941
rect 15016 2839 15068 2848
rect 15016 2805 15025 2839
rect 15025 2805 15059 2839
rect 15059 2805 15068 2839
rect 15016 2796 15068 2805
rect 16212 2796 16264 2848
rect 16764 2796 16816 2848
rect 17132 2796 17184 2848
rect 20812 2864 20864 2916
rect 19892 2796 19944 2848
rect 19984 2796 20036 2848
rect 20904 2796 20956 2848
rect 21456 2796 21508 2848
rect 21824 2796 21876 2848
rect 23296 2864 23348 2916
rect 22836 2796 22888 2848
rect 4366 2694 4418 2746
rect 4430 2694 4482 2746
rect 4494 2694 4546 2746
rect 4558 2694 4610 2746
rect 4622 2694 4674 2746
rect 4686 2694 4738 2746
rect 10366 2694 10418 2746
rect 10430 2694 10482 2746
rect 10494 2694 10546 2746
rect 10558 2694 10610 2746
rect 10622 2694 10674 2746
rect 10686 2694 10738 2746
rect 16366 2694 16418 2746
rect 16430 2694 16482 2746
rect 16494 2694 16546 2746
rect 16558 2694 16610 2746
rect 16622 2694 16674 2746
rect 16686 2694 16738 2746
rect 22366 2694 22418 2746
rect 22430 2694 22482 2746
rect 22494 2694 22546 2746
rect 22558 2694 22610 2746
rect 22622 2694 22674 2746
rect 22686 2694 22738 2746
rect 3332 2524 3384 2576
rect 3148 2363 3200 2372
rect 3148 2329 3157 2363
rect 3157 2329 3191 2363
rect 3191 2329 3200 2363
rect 3148 2320 3200 2329
rect 3424 2499 3476 2508
rect 3424 2465 3433 2499
rect 3433 2465 3467 2499
rect 3467 2465 3476 2499
rect 3424 2456 3476 2465
rect 5080 2592 5132 2644
rect 5540 2635 5592 2644
rect 5540 2601 5549 2635
rect 5549 2601 5583 2635
rect 5583 2601 5592 2635
rect 5540 2592 5592 2601
rect 5724 2592 5776 2644
rect 6552 2635 6604 2644
rect 6552 2601 6561 2635
rect 6561 2601 6595 2635
rect 6595 2601 6604 2635
rect 6552 2592 6604 2601
rect 7472 2592 7524 2644
rect 10784 2592 10836 2644
rect 11336 2592 11388 2644
rect 11520 2635 11572 2644
rect 11520 2601 11529 2635
rect 11529 2601 11563 2635
rect 11563 2601 11572 2635
rect 11520 2592 11572 2601
rect 11704 2592 11756 2644
rect 11796 2592 11848 2644
rect 11888 2592 11940 2644
rect 3884 2388 3936 2440
rect 6000 2456 6052 2508
rect 6828 2567 6880 2576
rect 6828 2533 6837 2567
rect 6837 2533 6871 2567
rect 6871 2533 6880 2567
rect 6828 2524 6880 2533
rect 6736 2456 6788 2508
rect 7748 2456 7800 2508
rect 9128 2524 9180 2576
rect 9588 2524 9640 2576
rect 9680 2524 9732 2576
rect 5816 2388 5868 2440
rect 7012 2431 7064 2440
rect 7012 2397 7021 2431
rect 7021 2397 7055 2431
rect 7055 2397 7064 2431
rect 7012 2388 7064 2397
rect 7104 2431 7156 2440
rect 7104 2397 7113 2431
rect 7113 2397 7147 2431
rect 7147 2397 7156 2431
rect 7104 2388 7156 2397
rect 8484 2499 8536 2508
rect 8484 2465 8493 2499
rect 8493 2465 8527 2499
rect 8527 2465 8536 2499
rect 8484 2456 8536 2465
rect 8760 2499 8812 2508
rect 8760 2465 8769 2499
rect 8769 2465 8803 2499
rect 8803 2465 8812 2499
rect 8760 2456 8812 2465
rect 8944 2388 8996 2440
rect 9496 2499 9548 2508
rect 9496 2465 9505 2499
rect 9505 2465 9539 2499
rect 9539 2465 9548 2499
rect 9496 2456 9548 2465
rect 10048 2499 10100 2508
rect 10048 2465 10057 2499
rect 10057 2465 10091 2499
rect 10091 2465 10100 2499
rect 10048 2456 10100 2465
rect 6184 2320 6236 2372
rect 3976 2252 4028 2304
rect 8300 2320 8352 2372
rect 9772 2320 9824 2372
rect 7840 2295 7892 2304
rect 7840 2261 7849 2295
rect 7849 2261 7883 2295
rect 7883 2261 7892 2295
rect 7840 2252 7892 2261
rect 8116 2252 8168 2304
rect 8760 2252 8812 2304
rect 9128 2252 9180 2304
rect 9404 2252 9456 2304
rect 10416 2499 10468 2508
rect 10416 2465 10425 2499
rect 10425 2465 10459 2499
rect 10459 2465 10468 2499
rect 10416 2456 10468 2465
rect 10968 2499 11020 2508
rect 10968 2465 10977 2499
rect 10977 2465 11011 2499
rect 11011 2465 11020 2499
rect 10968 2456 11020 2465
rect 11244 2388 11296 2440
rect 11704 2499 11756 2508
rect 11704 2465 11713 2499
rect 11713 2465 11747 2499
rect 11747 2465 11756 2499
rect 11704 2456 11756 2465
rect 12348 2592 12400 2644
rect 13544 2592 13596 2644
rect 12440 2567 12492 2576
rect 12440 2533 12449 2567
rect 12449 2533 12483 2567
rect 12483 2533 12492 2567
rect 12440 2524 12492 2533
rect 16580 2635 16632 2644
rect 16580 2601 16589 2635
rect 16589 2601 16623 2635
rect 16623 2601 16632 2635
rect 16580 2592 16632 2601
rect 16212 2524 16264 2576
rect 12164 2456 12216 2508
rect 12256 2456 12308 2508
rect 12532 2456 12584 2508
rect 12900 2499 12952 2508
rect 12900 2465 12909 2499
rect 12909 2465 12943 2499
rect 12943 2465 12952 2499
rect 12900 2456 12952 2465
rect 13084 2456 13136 2508
rect 11428 2320 11480 2372
rect 11520 2252 11572 2304
rect 12624 2295 12676 2304
rect 12624 2261 12633 2295
rect 12633 2261 12667 2295
rect 12667 2261 12676 2295
rect 12624 2252 12676 2261
rect 12900 2320 12952 2372
rect 13544 2499 13596 2508
rect 13544 2465 13553 2499
rect 13553 2465 13587 2499
rect 13587 2465 13596 2499
rect 13544 2456 13596 2465
rect 13728 2499 13780 2508
rect 13728 2465 13737 2499
rect 13737 2465 13771 2499
rect 13771 2465 13780 2499
rect 13728 2456 13780 2465
rect 13820 2499 13872 2508
rect 13820 2465 13829 2499
rect 13829 2465 13863 2499
rect 13863 2465 13872 2499
rect 13820 2456 13872 2465
rect 14556 2456 14608 2508
rect 15016 2499 15068 2508
rect 15016 2465 15025 2499
rect 15025 2465 15059 2499
rect 15059 2465 15068 2499
rect 15016 2456 15068 2465
rect 15200 2456 15252 2508
rect 15384 2499 15436 2508
rect 15384 2465 15393 2499
rect 15393 2465 15427 2499
rect 15427 2465 15436 2499
rect 15384 2456 15436 2465
rect 16304 2499 16356 2508
rect 16304 2465 16313 2499
rect 16313 2465 16347 2499
rect 16347 2465 16356 2499
rect 16304 2456 16356 2465
rect 16856 2524 16908 2576
rect 17776 2524 17828 2576
rect 16212 2388 16264 2440
rect 17040 2499 17092 2508
rect 17040 2465 17049 2499
rect 17049 2465 17083 2499
rect 17083 2465 17092 2499
rect 17040 2456 17092 2465
rect 16856 2388 16908 2440
rect 17684 2456 17736 2508
rect 18788 2499 18840 2508
rect 18788 2465 18797 2499
rect 18797 2465 18831 2499
rect 18831 2465 18840 2499
rect 18788 2456 18840 2465
rect 19156 2499 19208 2508
rect 19156 2465 19165 2499
rect 19165 2465 19199 2499
rect 19199 2465 19208 2499
rect 19156 2456 19208 2465
rect 15384 2320 15436 2372
rect 17868 2320 17920 2372
rect 14004 2252 14056 2304
rect 14096 2295 14148 2304
rect 14096 2261 14105 2295
rect 14105 2261 14139 2295
rect 14139 2261 14148 2295
rect 14096 2252 14148 2261
rect 16212 2252 16264 2304
rect 17040 2252 17092 2304
rect 17132 2252 17184 2304
rect 17408 2252 17460 2304
rect 19800 2320 19852 2372
rect 20720 2499 20772 2508
rect 20720 2465 20729 2499
rect 20729 2465 20763 2499
rect 20763 2465 20772 2499
rect 20720 2456 20772 2465
rect 20812 2388 20864 2440
rect 21456 2524 21508 2576
rect 21640 2499 21692 2508
rect 21640 2465 21649 2499
rect 21649 2465 21683 2499
rect 21683 2465 21692 2499
rect 21640 2456 21692 2465
rect 20260 2320 20312 2372
rect 22376 2592 22428 2644
rect 23112 2592 23164 2644
rect 22192 2499 22244 2508
rect 22192 2465 22201 2499
rect 22201 2465 22235 2499
rect 22235 2465 22244 2499
rect 22192 2456 22244 2465
rect 21916 2388 21968 2440
rect 22468 2499 22520 2508
rect 22468 2465 22477 2499
rect 22477 2465 22511 2499
rect 22511 2465 22520 2499
rect 22468 2456 22520 2465
rect 22928 2456 22980 2508
rect 18604 2252 18656 2304
rect 18880 2295 18932 2304
rect 18880 2261 18889 2295
rect 18889 2261 18923 2295
rect 18923 2261 18932 2295
rect 18880 2252 18932 2261
rect 18972 2252 19024 2304
rect 20444 2295 20496 2304
rect 20444 2261 20453 2295
rect 20453 2261 20487 2295
rect 20487 2261 20496 2295
rect 20444 2252 20496 2261
rect 20812 2252 20864 2304
rect 21364 2252 21416 2304
rect 21916 2295 21968 2304
rect 21916 2261 21925 2295
rect 21925 2261 21959 2295
rect 21959 2261 21968 2295
rect 21916 2252 21968 2261
rect 22100 2252 22152 2304
rect 22376 2252 22428 2304
rect 22560 2295 22612 2304
rect 22560 2261 22569 2295
rect 22569 2261 22603 2295
rect 22603 2261 22612 2295
rect 22560 2252 22612 2261
rect 1366 2150 1418 2202
rect 1430 2150 1482 2202
rect 1494 2150 1546 2202
rect 1558 2150 1610 2202
rect 1622 2150 1674 2202
rect 1686 2150 1738 2202
rect 7366 2150 7418 2202
rect 7430 2150 7482 2202
rect 7494 2150 7546 2202
rect 7558 2150 7610 2202
rect 7622 2150 7674 2202
rect 7686 2150 7738 2202
rect 13366 2150 13418 2202
rect 13430 2150 13482 2202
rect 13494 2150 13546 2202
rect 13558 2150 13610 2202
rect 13622 2150 13674 2202
rect 13686 2150 13738 2202
rect 19366 2150 19418 2202
rect 19430 2150 19482 2202
rect 19494 2150 19546 2202
rect 19558 2150 19610 2202
rect 19622 2150 19674 2202
rect 19686 2150 19738 2202
rect 3332 2048 3384 2100
rect 1860 1980 1912 2032
rect 3884 2023 3936 2032
rect 3884 1989 3893 2023
rect 3893 1989 3927 2023
rect 3927 1989 3936 2023
rect 3884 1980 3936 1989
rect 5816 2048 5868 2100
rect 7288 2048 7340 2100
rect 8760 2091 8812 2100
rect 8760 2057 8769 2091
rect 8769 2057 8803 2091
rect 8803 2057 8812 2091
rect 8760 2048 8812 2057
rect 8944 2048 8996 2100
rect 6644 1980 6696 2032
rect 2504 1912 2556 1964
rect 1952 1844 2004 1896
rect 3056 1887 3108 1896
rect 3056 1853 3065 1887
rect 3065 1853 3099 1887
rect 3099 1853 3108 1887
rect 3056 1844 3108 1853
rect 3424 1844 3476 1896
rect 2688 1751 2740 1760
rect 2688 1717 2697 1751
rect 2697 1717 2731 1751
rect 2731 1717 2740 1751
rect 2688 1708 2740 1717
rect 2780 1708 2832 1760
rect 3332 1776 3384 1828
rect 6184 1912 6236 1964
rect 6736 1912 6788 1964
rect 4988 1844 5040 1896
rect 5264 1887 5316 1896
rect 5264 1853 5273 1887
rect 5273 1853 5307 1887
rect 5307 1853 5316 1887
rect 5264 1844 5316 1853
rect 5724 1887 5776 1896
rect 5724 1853 5733 1887
rect 5733 1853 5767 1887
rect 5767 1853 5776 1887
rect 5724 1844 5776 1853
rect 6000 1844 6052 1896
rect 7012 1844 7064 1896
rect 7104 1844 7156 1896
rect 10048 1980 10100 2032
rect 10416 2091 10468 2100
rect 10416 2057 10425 2091
rect 10425 2057 10459 2091
rect 10459 2057 10468 2091
rect 10416 2048 10468 2057
rect 11612 2048 11664 2100
rect 11888 2091 11940 2100
rect 11888 2057 11897 2091
rect 11897 2057 11931 2091
rect 11931 2057 11940 2091
rect 11888 2048 11940 2057
rect 13268 2048 13320 2100
rect 14096 2048 14148 2100
rect 16580 2048 16632 2100
rect 17040 2048 17092 2100
rect 20076 2091 20128 2100
rect 20076 2057 20085 2091
rect 20085 2057 20119 2091
rect 20119 2057 20128 2091
rect 20076 2048 20128 2057
rect 22192 2048 22244 2100
rect 22376 2091 22428 2100
rect 22376 2057 22385 2091
rect 22385 2057 22419 2091
rect 22419 2057 22428 2091
rect 22376 2048 22428 2057
rect 22560 2048 22612 2100
rect 5448 1776 5500 1828
rect 3976 1708 4028 1760
rect 4160 1708 4212 1760
rect 4896 1708 4948 1760
rect 5908 1751 5960 1760
rect 5908 1717 5917 1751
rect 5917 1717 5951 1751
rect 5951 1717 5960 1751
rect 5908 1708 5960 1717
rect 7932 1708 7984 1760
rect 8484 1844 8536 1896
rect 14004 1980 14056 2032
rect 12440 1912 12492 1964
rect 14280 1912 14332 1964
rect 14372 1912 14424 1964
rect 9128 1887 9180 1896
rect 9128 1853 9137 1887
rect 9137 1853 9171 1887
rect 9171 1853 9180 1887
rect 9128 1844 9180 1853
rect 8668 1776 8720 1828
rect 9036 1776 9088 1828
rect 9312 1887 9364 1896
rect 9312 1853 9321 1887
rect 9321 1853 9355 1887
rect 9355 1853 9364 1887
rect 9312 1844 9364 1853
rect 9864 1887 9916 1896
rect 9864 1853 9873 1887
rect 9873 1853 9907 1887
rect 9907 1853 9916 1887
rect 9864 1844 9916 1853
rect 9956 1887 10008 1896
rect 9956 1853 9965 1887
rect 9965 1853 9999 1887
rect 9999 1853 10008 1887
rect 9956 1844 10008 1853
rect 10232 1887 10284 1896
rect 10232 1853 10241 1887
rect 10241 1853 10275 1887
rect 10275 1853 10284 1887
rect 10232 1844 10284 1853
rect 10324 1844 10376 1896
rect 10876 1887 10928 1896
rect 10876 1853 10904 1887
rect 10904 1853 10928 1887
rect 10876 1844 10928 1853
rect 11244 1887 11296 1896
rect 11244 1853 11253 1887
rect 11253 1853 11287 1887
rect 11287 1853 11296 1887
rect 11244 1844 11296 1853
rect 11428 1844 11480 1896
rect 11520 1887 11572 1896
rect 11520 1853 11529 1887
rect 11529 1853 11563 1887
rect 11563 1853 11572 1887
rect 11520 1844 11572 1853
rect 11612 1887 11664 1896
rect 11612 1853 11621 1887
rect 11621 1853 11655 1887
rect 11655 1853 11664 1887
rect 11612 1844 11664 1853
rect 11888 1844 11940 1896
rect 12348 1844 12400 1896
rect 12716 1844 12768 1896
rect 12900 1887 12952 1896
rect 12900 1853 12909 1887
rect 12909 1853 12943 1887
rect 12943 1853 12952 1887
rect 12900 1844 12952 1853
rect 14464 1844 14516 1896
rect 15568 1887 15620 1896
rect 15568 1853 15577 1887
rect 15577 1853 15611 1887
rect 15611 1853 15620 1887
rect 15568 1844 15620 1853
rect 15660 1887 15712 1896
rect 15660 1853 15669 1887
rect 15669 1853 15703 1887
rect 15703 1853 15712 1887
rect 15660 1844 15712 1853
rect 16120 1912 16172 1964
rect 18052 1955 18104 1964
rect 18052 1921 18061 1955
rect 18061 1921 18095 1955
rect 18095 1921 18104 1955
rect 18052 1912 18104 1921
rect 19984 1980 20036 2032
rect 17408 1844 17460 1896
rect 17776 1887 17828 1896
rect 17776 1853 17785 1887
rect 17785 1853 17819 1887
rect 17819 1853 17828 1887
rect 17776 1844 17828 1853
rect 18696 1887 18748 1896
rect 18696 1853 18705 1887
rect 18705 1853 18739 1887
rect 18739 1853 18748 1887
rect 18696 1844 18748 1853
rect 20260 1955 20312 1964
rect 20260 1921 20269 1955
rect 20269 1921 20303 1955
rect 20303 1921 20312 1955
rect 20260 1912 20312 1921
rect 13268 1776 13320 1828
rect 13728 1776 13780 1828
rect 15936 1776 15988 1828
rect 8852 1708 8904 1760
rect 9220 1708 9272 1760
rect 9588 1708 9640 1760
rect 10784 1751 10836 1760
rect 10784 1717 10793 1751
rect 10793 1717 10827 1751
rect 10827 1717 10836 1751
rect 10784 1708 10836 1717
rect 11244 1708 11296 1760
rect 11428 1751 11480 1760
rect 11428 1717 11437 1751
rect 11437 1717 11471 1751
rect 11471 1717 11480 1751
rect 11428 1708 11480 1717
rect 12624 1708 12676 1760
rect 13084 1751 13136 1760
rect 13084 1717 13093 1751
rect 13093 1717 13127 1751
rect 13127 1717 13136 1751
rect 13084 1708 13136 1717
rect 13176 1708 13228 1760
rect 13636 1708 13688 1760
rect 14648 1708 14700 1760
rect 15752 1708 15804 1760
rect 16856 1708 16908 1760
rect 18328 1776 18380 1828
rect 18972 1776 19024 1828
rect 20812 1844 20864 1896
rect 22008 1980 22060 2032
rect 22100 1980 22152 2032
rect 22376 1912 22428 1964
rect 21364 1887 21416 1896
rect 21364 1853 21373 1887
rect 21373 1853 21407 1887
rect 21407 1853 21416 1887
rect 21364 1844 21416 1853
rect 21548 1887 21600 1896
rect 21548 1853 21557 1887
rect 21557 1853 21591 1887
rect 21591 1853 21600 1887
rect 21548 1844 21600 1853
rect 21732 1887 21784 1896
rect 21732 1853 21741 1887
rect 21741 1853 21775 1887
rect 21775 1853 21784 1887
rect 21732 1844 21784 1853
rect 21640 1819 21692 1828
rect 21640 1785 21649 1819
rect 21649 1785 21683 1819
rect 21683 1785 21692 1819
rect 21640 1776 21692 1785
rect 19248 1708 19300 1760
rect 19340 1751 19392 1760
rect 19340 1717 19349 1751
rect 19349 1717 19383 1751
rect 19383 1717 19392 1751
rect 19340 1708 19392 1717
rect 19892 1751 19944 1760
rect 19892 1717 19901 1751
rect 19901 1717 19935 1751
rect 19935 1717 19944 1751
rect 19892 1708 19944 1717
rect 19984 1708 20036 1760
rect 21824 1708 21876 1760
rect 22192 1708 22244 1760
rect 22560 1887 22612 1896
rect 22560 1853 22569 1887
rect 22569 1853 22603 1887
rect 22603 1853 22612 1887
rect 22560 1844 22612 1853
rect 22744 1844 22796 1896
rect 23204 1844 23256 1896
rect 22928 1776 22980 1828
rect 23020 1708 23072 1760
rect 4366 1606 4418 1658
rect 4430 1606 4482 1658
rect 4494 1606 4546 1658
rect 4558 1606 4610 1658
rect 4622 1606 4674 1658
rect 4686 1606 4738 1658
rect 10366 1606 10418 1658
rect 10430 1606 10482 1658
rect 10494 1606 10546 1658
rect 10558 1606 10610 1658
rect 10622 1606 10674 1658
rect 10686 1606 10738 1658
rect 16366 1606 16418 1658
rect 16430 1606 16482 1658
rect 16494 1606 16546 1658
rect 16558 1606 16610 1658
rect 16622 1606 16674 1658
rect 16686 1606 16738 1658
rect 22366 1606 22418 1658
rect 22430 1606 22482 1658
rect 22494 1606 22546 1658
rect 22558 1606 22610 1658
rect 22622 1606 22674 1658
rect 22686 1606 22738 1658
rect 756 1504 808 1556
rect 572 1436 624 1488
rect 2228 1504 2280 1556
rect 2688 1436 2740 1488
rect 1860 1411 1912 1420
rect 1860 1377 1869 1411
rect 1869 1377 1903 1411
rect 1903 1377 1912 1411
rect 1860 1368 1912 1377
rect 1952 1368 2004 1420
rect 2780 1411 2832 1420
rect 2780 1377 2789 1411
rect 2789 1377 2823 1411
rect 2823 1377 2832 1411
rect 2780 1368 2832 1377
rect 3332 1411 3384 1420
rect 3332 1377 3341 1411
rect 3341 1377 3375 1411
rect 3375 1377 3384 1411
rect 3332 1368 3384 1377
rect 4252 1368 4304 1420
rect 5448 1479 5500 1488
rect 5448 1445 5457 1479
rect 5457 1445 5491 1479
rect 5491 1445 5500 1479
rect 5448 1436 5500 1445
rect 6644 1504 6696 1556
rect 8300 1547 8352 1556
rect 8300 1513 8309 1547
rect 8309 1513 8343 1547
rect 8343 1513 8352 1547
rect 8300 1504 8352 1513
rect 9312 1504 9364 1556
rect 12532 1504 12584 1556
rect 13084 1547 13136 1556
rect 13084 1513 13093 1547
rect 13093 1513 13127 1547
rect 13127 1513 13136 1547
rect 13084 1504 13136 1513
rect 5724 1368 5776 1420
rect 6000 1411 6052 1420
rect 6000 1377 6009 1411
rect 6009 1377 6043 1411
rect 6043 1377 6052 1411
rect 6000 1368 6052 1377
rect 6736 1411 6788 1420
rect 6736 1377 6745 1411
rect 6745 1377 6779 1411
rect 6779 1377 6788 1411
rect 6736 1368 6788 1377
rect 8576 1436 8628 1488
rect 7840 1368 7892 1420
rect 7932 1411 7984 1420
rect 7932 1377 7941 1411
rect 7941 1377 7975 1411
rect 7975 1377 7984 1411
rect 7932 1368 7984 1377
rect 8116 1411 8168 1420
rect 8116 1377 8125 1411
rect 8125 1377 8159 1411
rect 8159 1377 8168 1411
rect 8116 1368 8168 1377
rect 8484 1411 8536 1420
rect 8484 1377 8493 1411
rect 8493 1377 8527 1411
rect 8527 1377 8536 1411
rect 8484 1368 8536 1377
rect 9128 1436 9180 1488
rect 8944 1411 8996 1420
rect 8944 1377 8953 1411
rect 8953 1377 8987 1411
rect 8987 1377 8996 1411
rect 8944 1368 8996 1377
rect 9404 1411 9456 1420
rect 9404 1377 9413 1411
rect 9413 1377 9447 1411
rect 9447 1377 9456 1411
rect 9404 1368 9456 1377
rect 3608 1300 3660 1352
rect 6828 1343 6880 1352
rect 6828 1309 6837 1343
rect 6837 1309 6871 1343
rect 6871 1309 6880 1343
rect 6828 1300 6880 1309
rect 7104 1343 7156 1352
rect 7104 1309 7113 1343
rect 7113 1309 7147 1343
rect 7147 1309 7156 1343
rect 7104 1300 7156 1309
rect 6368 1275 6420 1284
rect 6368 1241 6377 1275
rect 6377 1241 6411 1275
rect 6411 1241 6420 1275
rect 6368 1232 6420 1241
rect 8024 1232 8076 1284
rect 9128 1300 9180 1352
rect 9496 1300 9548 1352
rect 1768 1164 1820 1216
rect 2964 1207 3016 1216
rect 2964 1173 2973 1207
rect 2973 1173 3007 1207
rect 3007 1173 3016 1207
rect 2964 1164 3016 1173
rect 6184 1164 6236 1216
rect 8484 1164 8536 1216
rect 9772 1368 9824 1420
rect 9956 1300 10008 1352
rect 10048 1300 10100 1352
rect 11336 1411 11388 1420
rect 11336 1377 11345 1411
rect 11345 1377 11379 1411
rect 11379 1377 11388 1411
rect 11336 1368 11388 1377
rect 11704 1411 11756 1420
rect 11704 1377 11713 1411
rect 11713 1377 11747 1411
rect 11747 1377 11756 1411
rect 11704 1368 11756 1377
rect 11980 1411 12032 1420
rect 11980 1377 11989 1411
rect 11989 1377 12023 1411
rect 12023 1377 12032 1411
rect 11980 1368 12032 1377
rect 12072 1411 12124 1420
rect 12072 1377 12081 1411
rect 12081 1377 12115 1411
rect 12115 1377 12124 1411
rect 12072 1368 12124 1377
rect 12808 1368 12860 1420
rect 12992 1411 13044 1420
rect 12992 1377 13001 1411
rect 13001 1377 13035 1411
rect 13035 1377 13044 1411
rect 12992 1368 13044 1377
rect 13084 1368 13136 1420
rect 13636 1411 13688 1420
rect 13636 1377 13645 1411
rect 13645 1377 13679 1411
rect 13679 1377 13688 1411
rect 13636 1368 13688 1377
rect 13728 1368 13780 1420
rect 13360 1343 13412 1352
rect 9680 1232 9732 1284
rect 9864 1232 9916 1284
rect 10784 1232 10836 1284
rect 10876 1232 10928 1284
rect 10140 1164 10192 1216
rect 11520 1164 11572 1216
rect 13360 1309 13369 1343
rect 13369 1309 13403 1343
rect 13403 1309 13412 1343
rect 13360 1300 13412 1309
rect 15660 1547 15712 1556
rect 15660 1513 15675 1547
rect 15675 1513 15709 1547
rect 15709 1513 15712 1547
rect 15660 1504 15712 1513
rect 16212 1504 16264 1556
rect 14372 1436 14424 1488
rect 14556 1368 14608 1420
rect 14924 1436 14976 1488
rect 15384 1479 15436 1488
rect 15384 1445 15393 1479
rect 15393 1445 15427 1479
rect 15427 1445 15436 1479
rect 15384 1436 15436 1445
rect 18512 1504 18564 1556
rect 18696 1504 18748 1556
rect 19892 1504 19944 1556
rect 22284 1504 22336 1556
rect 22376 1504 22428 1556
rect 23296 1504 23348 1556
rect 15108 1411 15160 1420
rect 15108 1377 15117 1411
rect 15117 1377 15151 1411
rect 15151 1377 15160 1411
rect 15108 1368 15160 1377
rect 15200 1411 15252 1420
rect 15200 1377 15209 1411
rect 15209 1377 15243 1411
rect 15243 1377 15252 1411
rect 15200 1368 15252 1377
rect 15752 1411 15804 1420
rect 15752 1377 15761 1411
rect 15761 1377 15795 1411
rect 15795 1377 15804 1411
rect 15752 1368 15804 1377
rect 15844 1411 15896 1420
rect 15844 1377 15853 1411
rect 15853 1377 15887 1411
rect 15887 1377 15896 1411
rect 15844 1368 15896 1377
rect 16120 1368 16172 1420
rect 16580 1411 16632 1420
rect 16580 1377 16589 1411
rect 16589 1377 16623 1411
rect 16623 1377 16632 1411
rect 16580 1368 16632 1377
rect 15568 1300 15620 1352
rect 17132 1411 17184 1420
rect 17132 1377 17141 1411
rect 17141 1377 17175 1411
rect 17175 1377 17184 1411
rect 17132 1368 17184 1377
rect 18604 1411 18656 1420
rect 18604 1377 18613 1411
rect 18613 1377 18647 1411
rect 18647 1377 18656 1411
rect 18604 1368 18656 1377
rect 18972 1411 19024 1420
rect 18972 1377 18981 1411
rect 18981 1377 19015 1411
rect 19015 1377 19024 1411
rect 18972 1368 19024 1377
rect 19064 1411 19116 1420
rect 19064 1377 19073 1411
rect 19073 1377 19107 1411
rect 19107 1377 19116 1411
rect 19064 1368 19116 1377
rect 19708 1411 19760 1420
rect 19708 1377 19717 1411
rect 19717 1377 19751 1411
rect 19751 1377 19760 1411
rect 19708 1368 19760 1377
rect 19800 1368 19852 1420
rect 20352 1411 20404 1420
rect 20352 1377 20361 1411
rect 20361 1377 20395 1411
rect 20395 1377 20404 1411
rect 20352 1368 20404 1377
rect 20720 1436 20772 1488
rect 21732 1436 21784 1488
rect 16856 1300 16908 1352
rect 12348 1232 12400 1284
rect 13084 1164 13136 1216
rect 14280 1275 14332 1284
rect 14280 1241 14289 1275
rect 14289 1241 14323 1275
rect 14323 1241 14332 1275
rect 14280 1232 14332 1241
rect 14464 1232 14516 1284
rect 17592 1343 17644 1352
rect 17592 1309 17601 1343
rect 17601 1309 17635 1343
rect 17635 1309 17644 1343
rect 17592 1300 17644 1309
rect 18604 1275 18656 1284
rect 18604 1241 18613 1275
rect 18613 1241 18647 1275
rect 18647 1241 18656 1275
rect 18604 1232 18656 1241
rect 18696 1232 18748 1284
rect 20076 1300 20128 1352
rect 20444 1300 20496 1352
rect 20628 1343 20680 1352
rect 20628 1309 20637 1343
rect 20637 1309 20671 1343
rect 20671 1309 20680 1343
rect 20628 1300 20680 1309
rect 20812 1368 20864 1420
rect 21548 1411 21600 1420
rect 21548 1377 21557 1411
rect 21557 1377 21591 1411
rect 21591 1377 21600 1411
rect 21548 1368 21600 1377
rect 22376 1368 22428 1420
rect 21916 1300 21968 1352
rect 23020 1436 23072 1488
rect 22928 1368 22980 1420
rect 23388 1300 23440 1352
rect 19892 1275 19944 1284
rect 19892 1241 19901 1275
rect 19901 1241 19935 1275
rect 19935 1241 19944 1275
rect 19892 1232 19944 1241
rect 13820 1207 13872 1216
rect 13820 1173 13829 1207
rect 13829 1173 13863 1207
rect 13863 1173 13872 1207
rect 13820 1164 13872 1173
rect 15016 1207 15068 1216
rect 15016 1173 15025 1207
rect 15025 1173 15059 1207
rect 15059 1173 15068 1207
rect 15016 1164 15068 1173
rect 15108 1164 15160 1216
rect 17684 1207 17736 1216
rect 17684 1173 17693 1207
rect 17693 1173 17727 1207
rect 17727 1173 17736 1207
rect 17684 1164 17736 1173
rect 17776 1207 17828 1216
rect 17776 1173 17785 1207
rect 17785 1173 17819 1207
rect 17819 1173 17828 1207
rect 17776 1164 17828 1173
rect 18328 1164 18380 1216
rect 19064 1164 19116 1216
rect 20076 1207 20128 1216
rect 20076 1173 20085 1207
rect 20085 1173 20119 1207
rect 20119 1173 20128 1207
rect 20076 1164 20128 1173
rect 20352 1164 20404 1216
rect 20444 1207 20496 1216
rect 20444 1173 20453 1207
rect 20453 1173 20487 1207
rect 20487 1173 20496 1207
rect 20444 1164 20496 1173
rect 20536 1207 20588 1216
rect 20536 1173 20545 1207
rect 20545 1173 20579 1207
rect 20579 1173 20588 1207
rect 20536 1164 20588 1173
rect 20812 1207 20864 1216
rect 20812 1173 20821 1207
rect 20821 1173 20855 1207
rect 20855 1173 20864 1207
rect 20812 1164 20864 1173
rect 20904 1164 20956 1216
rect 1366 1062 1418 1114
rect 1430 1062 1482 1114
rect 1494 1062 1546 1114
rect 1558 1062 1610 1114
rect 1622 1062 1674 1114
rect 1686 1062 1738 1114
rect 7366 1062 7418 1114
rect 7430 1062 7482 1114
rect 7494 1062 7546 1114
rect 7558 1062 7610 1114
rect 7622 1062 7674 1114
rect 7686 1062 7738 1114
rect 13366 1062 13418 1114
rect 13430 1062 13482 1114
rect 13494 1062 13546 1114
rect 13558 1062 13610 1114
rect 13622 1062 13674 1114
rect 13686 1062 13738 1114
rect 19366 1062 19418 1114
rect 19430 1062 19482 1114
rect 19494 1062 19546 1114
rect 19558 1062 19610 1114
rect 19622 1062 19674 1114
rect 19686 1062 19738 1114
rect 3332 960 3384 1012
rect 6000 960 6052 1012
rect 6092 960 6144 1012
rect 6828 1003 6880 1012
rect 6828 969 6837 1003
rect 6837 969 6871 1003
rect 6871 969 6880 1003
rect 6828 960 6880 969
rect 7840 960 7892 1012
rect 8484 960 8536 1012
rect 9956 960 10008 1012
rect 11336 1003 11388 1012
rect 11336 969 11345 1003
rect 11345 969 11379 1003
rect 11379 969 11388 1003
rect 11336 960 11388 969
rect 11520 960 11572 1012
rect 14188 960 14240 1012
rect 15016 960 15068 1012
rect 16580 960 16632 1012
rect 2596 892 2648 944
rect 3056 892 3108 944
rect 4068 892 4120 944
rect 5172 892 5224 944
rect 1216 799 1268 808
rect 1216 765 1225 799
rect 1225 765 1259 799
rect 1259 765 1268 799
rect 1216 756 1268 765
rect 1768 756 1820 808
rect 1952 799 2004 808
rect 1952 765 1961 799
rect 1961 765 1995 799
rect 1995 765 2004 799
rect 1952 756 2004 765
rect 3424 799 3476 808
rect 3424 765 3433 799
rect 3433 765 3467 799
rect 3467 765 3476 799
rect 3424 756 3476 765
rect 4160 799 4212 808
rect 4160 765 4169 799
rect 4169 765 4203 799
rect 4203 765 4212 799
rect 4160 756 4212 765
rect 4528 799 4580 808
rect 4528 765 4537 799
rect 4537 765 4571 799
rect 4571 765 4580 799
rect 4528 756 4580 765
rect 4896 799 4948 808
rect 4896 765 4905 799
rect 4905 765 4939 799
rect 4939 765 4948 799
rect 4896 756 4948 765
rect 7104 892 7156 944
rect 7932 824 7984 876
rect 5908 799 5960 808
rect 5908 765 5917 799
rect 5917 765 5951 799
rect 5951 765 5960 799
rect 5908 756 5960 765
rect 6184 799 6236 808
rect 6184 765 6193 799
rect 6193 765 6227 799
rect 6227 765 6236 799
rect 6184 756 6236 765
rect 7104 799 7156 808
rect 7104 765 7113 799
rect 7113 765 7147 799
rect 7147 765 7156 799
rect 7104 756 7156 765
rect 7196 799 7248 808
rect 7196 765 7205 799
rect 7205 765 7239 799
rect 7239 765 7248 799
rect 7196 756 7248 765
rect 7840 756 7892 808
rect 8116 756 8168 808
rect 9588 892 9640 944
rect 10968 892 11020 944
rect 11428 892 11480 944
rect 14924 892 14976 944
rect 9312 824 9364 876
rect 10692 824 10744 876
rect 4988 688 5040 740
rect 1124 620 1176 672
rect 1492 620 1544 672
rect 1860 620 1912 672
rect 3700 620 3752 672
rect 4252 620 4304 672
rect 4804 620 4856 672
rect 5540 688 5592 740
rect 6736 688 6788 740
rect 8852 756 8904 808
rect 5816 620 5868 672
rect 7748 663 7800 672
rect 7748 629 7757 663
rect 7757 629 7791 663
rect 7791 629 7800 663
rect 7748 620 7800 629
rect 9128 688 9180 740
rect 9772 799 9824 808
rect 9772 765 9781 799
rect 9781 765 9815 799
rect 9815 765 9824 799
rect 9772 756 9824 765
rect 10140 799 10192 808
rect 10140 765 10149 799
rect 10149 765 10183 799
rect 10183 765 10192 799
rect 10140 756 10192 765
rect 11060 799 11112 808
rect 11060 765 11069 799
rect 11069 765 11103 799
rect 11103 765 11112 799
rect 11060 756 11112 765
rect 9864 620 9916 672
rect 10232 620 10284 672
rect 11152 663 11204 672
rect 11152 629 11161 663
rect 11161 629 11195 663
rect 11195 629 11204 663
rect 11152 620 11204 629
rect 11336 731 11388 740
rect 11336 697 11345 731
rect 11345 697 11379 731
rect 11379 697 11388 731
rect 11336 688 11388 697
rect 11704 756 11756 808
rect 13176 824 13228 876
rect 14372 824 14424 876
rect 20260 960 20312 1012
rect 21824 1003 21876 1012
rect 21824 969 21833 1003
rect 21833 969 21867 1003
rect 21867 969 21876 1003
rect 21824 960 21876 969
rect 11888 799 11940 808
rect 11888 765 11897 799
rect 11897 765 11931 799
rect 11931 765 11940 799
rect 11888 756 11940 765
rect 11520 731 11572 740
rect 11520 697 11529 731
rect 11529 697 11563 731
rect 11563 697 11572 731
rect 11520 688 11572 697
rect 12624 799 12676 808
rect 12624 765 12633 799
rect 12633 765 12667 799
rect 12667 765 12676 799
rect 12624 756 12676 765
rect 13268 799 13320 808
rect 13268 765 13277 799
rect 13277 765 13311 799
rect 13311 765 13320 799
rect 13268 756 13320 765
rect 13820 799 13872 808
rect 13820 765 13829 799
rect 13829 765 13863 799
rect 13863 765 13872 799
rect 13820 756 13872 765
rect 14464 756 14516 808
rect 14556 799 14608 808
rect 14556 765 14565 799
rect 14565 765 14599 799
rect 14599 765 14608 799
rect 14556 756 14608 765
rect 14648 799 14700 808
rect 14648 765 14657 799
rect 14657 765 14691 799
rect 14691 765 14700 799
rect 14648 756 14700 765
rect 16212 756 16264 808
rect 16764 756 16816 808
rect 17684 824 17736 876
rect 19156 892 19208 944
rect 19800 892 19852 944
rect 20444 892 20496 944
rect 20996 892 21048 944
rect 17868 799 17920 808
rect 17868 765 17877 799
rect 17877 765 17911 799
rect 17911 765 17920 799
rect 17868 756 17920 765
rect 19984 824 20036 876
rect 12716 688 12768 740
rect 14372 688 14424 740
rect 19064 799 19116 808
rect 19064 765 19073 799
rect 19073 765 19107 799
rect 19107 765 19116 799
rect 19064 756 19116 765
rect 19248 756 19300 808
rect 19800 799 19852 808
rect 19800 765 19809 799
rect 19809 765 19843 799
rect 19843 765 19852 799
rect 19800 756 19852 765
rect 20168 756 20220 808
rect 20352 799 20404 808
rect 20352 765 20361 799
rect 20361 765 20395 799
rect 20395 765 20404 799
rect 20352 756 20404 765
rect 20536 824 20588 876
rect 21732 892 21784 944
rect 11428 620 11480 672
rect 11796 620 11848 672
rect 12164 620 12216 672
rect 12532 620 12584 672
rect 12900 620 12952 672
rect 13268 620 13320 672
rect 13728 620 13780 672
rect 14096 620 14148 672
rect 17684 663 17736 672
rect 17684 629 17693 663
rect 17693 629 17727 663
rect 17727 629 17736 663
rect 17684 620 17736 629
rect 18788 688 18840 740
rect 18144 620 18196 672
rect 18420 620 18472 672
rect 19524 688 19576 740
rect 20720 799 20772 808
rect 20720 765 20729 799
rect 20729 765 20763 799
rect 20763 765 20772 799
rect 20720 756 20772 765
rect 21916 756 21968 808
rect 22192 756 22244 808
rect 22468 756 22520 808
rect 23112 756 23164 808
rect 20628 620 20680 672
rect 21548 620 21600 672
rect 4366 518 4418 570
rect 4430 518 4482 570
rect 4494 518 4546 570
rect 4558 518 4610 570
rect 4622 518 4674 570
rect 4686 518 4738 570
rect 10366 518 10418 570
rect 10430 518 10482 570
rect 10494 518 10546 570
rect 10558 518 10610 570
rect 10622 518 10674 570
rect 10686 518 10738 570
rect 16366 518 16418 570
rect 16430 518 16482 570
rect 16494 518 16546 570
rect 16558 518 16610 570
rect 16622 518 16674 570
rect 16686 518 16738 570
rect 22366 518 22418 570
rect 22430 518 22482 570
rect 22494 518 22546 570
rect 22558 518 22610 570
rect 22622 518 22674 570
rect 22686 518 22738 570
rect 7196 416 7248 468
rect 9680 416 9732 468
rect 9864 416 9916 468
rect 10416 416 10468 468
rect 10600 416 10652 468
rect 11152 416 11204 468
rect 12072 416 12124 468
rect 1216 348 1268 400
rect 7748 348 7800 400
rect 3056 280 3108 332
rect 9312 348 9364 400
rect 10232 348 10284 400
rect 10784 348 10836 400
rect 17776 416 17828 468
rect 17868 416 17920 468
rect 18696 416 18748 468
rect 19800 416 19852 468
rect 19984 416 20036 468
rect 20444 416 20496 468
rect 12992 348 13044 400
rect 15108 348 15160 400
rect 17684 348 17736 400
rect 22192 348 22244 400
rect 8116 280 8168 332
rect 10048 280 10100 332
rect 3424 212 3476 264
rect 14280 280 14332 332
rect 14556 280 14608 332
rect 15568 280 15620 332
rect 18880 280 18932 332
rect 20904 280 20956 332
rect 11704 212 11756 264
rect 1952 144 2004 196
rect 4988 144 5040 196
rect 12992 144 13044 196
rect 9128 76 9180 128
rect 12072 76 12124 128
rect 16856 212 16908 264
rect 20812 212 20864 264
rect 18972 144 19024 196
rect 23388 144 23440 196
rect 12256 8 12308 60
rect 15200 76 15252 128
rect 20076 76 20128 128
rect 20168 8 20220 60
<< metal2 >>
rect 2228 23656 2280 23662
rect 2228 23598 2280 23604
rect 8298 23600 8354 24000
rect 8850 23600 8906 24000
rect 9402 23746 9458 24000
rect 9402 23718 9536 23746
rect 9402 23600 9458 23718
rect 2240 23186 2268 23598
rect 4160 23588 4212 23594
rect 4160 23530 4212 23536
rect 3056 23316 3108 23322
rect 3056 23258 3108 23264
rect 2228 23180 2280 23186
rect 2228 23122 2280 23128
rect 2412 23180 2464 23186
rect 2412 23122 2464 23128
rect 1768 22976 1820 22982
rect 1768 22918 1820 22924
rect 1364 22876 1740 22885
rect 1420 22874 1444 22876
rect 1500 22874 1524 22876
rect 1580 22874 1604 22876
rect 1660 22874 1684 22876
rect 1420 22822 1430 22874
rect 1674 22822 1684 22874
rect 1420 22820 1444 22822
rect 1500 22820 1524 22822
rect 1580 22820 1604 22822
rect 1660 22820 1684 22822
rect 1364 22811 1740 22820
rect 1780 22574 1808 22918
rect 1492 22568 1544 22574
rect 1492 22510 1544 22516
rect 1768 22568 1820 22574
rect 1768 22510 1820 22516
rect 1504 22234 1532 22510
rect 1768 22432 1820 22438
rect 1768 22374 1820 22380
rect 1492 22228 1544 22234
rect 1492 22170 1544 22176
rect 1364 21788 1740 21797
rect 1420 21786 1444 21788
rect 1500 21786 1524 21788
rect 1580 21786 1604 21788
rect 1660 21786 1684 21788
rect 1420 21734 1430 21786
rect 1674 21734 1684 21786
rect 1420 21732 1444 21734
rect 1500 21732 1524 21734
rect 1580 21732 1604 21734
rect 1660 21732 1684 21734
rect 1364 21723 1740 21732
rect 1364 20700 1740 20709
rect 1420 20698 1444 20700
rect 1500 20698 1524 20700
rect 1580 20698 1604 20700
rect 1660 20698 1684 20700
rect 1420 20646 1430 20698
rect 1674 20646 1684 20698
rect 1420 20644 1444 20646
rect 1500 20644 1524 20646
rect 1580 20644 1604 20646
rect 1660 20644 1684 20646
rect 1364 20635 1740 20644
rect 1400 20256 1452 20262
rect 1400 20198 1452 20204
rect 1412 19922 1440 20198
rect 1400 19916 1452 19922
rect 1400 19858 1452 19864
rect 1780 19854 1808 22374
rect 2240 22166 2268 23122
rect 2424 22234 2452 23122
rect 2964 22636 3016 22642
rect 2964 22578 3016 22584
rect 2976 22409 3004 22578
rect 2962 22400 3018 22409
rect 2962 22335 3018 22344
rect 2412 22228 2464 22234
rect 2412 22170 2464 22176
rect 2228 22160 2280 22166
rect 2228 22102 2280 22108
rect 1860 22092 1912 22098
rect 1860 22034 1912 22040
rect 2044 22092 2096 22098
rect 2044 22034 2096 22040
rect 2964 22092 3016 22098
rect 2964 22034 3016 22040
rect 1872 21690 1900 22034
rect 1952 21888 2004 21894
rect 1952 21830 2004 21836
rect 1860 21684 1912 21690
rect 1860 21626 1912 21632
rect 1964 21486 1992 21830
rect 1952 21480 2004 21486
rect 1952 21422 2004 21428
rect 2056 21350 2084 22034
rect 2228 22024 2280 22030
rect 2228 21966 2280 21972
rect 2872 22024 2924 22030
rect 2872 21966 2924 21972
rect 2136 21412 2188 21418
rect 2136 21354 2188 21360
rect 2044 21344 2096 21350
rect 2044 21286 2096 21292
rect 2148 21078 2176 21354
rect 2240 21146 2268 21966
rect 2780 21548 2832 21554
rect 2780 21490 2832 21496
rect 2504 21480 2556 21486
rect 2792 21457 2820 21490
rect 2504 21422 2556 21428
rect 2778 21448 2834 21457
rect 2516 21146 2544 21422
rect 2884 21418 2912 21966
rect 2976 21554 3004 22034
rect 3068 22030 3096 23258
rect 3240 23180 3292 23186
rect 3240 23122 3292 23128
rect 3332 23180 3384 23186
rect 3332 23122 3384 23128
rect 3056 22024 3108 22030
rect 3056 21966 3108 21972
rect 3252 21622 3280 23122
rect 3344 22234 3372 23122
rect 3976 22976 4028 22982
rect 3976 22918 4028 22924
rect 3988 22574 4016 22918
rect 4172 22574 4200 23530
rect 6092 23520 6144 23526
rect 6092 23462 6144 23468
rect 4364 23420 4740 23429
rect 4420 23418 4444 23420
rect 4500 23418 4524 23420
rect 4580 23418 4604 23420
rect 4660 23418 4684 23420
rect 4420 23366 4430 23418
rect 4674 23366 4684 23418
rect 4420 23364 4444 23366
rect 4500 23364 4524 23366
rect 4580 23364 4604 23366
rect 4660 23364 4684 23366
rect 4364 23355 4740 23364
rect 5448 23180 5500 23186
rect 5448 23122 5500 23128
rect 5724 23180 5776 23186
rect 5724 23122 5776 23128
rect 5080 23044 5132 23050
rect 5080 22986 5132 22992
rect 4896 22976 4948 22982
rect 4896 22918 4948 22924
rect 4804 22704 4856 22710
rect 4804 22646 4856 22652
rect 4252 22636 4304 22642
rect 4252 22578 4304 22584
rect 3700 22568 3752 22574
rect 3700 22510 3752 22516
rect 3976 22568 4028 22574
rect 3976 22510 4028 22516
rect 4160 22568 4212 22574
rect 4160 22510 4212 22516
rect 3332 22228 3384 22234
rect 3332 22170 3384 22176
rect 3712 22166 3740 22510
rect 3516 22160 3568 22166
rect 3516 22102 3568 22108
rect 3700 22160 3752 22166
rect 3700 22102 3752 22108
rect 3424 22092 3476 22098
rect 3424 22034 3476 22040
rect 3332 21888 3384 21894
rect 3332 21830 3384 21836
rect 3240 21616 3292 21622
rect 3240 21558 3292 21564
rect 2964 21548 3016 21554
rect 2964 21490 3016 21496
rect 3148 21480 3200 21486
rect 3148 21422 3200 21428
rect 2778 21383 2834 21392
rect 2872 21412 2924 21418
rect 2872 21354 2924 21360
rect 2596 21344 2648 21350
rect 2596 21286 2648 21292
rect 2228 21140 2280 21146
rect 2228 21082 2280 21088
rect 2504 21140 2556 21146
rect 2504 21082 2556 21088
rect 2136 21072 2188 21078
rect 2136 21014 2188 21020
rect 1860 21004 1912 21010
rect 1860 20946 1912 20952
rect 2228 21004 2280 21010
rect 2228 20946 2280 20952
rect 1872 20602 1900 20946
rect 1860 20596 1912 20602
rect 1860 20538 1912 20544
rect 1872 20398 1900 20538
rect 2134 20496 2190 20505
rect 2134 20431 2190 20440
rect 1860 20392 1912 20398
rect 2044 20392 2096 20398
rect 1860 20334 1912 20340
rect 2042 20360 2044 20369
rect 2096 20360 2098 20369
rect 2042 20295 2098 20304
rect 2044 20256 2096 20262
rect 2044 20198 2096 20204
rect 1952 20052 2004 20058
rect 1952 19994 2004 20000
rect 1768 19848 1820 19854
rect 1768 19790 1820 19796
rect 1364 19612 1740 19621
rect 1420 19610 1444 19612
rect 1500 19610 1524 19612
rect 1580 19610 1604 19612
rect 1660 19610 1684 19612
rect 1420 19558 1430 19610
rect 1674 19558 1684 19610
rect 1420 19556 1444 19558
rect 1500 19556 1524 19558
rect 1580 19556 1604 19558
rect 1660 19556 1684 19558
rect 1364 19547 1740 19556
rect 572 19372 624 19378
rect 572 19314 624 19320
rect 584 9518 612 19314
rect 1780 19310 1808 19790
rect 1860 19712 1912 19718
rect 1860 19654 1912 19660
rect 1872 19310 1900 19654
rect 1768 19304 1820 19310
rect 1768 19246 1820 19252
rect 1860 19304 1912 19310
rect 1964 19281 1992 19994
rect 2056 19922 2084 20198
rect 2044 19916 2096 19922
rect 2044 19858 2096 19864
rect 1860 19246 1912 19252
rect 1950 19272 2006 19281
rect 1950 19207 2006 19216
rect 1964 18766 1992 19207
rect 1952 18760 2004 18766
rect 1952 18702 2004 18708
rect 1364 18524 1740 18533
rect 1420 18522 1444 18524
rect 1500 18522 1524 18524
rect 1580 18522 1604 18524
rect 1660 18522 1684 18524
rect 1420 18470 1430 18522
rect 1674 18470 1684 18522
rect 1420 18468 1444 18470
rect 1500 18468 1524 18470
rect 1580 18468 1604 18470
rect 1660 18468 1684 18470
rect 1364 18459 1740 18468
rect 2148 18442 2176 20431
rect 2240 19310 2268 20946
rect 2504 20392 2556 20398
rect 2504 20334 2556 20340
rect 2516 19990 2544 20334
rect 2608 20330 2636 21286
rect 2780 21140 2832 21146
rect 2780 21082 2832 21088
rect 2792 20754 2820 21082
rect 2700 20726 2820 20754
rect 2700 20602 2728 20726
rect 2688 20596 2740 20602
rect 2688 20538 2740 20544
rect 2780 20392 2832 20398
rect 2780 20334 2832 20340
rect 2596 20324 2648 20330
rect 2596 20266 2648 20272
rect 2688 20256 2740 20262
rect 2688 20198 2740 20204
rect 2700 20058 2728 20198
rect 2688 20052 2740 20058
rect 2688 19994 2740 20000
rect 2504 19984 2556 19990
rect 2504 19926 2556 19932
rect 2516 19446 2544 19926
rect 2792 19922 2820 20334
rect 2884 19972 2912 21354
rect 2964 21344 3016 21350
rect 2964 21286 3016 21292
rect 2976 21078 3004 21286
rect 2964 21072 3016 21078
rect 2964 21014 3016 21020
rect 3160 20874 3188 21422
rect 3148 20868 3200 20874
rect 3148 20810 3200 20816
rect 3252 20466 3280 21558
rect 3344 21418 3372 21830
rect 3436 21690 3464 22034
rect 3424 21684 3476 21690
rect 3424 21626 3476 21632
rect 3332 21412 3384 21418
rect 3332 21354 3384 21360
rect 3528 21049 3556 22102
rect 3884 22094 3936 22098
rect 3988 22094 4016 22510
rect 4172 22094 4200 22510
rect 3884 22092 4016 22094
rect 3936 22066 4016 22092
rect 4080 22066 4200 22094
rect 3884 22034 3936 22040
rect 4080 22030 4108 22066
rect 4264 22030 4292 22578
rect 4364 22332 4740 22341
rect 4420 22330 4444 22332
rect 4500 22330 4524 22332
rect 4580 22330 4604 22332
rect 4660 22330 4684 22332
rect 4420 22278 4430 22330
rect 4674 22278 4684 22330
rect 4420 22276 4444 22278
rect 4500 22276 4524 22278
rect 4580 22276 4604 22278
rect 4660 22276 4684 22278
rect 4364 22267 4740 22276
rect 4816 22234 4844 22646
rect 4908 22574 4936 22918
rect 4896 22568 4948 22574
rect 4896 22510 4948 22516
rect 5092 22506 5120 22986
rect 5460 22982 5488 23122
rect 5540 23112 5592 23118
rect 5540 23054 5592 23060
rect 5448 22976 5500 22982
rect 5448 22918 5500 22924
rect 5080 22500 5132 22506
rect 5080 22442 5132 22448
rect 4804 22228 4856 22234
rect 4804 22170 4856 22176
rect 4712 22092 4764 22098
rect 4712 22034 4764 22040
rect 4068 22024 4120 22030
rect 4068 21966 4120 21972
rect 4252 22024 4304 22030
rect 4252 21966 4304 21972
rect 4724 21894 4752 22034
rect 5092 21962 5120 22442
rect 5264 22432 5316 22438
rect 5264 22374 5316 22380
rect 5356 22432 5408 22438
rect 5356 22374 5408 22380
rect 5276 22098 5304 22374
rect 5368 22137 5396 22374
rect 5460 22234 5488 22918
rect 5552 22778 5580 23054
rect 5736 22778 5764 23122
rect 5540 22772 5592 22778
rect 5540 22714 5592 22720
rect 5724 22772 5776 22778
rect 5724 22714 5776 22720
rect 5632 22704 5684 22710
rect 5632 22646 5684 22652
rect 5540 22500 5592 22506
rect 5540 22442 5592 22448
rect 5552 22234 5580 22442
rect 5448 22228 5500 22234
rect 5448 22170 5500 22176
rect 5540 22228 5592 22234
rect 5540 22170 5592 22176
rect 5354 22128 5410 22137
rect 5172 22092 5224 22098
rect 5172 22034 5224 22040
rect 5264 22092 5316 22098
rect 5354 22063 5410 22072
rect 5448 22092 5500 22098
rect 5264 22034 5316 22040
rect 5644 22080 5672 22646
rect 6104 22642 6132 23462
rect 8312 23322 8340 23600
rect 8300 23316 8352 23322
rect 8300 23258 8352 23264
rect 6736 23180 6788 23186
rect 6736 23122 6788 23128
rect 8208 23180 8260 23186
rect 8208 23122 8260 23128
rect 6368 23112 6420 23118
rect 6368 23054 6420 23060
rect 6092 22636 6144 22642
rect 6092 22578 6144 22584
rect 6104 22506 6132 22578
rect 6092 22500 6144 22506
rect 6092 22442 6144 22448
rect 6184 22432 6236 22438
rect 6184 22374 6236 22380
rect 5500 22052 5672 22080
rect 5448 22034 5500 22040
rect 5080 21956 5132 21962
rect 5080 21898 5132 21904
rect 3884 21888 3936 21894
rect 3884 21830 3936 21836
rect 4712 21888 4764 21894
rect 4712 21830 4764 21836
rect 4896 21888 4948 21894
rect 4896 21830 4948 21836
rect 3896 21593 3924 21830
rect 3882 21584 3938 21593
rect 4908 21554 4936 21830
rect 5184 21690 5212 22034
rect 5816 21956 5868 21962
rect 5816 21898 5868 21904
rect 5172 21684 5224 21690
rect 5172 21626 5224 21632
rect 5264 21616 5316 21622
rect 5264 21558 5316 21564
rect 3882 21519 3938 21528
rect 4896 21548 4948 21554
rect 3896 21486 3924 21519
rect 4896 21490 4948 21496
rect 3884 21480 3936 21486
rect 3884 21422 3936 21428
rect 4252 21480 4304 21486
rect 4252 21422 4304 21428
rect 5172 21480 5224 21486
rect 5172 21422 5224 21428
rect 3514 21040 3570 21049
rect 3514 20975 3516 20984
rect 3568 20975 3570 20984
rect 3516 20946 3568 20952
rect 4160 20936 4212 20942
rect 4066 20904 4122 20913
rect 4264 20890 4292 21422
rect 4896 21344 4948 21350
rect 4896 21286 4948 21292
rect 5080 21344 5132 21350
rect 5080 21286 5132 21292
rect 4364 21244 4740 21253
rect 4420 21242 4444 21244
rect 4500 21242 4524 21244
rect 4580 21242 4604 21244
rect 4660 21242 4684 21244
rect 4420 21190 4430 21242
rect 4674 21190 4684 21242
rect 4420 21188 4444 21190
rect 4500 21188 4524 21190
rect 4580 21188 4604 21190
rect 4660 21188 4684 21190
rect 4364 21179 4740 21188
rect 4908 21078 4936 21286
rect 4986 21176 5042 21185
rect 4986 21111 5042 21120
rect 4344 21072 4396 21078
rect 4344 21014 4396 21020
rect 4896 21072 4948 21078
rect 4896 21014 4948 21020
rect 4212 20884 4292 20890
rect 4160 20878 4292 20884
rect 4172 20862 4292 20878
rect 4066 20839 4122 20848
rect 4080 20806 4108 20839
rect 4068 20800 4120 20806
rect 4068 20742 4120 20748
rect 3240 20460 3292 20466
rect 3240 20402 3292 20408
rect 2964 19984 3016 19990
rect 2884 19944 2964 19972
rect 2964 19926 3016 19932
rect 2780 19916 2832 19922
rect 2780 19858 2832 19864
rect 2504 19440 2556 19446
rect 2504 19382 2556 19388
rect 2228 19304 2280 19310
rect 2228 19246 2280 19252
rect 2412 19304 2464 19310
rect 2412 19246 2464 19252
rect 2240 19145 2268 19246
rect 2226 19136 2282 19145
rect 2226 19071 2282 19080
rect 2424 18834 2452 19246
rect 2976 19242 3004 19926
rect 3252 19922 3280 20402
rect 4080 20398 4108 20742
rect 4068 20392 4120 20398
rect 4068 20334 4120 20340
rect 4264 19990 4292 20862
rect 4356 20262 4384 21014
rect 5000 21010 5028 21111
rect 4620 21004 4672 21010
rect 4620 20946 4672 20952
rect 4712 21004 4764 21010
rect 4712 20946 4764 20952
rect 4988 21004 5040 21010
rect 4988 20946 5040 20952
rect 4632 20466 4660 20946
rect 4724 20913 4752 20946
rect 4804 20936 4856 20942
rect 4710 20904 4766 20913
rect 4804 20878 4856 20884
rect 4710 20839 4766 20848
rect 4620 20460 4672 20466
rect 4620 20402 4672 20408
rect 4344 20256 4396 20262
rect 4344 20198 4396 20204
rect 4364 20156 4740 20165
rect 4420 20154 4444 20156
rect 4500 20154 4524 20156
rect 4580 20154 4604 20156
rect 4660 20154 4684 20156
rect 4420 20102 4430 20154
rect 4674 20102 4684 20154
rect 4420 20100 4444 20102
rect 4500 20100 4524 20102
rect 4580 20100 4604 20102
rect 4660 20100 4684 20102
rect 4364 20091 4740 20100
rect 4816 20058 4844 20878
rect 4988 20868 5040 20874
rect 4988 20810 5040 20816
rect 4896 20460 4948 20466
rect 4896 20402 4948 20408
rect 4804 20052 4856 20058
rect 4804 19994 4856 20000
rect 4252 19984 4304 19990
rect 4252 19926 4304 19932
rect 3240 19916 3292 19922
rect 3240 19858 3292 19864
rect 3424 19916 3476 19922
rect 3424 19858 3476 19864
rect 2964 19236 3016 19242
rect 2964 19178 3016 19184
rect 3056 19168 3108 19174
rect 3056 19110 3108 19116
rect 3068 18970 3096 19110
rect 3252 18970 3280 19858
rect 3436 19514 3464 19858
rect 3516 19712 3568 19718
rect 3516 19654 3568 19660
rect 4528 19712 4580 19718
rect 4528 19654 4580 19660
rect 3332 19508 3384 19514
rect 3332 19450 3384 19456
rect 3424 19508 3476 19514
rect 3424 19450 3476 19456
rect 3344 19394 3372 19450
rect 3422 19408 3478 19417
rect 3344 19366 3422 19394
rect 3422 19343 3478 19352
rect 3436 19310 3464 19343
rect 3528 19310 3556 19654
rect 4540 19310 4568 19654
rect 3424 19304 3476 19310
rect 3424 19246 3476 19252
rect 3516 19304 3568 19310
rect 3516 19246 3568 19252
rect 3792 19304 3844 19310
rect 3792 19246 3844 19252
rect 3976 19304 4028 19310
rect 4068 19304 4120 19310
rect 3976 19246 4028 19252
rect 4066 19272 4068 19281
rect 4528 19304 4580 19310
rect 4120 19272 4122 19281
rect 3804 19145 3832 19246
rect 3790 19136 3846 19145
rect 3790 19071 3846 19080
rect 3988 18970 4016 19246
rect 4528 19246 4580 19252
rect 4066 19207 4122 19216
rect 4252 19168 4304 19174
rect 4252 19110 4304 19116
rect 4804 19168 4856 19174
rect 4804 19110 4856 19116
rect 3056 18964 3108 18970
rect 3056 18906 3108 18912
rect 3240 18964 3292 18970
rect 3240 18906 3292 18912
rect 3976 18964 4028 18970
rect 3976 18906 4028 18912
rect 2412 18828 2464 18834
rect 2412 18770 2464 18776
rect 4264 18766 4292 19110
rect 4364 19068 4740 19077
rect 4420 19066 4444 19068
rect 4500 19066 4524 19068
rect 4580 19066 4604 19068
rect 4660 19066 4684 19068
rect 4420 19014 4430 19066
rect 4674 19014 4684 19066
rect 4420 19012 4444 19014
rect 4500 19012 4524 19014
rect 4580 19012 4604 19014
rect 4660 19012 4684 19014
rect 4364 19003 4740 19012
rect 4816 18766 4844 19110
rect 4908 18902 4936 20402
rect 5000 19854 5028 20810
rect 5092 19922 5120 21286
rect 5080 19916 5132 19922
rect 5080 19858 5132 19864
rect 4988 19848 5040 19854
rect 4988 19790 5040 19796
rect 5000 19514 5028 19790
rect 4988 19508 5040 19514
rect 4988 19450 5040 19456
rect 4896 18896 4948 18902
rect 4896 18838 4948 18844
rect 5000 18834 5028 19450
rect 5184 19174 5212 21422
rect 5276 21010 5304 21558
rect 5632 21480 5684 21486
rect 5632 21422 5684 21428
rect 5644 21146 5672 21422
rect 5828 21350 5856 21898
rect 6196 21894 6224 22374
rect 6184 21888 6236 21894
rect 6184 21830 6236 21836
rect 5908 21684 5960 21690
rect 5908 21626 5960 21632
rect 5920 21350 5948 21626
rect 6196 21486 6224 21830
rect 6184 21480 6236 21486
rect 6184 21422 6236 21428
rect 5816 21344 5868 21350
rect 5816 21286 5868 21292
rect 5908 21344 5960 21350
rect 5908 21286 5960 21292
rect 5632 21140 5684 21146
rect 5632 21082 5684 21088
rect 5264 21004 5316 21010
rect 5264 20946 5316 20952
rect 5540 21004 5592 21010
rect 5540 20946 5592 20952
rect 5816 21004 5868 21010
rect 5816 20946 5868 20952
rect 5276 20058 5304 20946
rect 5552 20534 5580 20946
rect 5540 20528 5592 20534
rect 5540 20470 5592 20476
rect 5540 20324 5592 20330
rect 5540 20266 5592 20272
rect 5356 20256 5408 20262
rect 5356 20198 5408 20204
rect 5264 20052 5316 20058
rect 5264 19994 5316 20000
rect 5276 19446 5304 19994
rect 5368 19990 5396 20198
rect 5356 19984 5408 19990
rect 5356 19926 5408 19932
rect 5446 19952 5502 19961
rect 5446 19887 5448 19896
rect 5500 19887 5502 19896
rect 5448 19858 5500 19864
rect 5460 19514 5488 19858
rect 5552 19514 5580 20266
rect 5828 20058 5856 20946
rect 5816 20052 5868 20058
rect 5816 19994 5868 20000
rect 5920 19854 5948 21286
rect 6090 21040 6146 21049
rect 6090 20975 6092 20984
rect 6144 20975 6146 20984
rect 6092 20946 6144 20952
rect 6196 20806 6224 21422
rect 6276 21140 6328 21146
rect 6276 21082 6328 21088
rect 6288 20913 6316 21082
rect 6274 20904 6330 20913
rect 6274 20839 6330 20848
rect 6184 20800 6236 20806
rect 6184 20742 6236 20748
rect 6380 20602 6408 23054
rect 6748 22778 6776 23122
rect 8116 22976 8168 22982
rect 8116 22918 8168 22924
rect 7364 22876 7740 22885
rect 7420 22874 7444 22876
rect 7500 22874 7524 22876
rect 7580 22874 7604 22876
rect 7660 22874 7684 22876
rect 7420 22822 7430 22874
rect 7674 22822 7684 22874
rect 7420 22820 7444 22822
rect 7500 22820 7524 22822
rect 7580 22820 7604 22822
rect 7660 22820 7684 22822
rect 7364 22811 7740 22820
rect 6736 22772 6788 22778
rect 6736 22714 6788 22720
rect 8128 22642 8156 22918
rect 7840 22636 7892 22642
rect 7840 22578 7892 22584
rect 8116 22636 8168 22642
rect 8116 22578 8168 22584
rect 7288 22568 7340 22574
rect 7288 22510 7340 22516
rect 7196 22432 7248 22438
rect 7196 22374 7248 22380
rect 7208 22234 7236 22374
rect 7196 22228 7248 22234
rect 7196 22170 7248 22176
rect 6460 22160 6512 22166
rect 6460 22102 6512 22108
rect 6472 22030 6500 22102
rect 7196 22092 7248 22098
rect 7196 22034 7248 22040
rect 6460 22024 6512 22030
rect 6460 21966 6512 21972
rect 6552 21888 6604 21894
rect 6552 21830 6604 21836
rect 7104 21888 7156 21894
rect 7104 21830 7156 21836
rect 6460 21004 6512 21010
rect 6460 20946 6512 20952
rect 6368 20596 6420 20602
rect 6368 20538 6420 20544
rect 6184 20324 6236 20330
rect 6184 20266 6236 20272
rect 6196 20058 6224 20266
rect 6184 20052 6236 20058
rect 6184 19994 6236 20000
rect 6184 19916 6236 19922
rect 6184 19858 6236 19864
rect 5908 19848 5960 19854
rect 5908 19790 5960 19796
rect 5448 19508 5500 19514
rect 5448 19450 5500 19456
rect 5540 19508 5592 19514
rect 5540 19450 5592 19456
rect 5264 19440 5316 19446
rect 5264 19382 5316 19388
rect 5172 19168 5224 19174
rect 5172 19110 5224 19116
rect 5184 18834 5212 19110
rect 5264 18896 5316 18902
rect 5264 18838 5316 18844
rect 4988 18828 5040 18834
rect 4988 18770 5040 18776
rect 5172 18828 5224 18834
rect 5172 18770 5224 18776
rect 2596 18760 2648 18766
rect 2596 18702 2648 18708
rect 4252 18760 4304 18766
rect 4252 18702 4304 18708
rect 4804 18760 4856 18766
rect 4804 18702 4856 18708
rect 1872 18414 2176 18442
rect 2320 18420 2372 18426
rect 1768 18080 1820 18086
rect 1768 18022 1820 18028
rect 1216 17740 1268 17746
rect 1216 17682 1268 17688
rect 848 17672 900 17678
rect 848 17614 900 17620
rect 860 16658 888 17614
rect 1228 17338 1256 17682
rect 1364 17436 1740 17445
rect 1420 17434 1444 17436
rect 1500 17434 1524 17436
rect 1580 17434 1604 17436
rect 1660 17434 1684 17436
rect 1420 17382 1430 17434
rect 1674 17382 1684 17434
rect 1420 17380 1444 17382
rect 1500 17380 1524 17382
rect 1580 17380 1604 17382
rect 1660 17380 1684 17382
rect 1364 17371 1740 17380
rect 1216 17332 1268 17338
rect 1216 17274 1268 17280
rect 1780 17218 1808 18022
rect 1688 17190 1808 17218
rect 1688 17134 1716 17190
rect 1676 17128 1728 17134
rect 1676 17070 1728 17076
rect 1124 16992 1176 16998
rect 1124 16934 1176 16940
rect 848 16652 900 16658
rect 848 16594 900 16600
rect 860 16114 888 16594
rect 848 16108 900 16114
rect 848 16050 900 16056
rect 1136 16046 1164 16934
rect 1364 16348 1740 16357
rect 1420 16346 1444 16348
rect 1500 16346 1524 16348
rect 1580 16346 1604 16348
rect 1660 16346 1684 16348
rect 1420 16294 1430 16346
rect 1674 16294 1684 16346
rect 1420 16292 1444 16294
rect 1500 16292 1524 16294
rect 1580 16292 1604 16294
rect 1660 16292 1684 16294
rect 1364 16283 1740 16292
rect 1124 16040 1176 16046
rect 1124 15982 1176 15988
rect 1214 16008 1270 16017
rect 1214 15943 1270 15952
rect 1228 15638 1256 15943
rect 1872 15722 1900 18414
rect 2320 18362 2372 18368
rect 2044 18352 2096 18358
rect 2044 18294 2096 18300
rect 1952 18216 2004 18222
rect 1952 18158 2004 18164
rect 1964 17134 1992 18158
rect 2056 17134 2084 18294
rect 2228 18148 2280 18154
rect 2228 18090 2280 18096
rect 1952 17128 2004 17134
rect 1952 17070 2004 17076
rect 2044 17128 2096 17134
rect 2044 17070 2096 17076
rect 2240 16674 2268 18090
rect 2332 17882 2360 18362
rect 2320 17876 2372 17882
rect 2320 17818 2372 17824
rect 2504 17536 2556 17542
rect 2504 17478 2556 17484
rect 2516 17338 2544 17478
rect 2504 17332 2556 17338
rect 2504 17274 2556 17280
rect 2516 17066 2544 17274
rect 2504 17060 2556 17066
rect 2504 17002 2556 17008
rect 2410 16688 2466 16697
rect 2240 16646 2410 16674
rect 2410 16623 2412 16632
rect 2464 16623 2466 16632
rect 2504 16652 2556 16658
rect 2412 16594 2464 16600
rect 2504 16594 2556 16600
rect 2516 16561 2544 16594
rect 2502 16552 2558 16561
rect 2502 16487 2558 16496
rect 2320 16448 2372 16454
rect 2320 16390 2372 16396
rect 2332 16250 2360 16390
rect 2320 16244 2372 16250
rect 2320 16186 2372 16192
rect 1872 15694 2176 15722
rect 940 15632 992 15638
rect 940 15574 992 15580
rect 1216 15632 1268 15638
rect 1216 15574 1268 15580
rect 848 13864 900 13870
rect 848 13806 900 13812
rect 860 13394 888 13806
rect 848 13388 900 13394
rect 848 13330 900 13336
rect 860 12986 888 13330
rect 848 12980 900 12986
rect 848 12922 900 12928
rect 756 12912 808 12918
rect 756 12854 808 12860
rect 664 12844 716 12850
rect 664 12786 716 12792
rect 572 9512 624 9518
rect 572 9454 624 9460
rect 676 4690 704 12786
rect 768 11694 796 12854
rect 848 12164 900 12170
rect 848 12106 900 12112
rect 756 11688 808 11694
rect 756 11630 808 11636
rect 860 11626 888 12106
rect 952 11830 980 15574
rect 1676 15564 1728 15570
rect 1952 15564 2004 15570
rect 1728 15524 1808 15552
rect 1676 15506 1728 15512
rect 1364 15260 1740 15269
rect 1420 15258 1444 15260
rect 1500 15258 1524 15260
rect 1580 15258 1604 15260
rect 1660 15258 1684 15260
rect 1420 15206 1430 15258
rect 1674 15206 1684 15258
rect 1420 15204 1444 15206
rect 1500 15204 1524 15206
rect 1580 15204 1604 15206
rect 1660 15204 1684 15206
rect 1364 15195 1740 15204
rect 1216 14952 1268 14958
rect 1216 14894 1268 14900
rect 1032 14476 1084 14482
rect 1032 14418 1084 14424
rect 1124 14476 1176 14482
rect 1124 14418 1176 14424
rect 1044 13802 1072 14418
rect 1136 13870 1164 14418
rect 1228 13870 1256 14894
rect 1584 14816 1636 14822
rect 1584 14758 1636 14764
rect 1596 14482 1624 14758
rect 1780 14550 1808 15524
rect 1952 15506 2004 15512
rect 1860 15428 1912 15434
rect 1860 15370 1912 15376
rect 1872 14618 1900 15370
rect 1964 14822 1992 15506
rect 1952 14816 2004 14822
rect 1952 14758 2004 14764
rect 1860 14612 1912 14618
rect 1860 14554 1912 14560
rect 1768 14544 1820 14550
rect 1768 14486 1820 14492
rect 1584 14476 1636 14482
rect 1584 14418 1636 14424
rect 1364 14172 1740 14181
rect 1420 14170 1444 14172
rect 1500 14170 1524 14172
rect 1580 14170 1604 14172
rect 1660 14170 1684 14172
rect 1420 14118 1430 14170
rect 1674 14118 1684 14170
rect 1420 14116 1444 14118
rect 1500 14116 1524 14118
rect 1580 14116 1604 14118
rect 1660 14116 1684 14118
rect 1364 14107 1740 14116
rect 1124 13864 1176 13870
rect 1124 13806 1176 13812
rect 1216 13864 1268 13870
rect 1216 13806 1268 13812
rect 1032 13796 1084 13802
rect 1032 13738 1084 13744
rect 1124 13456 1176 13462
rect 1124 13398 1176 13404
rect 1032 12776 1084 12782
rect 1032 12718 1084 12724
rect 1044 12442 1072 12718
rect 1032 12436 1084 12442
rect 1032 12378 1084 12384
rect 1044 12170 1072 12378
rect 1032 12164 1084 12170
rect 1032 12106 1084 12112
rect 940 11824 992 11830
rect 940 11766 992 11772
rect 1136 11762 1164 13398
rect 1228 12306 1256 13806
rect 1308 13728 1360 13734
rect 1308 13670 1360 13676
rect 1320 13530 1348 13670
rect 1308 13524 1360 13530
rect 1308 13466 1360 13472
rect 1780 13394 1808 14486
rect 2044 14476 2096 14482
rect 2044 14418 2096 14424
rect 1860 14272 1912 14278
rect 1860 14214 1912 14220
rect 1872 13870 1900 14214
rect 1860 13864 1912 13870
rect 1860 13806 1912 13812
rect 2056 13530 2084 14418
rect 2044 13524 2096 13530
rect 2044 13466 2096 13472
rect 1768 13388 1820 13394
rect 1768 13330 1820 13336
rect 2148 13190 2176 15694
rect 2332 15570 2360 16186
rect 2608 16153 2636 18702
rect 4896 18624 4948 18630
rect 4896 18566 4948 18572
rect 3976 18420 4028 18426
rect 3976 18362 4028 18368
rect 2964 18284 3016 18290
rect 2964 18226 3016 18232
rect 2780 18216 2832 18222
rect 2780 18158 2832 18164
rect 2688 18148 2740 18154
rect 2688 18090 2740 18096
rect 2700 17882 2728 18090
rect 2688 17876 2740 17882
rect 2688 17818 2740 17824
rect 2688 17672 2740 17678
rect 2686 17640 2688 17649
rect 2740 17640 2742 17649
rect 2686 17575 2742 17584
rect 2792 17338 2820 18158
rect 2872 17740 2924 17746
rect 2872 17682 2924 17688
rect 2884 17338 2912 17682
rect 2780 17332 2832 17338
rect 2700 17292 2780 17320
rect 2700 16658 2728 17292
rect 2780 17274 2832 17280
rect 2872 17332 2924 17338
rect 2872 17274 2924 17280
rect 2976 17134 3004 18226
rect 3056 18080 3108 18086
rect 3056 18022 3108 18028
rect 3884 18080 3936 18086
rect 3884 18022 3936 18028
rect 3068 17746 3096 18022
rect 3896 17814 3924 18022
rect 3884 17808 3936 17814
rect 3884 17750 3936 17756
rect 3056 17740 3108 17746
rect 3056 17682 3108 17688
rect 3884 17672 3936 17678
rect 3620 17598 3832 17626
rect 3884 17614 3936 17620
rect 3056 17332 3108 17338
rect 3056 17274 3108 17280
rect 2872 17128 2924 17134
rect 2872 17070 2924 17076
rect 2964 17128 3016 17134
rect 3068 17105 3096 17274
rect 3620 17202 3648 17598
rect 3804 17542 3832 17598
rect 3700 17536 3752 17542
rect 3700 17478 3752 17484
rect 3792 17536 3844 17542
rect 3792 17478 3844 17484
rect 3608 17196 3660 17202
rect 3608 17138 3660 17144
rect 2964 17070 3016 17076
rect 3054 17096 3110 17105
rect 2884 16998 2912 17070
rect 3054 17031 3110 17040
rect 3712 16998 3740 17478
rect 3790 17232 3846 17241
rect 3790 17167 3846 17176
rect 2872 16992 2924 16998
rect 2872 16934 2924 16940
rect 3700 16992 3752 16998
rect 3700 16934 3752 16940
rect 3712 16726 3740 16934
rect 3700 16720 3752 16726
rect 3804 16697 3832 17167
rect 3896 16794 3924 17614
rect 3988 16794 4016 18362
rect 4908 18358 4936 18566
rect 4896 18352 4948 18358
rect 4896 18294 4948 18300
rect 5078 18320 5134 18329
rect 4160 18284 4212 18290
rect 5184 18290 5212 18770
rect 5276 18698 5304 18838
rect 5264 18692 5316 18698
rect 5264 18634 5316 18640
rect 5448 18692 5500 18698
rect 5448 18634 5500 18640
rect 5078 18255 5134 18264
rect 5172 18284 5224 18290
rect 4160 18226 4212 18232
rect 4068 18216 4120 18222
rect 4066 18184 4068 18193
rect 4120 18184 4122 18193
rect 4066 18119 4122 18128
rect 3884 16788 3936 16794
rect 3884 16730 3936 16736
rect 3976 16788 4028 16794
rect 3976 16730 4028 16736
rect 3700 16662 3752 16668
rect 3790 16688 3846 16697
rect 2688 16652 2740 16658
rect 3516 16652 3568 16658
rect 2740 16612 2820 16640
rect 2688 16594 2740 16600
rect 2688 16448 2740 16454
rect 2688 16390 2740 16396
rect 2594 16144 2650 16153
rect 2700 16114 2728 16390
rect 2594 16079 2650 16088
rect 2688 16108 2740 16114
rect 2608 15994 2636 16079
rect 2688 16050 2740 16056
rect 2792 16046 2820 16612
rect 3516 16594 3568 16600
rect 3608 16652 3660 16658
rect 3790 16623 3792 16632
rect 3608 16594 3660 16600
rect 3844 16623 3846 16632
rect 3792 16594 3844 16600
rect 3528 16561 3556 16594
rect 2962 16552 3018 16561
rect 3514 16552 3570 16561
rect 2962 16487 3018 16496
rect 3332 16516 3384 16522
rect 2872 16176 2924 16182
rect 2872 16118 2924 16124
rect 2424 15966 2636 15994
rect 2780 16040 2832 16046
rect 2780 15982 2832 15988
rect 2320 15564 2372 15570
rect 2320 15506 2372 15512
rect 2424 14414 2452 15966
rect 2504 15904 2556 15910
rect 2504 15846 2556 15852
rect 2780 15904 2832 15910
rect 2780 15846 2832 15852
rect 2516 15162 2544 15846
rect 2792 15638 2820 15846
rect 2780 15632 2832 15638
rect 2780 15574 2832 15580
rect 2884 15473 2912 16118
rect 2976 15706 3004 16487
rect 3514 16487 3570 16496
rect 3332 16458 3384 16464
rect 3056 16108 3108 16114
rect 3056 16050 3108 16056
rect 2964 15700 3016 15706
rect 2964 15642 3016 15648
rect 2870 15464 2926 15473
rect 2870 15399 2926 15408
rect 3068 15366 3096 16050
rect 3344 16046 3372 16458
rect 3240 16040 3292 16046
rect 3240 15982 3292 15988
rect 3332 16040 3384 16046
rect 3332 15982 3384 15988
rect 3252 15638 3280 15982
rect 3240 15632 3292 15638
rect 3240 15574 3292 15580
rect 3148 15428 3200 15434
rect 3148 15370 3200 15376
rect 3056 15360 3108 15366
rect 3056 15302 3108 15308
rect 2504 15156 2556 15162
rect 2504 15098 2556 15104
rect 2516 15026 2544 15098
rect 2504 15020 2556 15026
rect 2504 14962 2556 14968
rect 2872 15020 2924 15026
rect 2872 14962 2924 14968
rect 2596 14952 2648 14958
rect 2596 14894 2648 14900
rect 2608 14550 2636 14894
rect 2596 14544 2648 14550
rect 2596 14486 2648 14492
rect 2884 14414 2912 14962
rect 3160 14482 3188 15370
rect 3252 15094 3280 15574
rect 3620 15570 3648 16594
rect 3792 16448 3844 16454
rect 3792 16390 3844 16396
rect 3804 15706 3832 16390
rect 3792 15700 3844 15706
rect 3792 15642 3844 15648
rect 3608 15564 3660 15570
rect 3608 15506 3660 15512
rect 3332 15496 3384 15502
rect 3330 15464 3332 15473
rect 3384 15464 3386 15473
rect 3330 15399 3386 15408
rect 3240 15088 3292 15094
rect 3240 15030 3292 15036
rect 3424 14884 3476 14890
rect 3424 14826 3476 14832
rect 3884 14884 3936 14890
rect 3884 14826 3936 14832
rect 3436 14618 3464 14826
rect 3700 14816 3752 14822
rect 3700 14758 3752 14764
rect 3792 14816 3844 14822
rect 3792 14758 3844 14764
rect 3424 14612 3476 14618
rect 3424 14554 3476 14560
rect 3712 14550 3740 14758
rect 3700 14544 3752 14550
rect 3700 14486 3752 14492
rect 2964 14476 3016 14482
rect 2964 14418 3016 14424
rect 3148 14476 3200 14482
rect 3148 14418 3200 14424
rect 2412 14408 2464 14414
rect 2412 14350 2464 14356
rect 2872 14408 2924 14414
rect 2872 14350 2924 14356
rect 2976 14074 3004 14418
rect 3516 14340 3568 14346
rect 3516 14282 3568 14288
rect 3148 14272 3200 14278
rect 3148 14214 3200 14220
rect 2964 14068 3016 14074
rect 2964 14010 3016 14016
rect 2688 14000 2740 14006
rect 2688 13942 2740 13948
rect 2412 13796 2464 13802
rect 2412 13738 2464 13744
rect 2424 13394 2452 13738
rect 2596 13728 2648 13734
rect 2596 13670 2648 13676
rect 2608 13530 2636 13670
rect 2596 13524 2648 13530
rect 2596 13466 2648 13472
rect 2412 13388 2464 13394
rect 2412 13330 2464 13336
rect 2504 13320 2556 13326
rect 2504 13262 2556 13268
rect 1768 13184 1820 13190
rect 1768 13126 1820 13132
rect 2136 13184 2188 13190
rect 2136 13126 2188 13132
rect 1364 13084 1740 13093
rect 1420 13082 1444 13084
rect 1500 13082 1524 13084
rect 1580 13082 1604 13084
rect 1660 13082 1684 13084
rect 1420 13030 1430 13082
rect 1674 13030 1684 13082
rect 1420 13028 1444 13030
rect 1500 13028 1524 13030
rect 1580 13028 1604 13030
rect 1660 13028 1684 13030
rect 1364 13019 1740 13028
rect 1676 12912 1728 12918
rect 1676 12854 1728 12860
rect 1492 12708 1544 12714
rect 1492 12650 1544 12656
rect 1216 12300 1268 12306
rect 1216 12242 1268 12248
rect 1124 11756 1176 11762
rect 1124 11698 1176 11704
rect 848 11620 900 11626
rect 1124 11620 1176 11626
rect 848 11562 900 11568
rect 1044 11580 1124 11608
rect 940 11552 992 11558
rect 940 11494 992 11500
rect 848 11144 900 11150
rect 848 11086 900 11092
rect 860 10130 888 11086
rect 952 10606 980 11494
rect 1044 10742 1072 11580
rect 1124 11562 1176 11568
rect 1228 11506 1256 12242
rect 1504 12209 1532 12650
rect 1688 12374 1716 12854
rect 1780 12434 1808 13126
rect 2044 12776 2096 12782
rect 2044 12718 2096 12724
rect 1952 12640 2004 12646
rect 1952 12582 2004 12588
rect 1964 12442 1992 12582
rect 1952 12436 2004 12442
rect 1780 12406 1900 12434
rect 1676 12368 1728 12374
rect 1728 12328 1808 12356
rect 1676 12310 1728 12316
rect 1490 12200 1546 12209
rect 1490 12135 1546 12144
rect 1364 11996 1740 12005
rect 1420 11994 1444 11996
rect 1500 11994 1524 11996
rect 1580 11994 1604 11996
rect 1660 11994 1684 11996
rect 1420 11942 1430 11994
rect 1674 11942 1684 11994
rect 1420 11940 1444 11942
rect 1500 11940 1524 11942
rect 1580 11940 1604 11942
rect 1660 11940 1684 11942
rect 1364 11931 1740 11940
rect 1780 11880 1808 12328
rect 1596 11852 1808 11880
rect 1308 11824 1360 11830
rect 1308 11766 1360 11772
rect 1320 11626 1348 11766
rect 1596 11762 1624 11852
rect 1584 11756 1636 11762
rect 1584 11698 1636 11704
rect 1676 11756 1728 11762
rect 1676 11698 1728 11704
rect 1308 11620 1360 11626
rect 1308 11562 1360 11568
rect 1136 11478 1256 11506
rect 1136 11218 1164 11478
rect 1688 11354 1716 11698
rect 1768 11620 1820 11626
rect 1768 11562 1820 11568
rect 1676 11348 1728 11354
rect 1676 11290 1728 11296
rect 1124 11212 1176 11218
rect 1124 11154 1176 11160
rect 1308 11212 1360 11218
rect 1308 11154 1360 11160
rect 1320 10996 1348 11154
rect 1228 10968 1348 10996
rect 1228 10810 1256 10968
rect 1364 10908 1740 10917
rect 1420 10906 1444 10908
rect 1500 10906 1524 10908
rect 1580 10906 1604 10908
rect 1660 10906 1684 10908
rect 1420 10854 1430 10906
rect 1674 10854 1684 10906
rect 1420 10852 1444 10854
rect 1500 10852 1524 10854
rect 1580 10852 1604 10854
rect 1660 10852 1684 10854
rect 1364 10843 1740 10852
rect 1780 10810 1808 11562
rect 1216 10804 1268 10810
rect 1216 10746 1268 10752
rect 1768 10804 1820 10810
rect 1768 10746 1820 10752
rect 1032 10736 1084 10742
rect 1032 10678 1084 10684
rect 940 10600 992 10606
rect 940 10542 992 10548
rect 848 10124 900 10130
rect 848 10066 900 10072
rect 1124 10124 1176 10130
rect 1124 10066 1176 10072
rect 1136 9178 1164 10066
rect 1364 9820 1740 9829
rect 1420 9818 1444 9820
rect 1500 9818 1524 9820
rect 1580 9818 1604 9820
rect 1660 9818 1684 9820
rect 1420 9766 1430 9818
rect 1674 9766 1684 9818
rect 1420 9764 1444 9766
rect 1500 9764 1524 9766
rect 1580 9764 1604 9766
rect 1660 9764 1684 9766
rect 1364 9755 1740 9764
rect 1676 9648 1728 9654
rect 1676 9590 1728 9596
rect 1400 9512 1452 9518
rect 1398 9480 1400 9489
rect 1452 9480 1454 9489
rect 1228 9438 1398 9466
rect 1124 9172 1176 9178
rect 1124 9114 1176 9120
rect 1124 9036 1176 9042
rect 1124 8978 1176 8984
rect 1032 8968 1084 8974
rect 1032 8910 1084 8916
rect 1044 7750 1072 8910
rect 1136 7954 1164 8978
rect 1124 7948 1176 7954
rect 1124 7890 1176 7896
rect 1228 7868 1256 9438
rect 1398 9415 1454 9424
rect 1582 9208 1638 9217
rect 1582 9143 1584 9152
rect 1636 9143 1638 9152
rect 1584 9114 1636 9120
rect 1688 8974 1716 9590
rect 1872 9110 1900 12406
rect 1952 12378 2004 12384
rect 1950 12200 2006 12209
rect 2056 12170 2084 12718
rect 1950 12135 2006 12144
rect 2044 12164 2096 12170
rect 1964 11762 1992 12135
rect 2044 12106 2096 12112
rect 2148 12084 2176 13126
rect 2320 12912 2372 12918
rect 2318 12880 2320 12889
rect 2372 12880 2374 12889
rect 2318 12815 2374 12824
rect 2332 12714 2360 12815
rect 2228 12708 2280 12714
rect 2228 12650 2280 12656
rect 2320 12708 2372 12714
rect 2320 12650 2372 12656
rect 2240 12442 2268 12650
rect 2412 12640 2464 12646
rect 2412 12582 2464 12588
rect 2228 12436 2280 12442
rect 2280 12406 2360 12434
rect 2228 12378 2280 12384
rect 2228 12096 2280 12102
rect 2148 12056 2228 12084
rect 2228 12038 2280 12044
rect 1952 11756 2004 11762
rect 1952 11698 2004 11704
rect 1964 11642 1992 11698
rect 1964 11614 2084 11642
rect 1952 11552 2004 11558
rect 1952 11494 2004 11500
rect 1964 10538 1992 11494
rect 1952 10532 2004 10538
rect 1952 10474 2004 10480
rect 1952 10124 2004 10130
rect 1952 10066 2004 10072
rect 1964 9722 1992 10066
rect 1952 9716 2004 9722
rect 1952 9658 2004 9664
rect 2056 9466 2084 11614
rect 2332 11354 2360 12406
rect 2424 12374 2452 12582
rect 2412 12368 2464 12374
rect 2412 12310 2464 12316
rect 2320 11348 2372 11354
rect 2320 11290 2372 11296
rect 2228 10600 2280 10606
rect 2228 10542 2280 10548
rect 2136 9920 2188 9926
rect 2136 9862 2188 9868
rect 1964 9438 2084 9466
rect 1964 9217 1992 9438
rect 2044 9376 2096 9382
rect 2044 9318 2096 9324
rect 1950 9208 2006 9217
rect 1950 9143 2006 9152
rect 1860 9104 1912 9110
rect 1860 9046 1912 9052
rect 1768 9036 1820 9042
rect 1768 8978 1820 8984
rect 1676 8968 1728 8974
rect 1676 8910 1728 8916
rect 1364 8732 1740 8741
rect 1420 8730 1444 8732
rect 1500 8730 1524 8732
rect 1580 8730 1604 8732
rect 1660 8730 1684 8732
rect 1420 8678 1430 8730
rect 1674 8678 1684 8730
rect 1420 8676 1444 8678
rect 1500 8676 1524 8678
rect 1580 8676 1604 8678
rect 1660 8676 1684 8678
rect 1364 8667 1740 8676
rect 1780 8090 1808 8978
rect 2056 8838 2084 9318
rect 2044 8832 2096 8838
rect 2044 8774 2096 8780
rect 1952 8628 2004 8634
rect 1952 8570 2004 8576
rect 1768 8084 1820 8090
rect 1768 8026 1820 8032
rect 1308 7880 1360 7886
rect 1228 7840 1308 7868
rect 1308 7822 1360 7828
rect 848 7744 900 7750
rect 848 7686 900 7692
rect 1032 7744 1084 7750
rect 1032 7686 1084 7692
rect 860 5710 888 7686
rect 848 5704 900 5710
rect 848 5646 900 5652
rect 664 4684 716 4690
rect 664 4626 716 4632
rect 1044 3058 1072 7686
rect 1364 7644 1740 7653
rect 1420 7642 1444 7644
rect 1500 7642 1524 7644
rect 1580 7642 1604 7644
rect 1660 7642 1684 7644
rect 1420 7590 1430 7642
rect 1674 7590 1684 7642
rect 1420 7588 1444 7590
rect 1500 7588 1524 7590
rect 1580 7588 1604 7590
rect 1660 7588 1684 7590
rect 1364 7579 1740 7588
rect 1780 7410 1808 8026
rect 1860 7948 1912 7954
rect 1860 7890 1912 7896
rect 1768 7404 1820 7410
rect 1768 7346 1820 7352
rect 1124 7336 1176 7342
rect 1124 7278 1176 7284
rect 1492 7336 1544 7342
rect 1492 7278 1544 7284
rect 1136 6798 1164 7278
rect 1504 7002 1532 7278
rect 1780 7002 1808 7346
rect 1872 7206 1900 7890
rect 1964 7546 1992 8570
rect 2056 8430 2084 8774
rect 2044 8424 2096 8430
rect 2044 8366 2096 8372
rect 2148 7954 2176 9862
rect 2240 8514 2268 10542
rect 2332 8673 2360 11290
rect 2412 11008 2464 11014
rect 2412 10950 2464 10956
rect 2424 10674 2452 10950
rect 2412 10668 2464 10674
rect 2412 10610 2464 10616
rect 2318 8664 2374 8673
rect 2318 8599 2374 8608
rect 2240 8486 2360 8514
rect 2228 8424 2280 8430
rect 2228 8366 2280 8372
rect 2240 8090 2268 8366
rect 2228 8084 2280 8090
rect 2228 8026 2280 8032
rect 2136 7948 2188 7954
rect 2136 7890 2188 7896
rect 2136 7812 2188 7818
rect 2136 7754 2188 7760
rect 1952 7540 2004 7546
rect 1952 7482 2004 7488
rect 2148 7274 2176 7754
rect 2136 7268 2188 7274
rect 2136 7210 2188 7216
rect 1860 7200 1912 7206
rect 1860 7142 1912 7148
rect 1492 6996 1544 7002
rect 1492 6938 1544 6944
rect 1768 6996 1820 7002
rect 1768 6938 1820 6944
rect 1780 6866 1808 6938
rect 1872 6866 1900 7142
rect 2148 6866 2176 7210
rect 1768 6860 1820 6866
rect 1768 6802 1820 6808
rect 1860 6860 1912 6866
rect 1860 6802 1912 6808
rect 2136 6860 2188 6866
rect 2136 6802 2188 6808
rect 1124 6792 1176 6798
rect 1124 6734 1176 6740
rect 1136 4826 1164 6734
rect 1364 6556 1740 6565
rect 1420 6554 1444 6556
rect 1500 6554 1524 6556
rect 1580 6554 1604 6556
rect 1660 6554 1684 6556
rect 1420 6502 1430 6554
rect 1674 6502 1684 6554
rect 1420 6500 1444 6502
rect 1500 6500 1524 6502
rect 1580 6500 1604 6502
rect 1660 6500 1684 6502
rect 1364 6491 1740 6500
rect 1768 6248 1820 6254
rect 1768 6190 1820 6196
rect 1780 5778 1808 6190
rect 1768 5772 1820 5778
rect 1768 5714 1820 5720
rect 1364 5468 1740 5477
rect 1420 5466 1444 5468
rect 1500 5466 1524 5468
rect 1580 5466 1604 5468
rect 1660 5466 1684 5468
rect 1420 5414 1430 5466
rect 1674 5414 1684 5466
rect 1420 5412 1444 5414
rect 1500 5412 1524 5414
rect 1580 5412 1604 5414
rect 1660 5412 1684 5414
rect 1364 5403 1740 5412
rect 1780 5370 1808 5714
rect 1872 5370 1900 6802
rect 2044 6248 2096 6254
rect 2044 6190 2096 6196
rect 2136 6248 2188 6254
rect 2136 6190 2188 6196
rect 1952 6112 2004 6118
rect 1952 6054 2004 6060
rect 1964 5778 1992 6054
rect 1952 5772 2004 5778
rect 1952 5714 2004 5720
rect 1952 5636 2004 5642
rect 1952 5578 2004 5584
rect 1768 5364 1820 5370
rect 1768 5306 1820 5312
rect 1860 5364 1912 5370
rect 1860 5306 1912 5312
rect 1676 5296 1728 5302
rect 1676 5238 1728 5244
rect 1688 5166 1716 5238
rect 1860 5228 1912 5234
rect 1860 5170 1912 5176
rect 1492 5160 1544 5166
rect 1492 5102 1544 5108
rect 1676 5160 1728 5166
rect 1676 5102 1728 5108
rect 1308 5024 1360 5030
rect 1308 4966 1360 4972
rect 1124 4820 1176 4826
rect 1124 4762 1176 4768
rect 1320 4690 1348 4966
rect 1504 4758 1532 5102
rect 1688 5030 1716 5102
rect 1676 5024 1728 5030
rect 1676 4966 1728 4972
rect 1492 4752 1544 4758
rect 1492 4694 1544 4700
rect 1872 4690 1900 5170
rect 1308 4684 1360 4690
rect 1228 4644 1308 4672
rect 1124 4616 1176 4622
rect 1124 4558 1176 4564
rect 1136 3466 1164 4558
rect 1228 3670 1256 4644
rect 1308 4626 1360 4632
rect 1860 4684 1912 4690
rect 1860 4626 1912 4632
rect 1768 4548 1820 4554
rect 1768 4490 1820 4496
rect 1364 4380 1740 4389
rect 1420 4378 1444 4380
rect 1500 4378 1524 4380
rect 1580 4378 1604 4380
rect 1660 4378 1684 4380
rect 1420 4326 1430 4378
rect 1674 4326 1684 4378
rect 1420 4324 1444 4326
rect 1500 4324 1524 4326
rect 1580 4324 1604 4326
rect 1660 4324 1684 4326
rect 1364 4315 1740 4324
rect 1676 4140 1728 4146
rect 1676 4082 1728 4088
rect 1688 3738 1716 4082
rect 1780 4078 1808 4490
rect 1768 4072 1820 4078
rect 1768 4014 1820 4020
rect 1676 3732 1728 3738
rect 1676 3674 1728 3680
rect 1216 3664 1268 3670
rect 1216 3606 1268 3612
rect 1124 3460 1176 3466
rect 1124 3402 1176 3408
rect 1364 3292 1740 3301
rect 1420 3290 1444 3292
rect 1500 3290 1524 3292
rect 1580 3290 1604 3292
rect 1660 3290 1684 3292
rect 1420 3238 1430 3290
rect 1674 3238 1684 3290
rect 1420 3236 1444 3238
rect 1500 3236 1524 3238
rect 1580 3236 1604 3238
rect 1660 3236 1684 3238
rect 1364 3227 1740 3236
rect 1964 3126 1992 5578
rect 2056 5370 2084 6190
rect 2044 5364 2096 5370
rect 2044 5306 2096 5312
rect 2148 5166 2176 6190
rect 2228 6112 2280 6118
rect 2228 6054 2280 6060
rect 2136 5160 2188 5166
rect 2136 5102 2188 5108
rect 2240 5098 2268 6054
rect 2228 5092 2280 5098
rect 2228 5034 2280 5040
rect 2240 4758 2268 5034
rect 2332 4826 2360 8486
rect 2424 6254 2452 10610
rect 2516 8634 2544 13262
rect 2608 10130 2636 13466
rect 2700 13326 2728 13942
rect 3056 13932 3108 13938
rect 3056 13874 3108 13880
rect 3068 13462 3096 13874
rect 3056 13456 3108 13462
rect 3056 13398 3108 13404
rect 2688 13320 2740 13326
rect 2688 13262 2740 13268
rect 2964 12776 3016 12782
rect 2964 12718 3016 12724
rect 2780 12096 2832 12102
rect 2780 12038 2832 12044
rect 2792 11694 2820 12038
rect 2780 11688 2832 11694
rect 2780 11630 2832 11636
rect 2688 11552 2740 11558
rect 2688 11494 2740 11500
rect 2596 10124 2648 10130
rect 2596 10066 2648 10072
rect 2608 9518 2636 10066
rect 2596 9512 2648 9518
rect 2596 9454 2648 9460
rect 2608 9178 2636 9454
rect 2596 9172 2648 9178
rect 2596 9114 2648 9120
rect 2700 9058 2728 11494
rect 2792 11218 2820 11630
rect 2976 11354 3004 12718
rect 3160 12434 3188 14214
rect 3332 12708 3384 12714
rect 3332 12650 3384 12656
rect 3068 12406 3188 12434
rect 2964 11348 3016 11354
rect 2964 11290 3016 11296
rect 2780 11212 2832 11218
rect 2780 11154 2832 11160
rect 2964 9920 3016 9926
rect 2964 9862 3016 9868
rect 2608 9030 2728 9058
rect 2872 9104 2924 9110
rect 2872 9046 2924 9052
rect 2780 9036 2832 9042
rect 2504 8628 2556 8634
rect 2504 8570 2556 8576
rect 2504 7948 2556 7954
rect 2504 7890 2556 7896
rect 2516 7546 2544 7890
rect 2504 7540 2556 7546
rect 2504 7482 2556 7488
rect 2504 6860 2556 6866
rect 2504 6802 2556 6808
rect 2412 6248 2464 6254
rect 2412 6190 2464 6196
rect 2412 6112 2464 6118
rect 2412 6054 2464 6060
rect 2424 5710 2452 6054
rect 2516 5778 2544 6802
rect 2504 5772 2556 5778
rect 2504 5714 2556 5720
rect 2412 5704 2464 5710
rect 2412 5646 2464 5652
rect 2320 4820 2372 4826
rect 2320 4762 2372 4768
rect 2228 4752 2280 4758
rect 2228 4694 2280 4700
rect 2044 4684 2096 4690
rect 2044 4626 2096 4632
rect 2320 4684 2372 4690
rect 2320 4626 2372 4632
rect 2056 3194 2084 4626
rect 2332 4282 2360 4626
rect 2320 4276 2372 4282
rect 2320 4218 2372 4224
rect 2044 3188 2096 3194
rect 2044 3130 2096 3136
rect 1952 3120 2004 3126
rect 1952 3062 2004 3068
rect 1032 3052 1084 3058
rect 1032 2994 1084 3000
rect 2056 2774 2084 3130
rect 1964 2746 2084 2774
rect 1364 2204 1740 2213
rect 1420 2202 1444 2204
rect 1500 2202 1524 2204
rect 1580 2202 1604 2204
rect 1660 2202 1684 2204
rect 1420 2150 1430 2202
rect 1674 2150 1684 2202
rect 1420 2148 1444 2150
rect 1500 2148 1524 2150
rect 1580 2148 1604 2150
rect 1660 2148 1684 2150
rect 1364 2139 1740 2148
rect 1860 2032 1912 2038
rect 1860 1974 1912 1980
rect 756 1556 808 1562
rect 756 1498 808 1504
rect 572 1488 624 1494
rect 572 1430 624 1436
rect 584 626 612 1430
rect 400 598 612 626
rect 400 400 428 598
rect 768 400 796 1498
rect 1872 1426 1900 1974
rect 1964 1902 1992 2746
rect 2516 1970 2544 5714
rect 2608 4554 2636 9030
rect 2780 8978 2832 8984
rect 2792 8922 2820 8978
rect 2700 8894 2820 8922
rect 2700 7954 2728 8894
rect 2884 8072 2912 9046
rect 2976 9042 3004 9862
rect 3068 9674 3096 12406
rect 3344 11218 3372 12650
rect 3424 12300 3476 12306
rect 3424 12242 3476 12248
rect 3436 11694 3464 12242
rect 3424 11688 3476 11694
rect 3424 11630 3476 11636
rect 3424 11280 3476 11286
rect 3424 11222 3476 11228
rect 3332 11212 3384 11218
rect 3332 11154 3384 11160
rect 3148 11144 3200 11150
rect 3200 11092 3280 11098
rect 3148 11086 3280 11092
rect 3160 11070 3280 11086
rect 3148 11008 3200 11014
rect 3148 10950 3200 10956
rect 3160 10130 3188 10950
rect 3148 10124 3200 10130
rect 3148 10066 3200 10072
rect 3068 9646 3188 9674
rect 3056 9376 3108 9382
rect 3056 9318 3108 9324
rect 3068 9042 3096 9318
rect 2964 9036 3016 9042
rect 2964 8978 3016 8984
rect 3056 9036 3108 9042
rect 3056 8978 3108 8984
rect 3160 8430 3188 9646
rect 3148 8424 3200 8430
rect 3146 8392 3148 8401
rect 3200 8392 3202 8401
rect 3146 8327 3202 8336
rect 2792 8044 2912 8072
rect 2792 7954 2820 8044
rect 3146 7984 3202 7993
rect 2688 7948 2740 7954
rect 2688 7890 2740 7896
rect 2780 7948 2832 7954
rect 2780 7890 2832 7896
rect 2872 7948 2924 7954
rect 3146 7919 3148 7928
rect 2872 7890 2924 7896
rect 3200 7919 3202 7928
rect 3148 7890 3200 7896
rect 2700 6866 2728 7890
rect 2688 6860 2740 6866
rect 2688 6802 2740 6808
rect 2700 4826 2728 6802
rect 2884 6746 2912 7890
rect 2964 7880 3016 7886
rect 2964 7822 3016 7828
rect 2976 7410 3004 7822
rect 3056 7812 3108 7818
rect 3056 7754 3108 7760
rect 2964 7404 3016 7410
rect 2964 7346 3016 7352
rect 2976 6934 3004 7346
rect 2964 6928 3016 6934
rect 2964 6870 3016 6876
rect 3068 6798 3096 7754
rect 3160 7410 3188 7890
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 2792 6730 2912 6746
rect 3056 6792 3108 6798
rect 3056 6734 3108 6740
rect 2780 6724 2912 6730
rect 2832 6718 2912 6724
rect 2780 6666 2832 6672
rect 2872 5704 2924 5710
rect 2872 5646 2924 5652
rect 2884 5166 2912 5646
rect 2872 5160 2924 5166
rect 2872 5102 2924 5108
rect 3252 4826 3280 11070
rect 3344 10674 3372 11154
rect 3332 10668 3384 10674
rect 3332 10610 3384 10616
rect 3436 9926 3464 11222
rect 3424 9920 3476 9926
rect 3424 9862 3476 9868
rect 3424 9580 3476 9586
rect 3424 9522 3476 9528
rect 3330 9480 3386 9489
rect 3330 9415 3386 9424
rect 3344 9382 3372 9415
rect 3332 9376 3384 9382
rect 3332 9318 3384 9324
rect 3332 9172 3384 9178
rect 3332 9114 3384 9120
rect 3344 7954 3372 9114
rect 3436 8022 3464 9522
rect 3528 9042 3556 14282
rect 3608 13864 3660 13870
rect 3608 13806 3660 13812
rect 3620 13394 3648 13806
rect 3608 13388 3660 13394
rect 3660 13348 3740 13376
rect 3608 13330 3660 13336
rect 3608 12640 3660 12646
rect 3608 12582 3660 12588
rect 3620 12306 3648 12582
rect 3712 12442 3740 13348
rect 3700 12436 3752 12442
rect 3700 12378 3752 12384
rect 3804 12322 3832 14758
rect 3896 14521 3924 14826
rect 3882 14512 3938 14521
rect 3882 14447 3884 14456
rect 3936 14447 3938 14456
rect 3884 14418 3936 14424
rect 3988 13954 4016 16730
rect 4080 16658 4108 18119
rect 4172 17882 4200 18226
rect 4252 18148 4304 18154
rect 4252 18090 4304 18096
rect 4160 17876 4212 17882
rect 4160 17818 4212 17824
rect 4068 16652 4120 16658
rect 4068 16594 4120 16600
rect 4172 16538 4200 17818
rect 4264 16658 4292 18090
rect 4804 18080 4856 18086
rect 4804 18022 4856 18028
rect 4896 18080 4948 18086
rect 4896 18022 4948 18028
rect 4988 18080 5040 18086
rect 4988 18022 5040 18028
rect 4364 17980 4740 17989
rect 4420 17978 4444 17980
rect 4500 17978 4524 17980
rect 4580 17978 4604 17980
rect 4660 17978 4684 17980
rect 4420 17926 4430 17978
rect 4674 17926 4684 17978
rect 4420 17924 4444 17926
rect 4500 17924 4524 17926
rect 4580 17924 4604 17926
rect 4660 17924 4684 17926
rect 4364 17915 4740 17924
rect 4816 17746 4844 18022
rect 4804 17740 4856 17746
rect 4804 17682 4856 17688
rect 4908 17354 4936 18022
rect 4816 17326 4936 17354
rect 4364 16892 4740 16901
rect 4420 16890 4444 16892
rect 4500 16890 4524 16892
rect 4580 16890 4604 16892
rect 4660 16890 4684 16892
rect 4420 16838 4430 16890
rect 4674 16838 4684 16890
rect 4420 16836 4444 16838
rect 4500 16836 4524 16838
rect 4580 16836 4604 16838
rect 4660 16836 4684 16838
rect 4364 16827 4740 16836
rect 4344 16788 4396 16794
rect 4344 16730 4396 16736
rect 4528 16788 4580 16794
rect 4528 16730 4580 16736
rect 4252 16652 4304 16658
rect 4252 16594 4304 16600
rect 4356 16538 4384 16730
rect 4172 16510 4384 16538
rect 4172 15026 4200 16510
rect 4540 15892 4568 16730
rect 4816 16561 4844 17326
rect 4802 16552 4858 16561
rect 4802 16487 4804 16496
rect 4856 16487 4858 16496
rect 4804 16458 4856 16464
rect 5000 16250 5028 18022
rect 5092 17241 5120 18255
rect 5172 18226 5224 18232
rect 5264 18284 5316 18290
rect 5264 18226 5316 18232
rect 5078 17232 5134 17241
rect 5078 17167 5134 17176
rect 5080 17128 5132 17134
rect 5080 17070 5132 17076
rect 5092 16794 5120 17070
rect 5080 16788 5132 16794
rect 5080 16730 5132 16736
rect 5184 16658 5212 18226
rect 5276 17814 5304 18226
rect 5460 17882 5488 18634
rect 5448 17876 5500 17882
rect 5448 17818 5500 17824
rect 5264 17808 5316 17814
rect 5264 17750 5316 17756
rect 5356 17672 5408 17678
rect 5356 17614 5408 17620
rect 5262 17096 5318 17105
rect 5262 17031 5318 17040
rect 5276 16794 5304 17031
rect 5264 16788 5316 16794
rect 5264 16730 5316 16736
rect 5172 16652 5224 16658
rect 5172 16594 5224 16600
rect 4988 16244 5040 16250
rect 4988 16186 5040 16192
rect 4896 16108 4948 16114
rect 4896 16050 4948 16056
rect 4804 15972 4856 15978
rect 4804 15914 4856 15920
rect 4264 15864 4568 15892
rect 4264 15314 4292 15864
rect 4364 15804 4740 15813
rect 4420 15802 4444 15804
rect 4500 15802 4524 15804
rect 4580 15802 4604 15804
rect 4660 15802 4684 15804
rect 4420 15750 4430 15802
rect 4674 15750 4684 15802
rect 4420 15748 4444 15750
rect 4500 15748 4524 15750
rect 4580 15748 4604 15750
rect 4660 15748 4684 15750
rect 4364 15739 4740 15748
rect 4264 15286 4384 15314
rect 4250 15192 4306 15201
rect 4250 15127 4306 15136
rect 4160 15020 4212 15026
rect 4160 14962 4212 14968
rect 4068 14952 4120 14958
rect 4068 14894 4120 14900
rect 4080 14618 4108 14894
rect 4264 14618 4292 15127
rect 4356 14958 4384 15286
rect 4712 15156 4764 15162
rect 4816 15144 4844 15914
rect 4764 15116 4844 15144
rect 4712 15098 4764 15104
rect 4434 15056 4490 15065
rect 4908 15026 4936 16050
rect 5000 16046 5028 16186
rect 4988 16040 5040 16046
rect 5040 15988 5120 15994
rect 4988 15982 5120 15988
rect 5000 15966 5120 15982
rect 4988 15904 5040 15910
rect 4988 15846 5040 15852
rect 5000 15473 5028 15846
rect 4986 15464 5042 15473
rect 4986 15399 5042 15408
rect 4434 14991 4490 15000
rect 4896 15020 4948 15026
rect 4344 14952 4396 14958
rect 4344 14894 4396 14900
rect 4448 14890 4476 14991
rect 4896 14962 4948 14968
rect 4804 14952 4856 14958
rect 4710 14920 4766 14929
rect 4436 14884 4488 14890
rect 4804 14894 4856 14900
rect 4710 14855 4712 14864
rect 4436 14826 4488 14832
rect 4764 14855 4766 14864
rect 4712 14826 4764 14832
rect 4364 14716 4740 14725
rect 4420 14714 4444 14716
rect 4500 14714 4524 14716
rect 4580 14714 4604 14716
rect 4660 14714 4684 14716
rect 4420 14662 4430 14714
rect 4674 14662 4684 14714
rect 4420 14660 4444 14662
rect 4500 14660 4524 14662
rect 4580 14660 4604 14662
rect 4660 14660 4684 14662
rect 4364 14651 4740 14660
rect 4816 14634 4844 14894
rect 4908 14890 4936 14962
rect 4896 14884 4948 14890
rect 4896 14826 4948 14832
rect 4816 14618 4936 14634
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 4252 14612 4304 14618
rect 4816 14612 4948 14618
rect 4816 14606 4896 14612
rect 4252 14554 4304 14560
rect 4896 14554 4948 14560
rect 4080 14074 4108 14554
rect 4804 14544 4856 14550
rect 4804 14486 4856 14492
rect 4528 14476 4580 14482
rect 4528 14418 4580 14424
rect 4620 14476 4672 14482
rect 4620 14418 4672 14424
rect 4068 14068 4120 14074
rect 4068 14010 4120 14016
rect 4540 14006 4568 14418
rect 4632 14385 4660 14418
rect 4618 14376 4674 14385
rect 4618 14311 4674 14320
rect 4528 14000 4580 14006
rect 3988 13926 4108 13954
rect 4528 13942 4580 13948
rect 3976 13864 4028 13870
rect 3976 13806 4028 13812
rect 3884 13728 3936 13734
rect 3884 13670 3936 13676
rect 3896 12782 3924 13670
rect 3988 13190 4016 13806
rect 3976 13184 4028 13190
rect 3976 13126 4028 13132
rect 3884 12776 3936 12782
rect 3884 12718 3936 12724
rect 3976 12708 4028 12714
rect 3976 12650 4028 12656
rect 3608 12300 3660 12306
rect 3608 12242 3660 12248
rect 3712 12294 3832 12322
rect 3884 12300 3936 12306
rect 3620 11626 3648 12242
rect 3712 11642 3740 12294
rect 3884 12242 3936 12248
rect 3792 12096 3844 12102
rect 3792 12038 3844 12044
rect 3804 11762 3832 12038
rect 3792 11756 3844 11762
rect 3792 11698 3844 11704
rect 3608 11620 3660 11626
rect 3712 11614 3832 11642
rect 3608 11562 3660 11568
rect 3700 11348 3752 11354
rect 3700 11290 3752 11296
rect 3712 11218 3740 11290
rect 3700 11212 3752 11218
rect 3700 11154 3752 11160
rect 3608 10600 3660 10606
rect 3608 10542 3660 10548
rect 3620 10266 3648 10542
rect 3608 10260 3660 10266
rect 3608 10202 3660 10208
rect 3608 9988 3660 9994
rect 3608 9930 3660 9936
rect 3620 9518 3648 9930
rect 3608 9512 3660 9518
rect 3606 9480 3608 9489
rect 3660 9480 3662 9489
rect 3606 9415 3662 9424
rect 3516 9036 3568 9042
rect 3516 8978 3568 8984
rect 3516 8832 3568 8838
rect 3516 8774 3568 8780
rect 3528 8634 3556 8774
rect 3516 8628 3568 8634
rect 3516 8570 3568 8576
rect 3528 8430 3556 8570
rect 3516 8424 3568 8430
rect 3516 8366 3568 8372
rect 3516 8288 3568 8294
rect 3516 8230 3568 8236
rect 3424 8016 3476 8022
rect 3424 7958 3476 7964
rect 3332 7948 3384 7954
rect 3332 7890 3384 7896
rect 3424 7744 3476 7750
rect 3424 7686 3476 7692
rect 3332 7472 3384 7478
rect 3332 7414 3384 7420
rect 3344 5302 3372 7414
rect 3436 7410 3464 7686
rect 3424 7404 3476 7410
rect 3424 7346 3476 7352
rect 3332 5296 3384 5302
rect 3332 5238 3384 5244
rect 2688 4820 2740 4826
rect 2688 4762 2740 4768
rect 2780 4820 2832 4826
rect 2780 4762 2832 4768
rect 3240 4820 3292 4826
rect 3240 4762 3292 4768
rect 2596 4548 2648 4554
rect 2596 4490 2648 4496
rect 2792 4078 2820 4762
rect 2964 4684 3016 4690
rect 2964 4626 3016 4632
rect 2976 4486 3004 4626
rect 2964 4480 3016 4486
rect 2964 4422 3016 4428
rect 2780 4072 2832 4078
rect 2780 4014 2832 4020
rect 2976 4010 3004 4422
rect 3056 4208 3108 4214
rect 3056 4150 3108 4156
rect 2964 4004 3016 4010
rect 2964 3946 3016 3952
rect 3068 3534 3096 4150
rect 3436 4078 3464 7346
rect 3528 6984 3556 8230
rect 3608 7948 3660 7954
rect 3608 7890 3660 7896
rect 3620 7410 3648 7890
rect 3608 7404 3660 7410
rect 3608 7346 3660 7352
rect 3528 6956 3648 6984
rect 3516 6860 3568 6866
rect 3516 6802 3568 6808
rect 3528 6254 3556 6802
rect 3516 6248 3568 6254
rect 3516 6190 3568 6196
rect 3528 5030 3556 6190
rect 3620 5681 3648 6956
rect 3712 6866 3740 11154
rect 3804 9178 3832 11614
rect 3792 9172 3844 9178
rect 3792 9114 3844 9120
rect 3804 8974 3832 9114
rect 3792 8968 3844 8974
rect 3792 8910 3844 8916
rect 3790 8392 3846 8401
rect 3790 8327 3846 8336
rect 3804 8294 3832 8327
rect 3792 8288 3844 8294
rect 3792 8230 3844 8236
rect 3896 7800 3924 12242
rect 3988 12102 4016 12650
rect 4080 12434 4108 13926
rect 4364 13628 4740 13637
rect 4420 13626 4444 13628
rect 4500 13626 4524 13628
rect 4580 13626 4604 13628
rect 4660 13626 4684 13628
rect 4420 13574 4430 13626
rect 4674 13574 4684 13626
rect 4420 13572 4444 13574
rect 4500 13572 4524 13574
rect 4580 13572 4604 13574
rect 4660 13572 4684 13574
rect 4364 13563 4740 13572
rect 4620 13456 4672 13462
rect 4250 13424 4306 13433
rect 4620 13398 4672 13404
rect 4250 13359 4252 13368
rect 4304 13359 4306 13368
rect 4252 13330 4304 13336
rect 4160 13320 4212 13326
rect 4160 13262 4212 13268
rect 4172 12782 4200 13262
rect 4160 12776 4212 12782
rect 4160 12718 4212 12724
rect 4264 12714 4292 13330
rect 4632 12782 4660 13398
rect 4620 12776 4672 12782
rect 4620 12718 4672 12724
rect 4252 12708 4304 12714
rect 4252 12650 4304 12656
rect 4816 12696 4844 14486
rect 5092 14006 5120 15966
rect 5264 15904 5316 15910
rect 5368 15881 5396 17614
rect 5552 17202 5580 19450
rect 5816 19236 5868 19242
rect 5816 19178 5868 19184
rect 5828 18834 5856 19178
rect 6196 18970 6224 19858
rect 6472 19334 6500 20946
rect 6564 20777 6592 21830
rect 6828 21684 6880 21690
rect 6828 21626 6880 21632
rect 6644 21616 6696 21622
rect 6696 21564 6776 21570
rect 6644 21558 6776 21564
rect 6656 21542 6776 21558
rect 6644 21480 6696 21486
rect 6644 21422 6696 21428
rect 6550 20768 6606 20777
rect 6550 20703 6606 20712
rect 6656 20602 6684 21422
rect 6644 20596 6696 20602
rect 6644 20538 6696 20544
rect 6550 20088 6606 20097
rect 6550 20023 6606 20032
rect 6380 19306 6500 19334
rect 6380 19242 6408 19306
rect 6368 19236 6420 19242
rect 6368 19178 6420 19184
rect 6184 18964 6236 18970
rect 6184 18906 6236 18912
rect 5632 18828 5684 18834
rect 5632 18770 5684 18776
rect 5816 18828 5868 18834
rect 5816 18770 5868 18776
rect 5644 17762 5672 18770
rect 6460 18760 6512 18766
rect 6104 18686 6316 18714
rect 6460 18702 6512 18708
rect 6104 18630 6132 18686
rect 5724 18624 5776 18630
rect 5722 18592 5724 18601
rect 6092 18624 6144 18630
rect 5776 18592 5778 18601
rect 6092 18566 6144 18572
rect 6184 18624 6236 18630
rect 6184 18566 6236 18572
rect 5722 18527 5778 18536
rect 5828 18414 6040 18442
rect 5828 18358 5856 18414
rect 5816 18352 5868 18358
rect 5816 18294 5868 18300
rect 5908 18352 5960 18358
rect 5908 18294 5960 18300
rect 5724 18080 5776 18086
rect 5724 18022 5776 18028
rect 5816 18080 5868 18086
rect 5816 18022 5868 18028
rect 5736 17882 5764 18022
rect 5724 17876 5776 17882
rect 5724 17818 5776 17824
rect 5644 17734 5764 17762
rect 5632 17264 5684 17270
rect 5632 17206 5684 17212
rect 5540 17196 5592 17202
rect 5540 17138 5592 17144
rect 5448 17060 5500 17066
rect 5448 17002 5500 17008
rect 5460 16250 5488 17002
rect 5448 16244 5500 16250
rect 5448 16186 5500 16192
rect 5448 15904 5500 15910
rect 5264 15846 5316 15852
rect 5354 15872 5410 15881
rect 5276 14929 5304 15846
rect 5448 15846 5500 15852
rect 5354 15807 5410 15816
rect 5460 15706 5488 15846
rect 5448 15700 5500 15706
rect 5448 15642 5500 15648
rect 5552 15638 5580 17138
rect 5644 16658 5672 17206
rect 5632 16652 5684 16658
rect 5632 16594 5684 16600
rect 5644 16182 5672 16594
rect 5632 16176 5684 16182
rect 5632 16118 5684 16124
rect 5736 16114 5764 17734
rect 5828 17649 5856 18022
rect 5814 17640 5870 17649
rect 5814 17575 5870 17584
rect 5816 17128 5868 17134
rect 5814 17096 5816 17105
rect 5868 17096 5870 17105
rect 5814 17031 5870 17040
rect 5920 16658 5948 18294
rect 5908 16652 5960 16658
rect 5908 16594 5960 16600
rect 5724 16108 5776 16114
rect 5724 16050 5776 16056
rect 5736 15910 5764 16050
rect 5724 15904 5776 15910
rect 5724 15846 5776 15852
rect 6012 15745 6040 18414
rect 6196 18222 6224 18566
rect 6092 18216 6144 18222
rect 6092 18158 6144 18164
rect 6184 18216 6236 18222
rect 6184 18158 6236 18164
rect 6104 17746 6132 18158
rect 6288 18086 6316 18686
rect 6472 18426 6500 18702
rect 6460 18420 6512 18426
rect 6460 18362 6512 18368
rect 6564 18306 6592 20023
rect 6748 19718 6776 21542
rect 6840 20806 6868 21626
rect 6920 21480 6972 21486
rect 6920 21422 6972 21428
rect 7012 21480 7064 21486
rect 7012 21422 7064 21428
rect 6932 21146 6960 21422
rect 6920 21140 6972 21146
rect 7024 21128 7052 21422
rect 7116 21321 7144 21830
rect 7208 21486 7236 22034
rect 7196 21480 7248 21486
rect 7196 21422 7248 21428
rect 7102 21312 7158 21321
rect 7102 21247 7158 21256
rect 7024 21100 7144 21128
rect 6920 21082 6972 21088
rect 6828 20800 6880 20806
rect 6828 20742 6880 20748
rect 6932 20534 6960 21082
rect 7116 21010 7144 21100
rect 7104 21004 7156 21010
rect 7104 20946 7156 20952
rect 7012 20936 7064 20942
rect 7012 20878 7064 20884
rect 6920 20528 6972 20534
rect 6920 20470 6972 20476
rect 6920 20392 6972 20398
rect 6920 20334 6972 20340
rect 6932 20233 6960 20334
rect 7024 20262 7052 20878
rect 7104 20800 7156 20806
rect 7104 20742 7156 20748
rect 7012 20256 7064 20262
rect 6918 20224 6974 20233
rect 7012 20198 7064 20204
rect 6918 20159 6974 20168
rect 6736 19712 6788 19718
rect 6736 19654 6788 19660
rect 6828 19304 6880 19310
rect 6828 19246 6880 19252
rect 6918 19272 6974 19281
rect 6840 19145 6868 19246
rect 6918 19207 6920 19216
rect 6972 19207 6974 19216
rect 6920 19178 6972 19184
rect 6826 19136 6882 19145
rect 6826 19071 6882 19080
rect 7024 18601 7052 20198
rect 7116 19718 7144 20742
rect 7208 20602 7236 21422
rect 7300 20942 7328 22510
rect 7748 22500 7800 22506
rect 7748 22442 7800 22448
rect 7760 22166 7788 22442
rect 7748 22160 7800 22166
rect 7748 22102 7800 22108
rect 7364 21788 7740 21797
rect 7420 21786 7444 21788
rect 7500 21786 7524 21788
rect 7580 21786 7604 21788
rect 7660 21786 7684 21788
rect 7420 21734 7430 21786
rect 7674 21734 7684 21786
rect 7420 21732 7444 21734
rect 7500 21732 7524 21734
rect 7580 21732 7604 21734
rect 7660 21732 7684 21734
rect 7364 21723 7740 21732
rect 7472 21684 7524 21690
rect 7472 21626 7524 21632
rect 7380 21480 7432 21486
rect 7380 21422 7432 21428
rect 7392 21049 7420 21422
rect 7484 21350 7512 21626
rect 7656 21480 7708 21486
rect 7656 21422 7708 21428
rect 7472 21344 7524 21350
rect 7472 21286 7524 21292
rect 7378 21040 7434 21049
rect 7378 20975 7434 20984
rect 7288 20936 7340 20942
rect 7288 20878 7340 20884
rect 7668 20806 7696 21422
rect 7852 21146 7880 22578
rect 8220 22094 8248 23122
rect 8576 22976 8628 22982
rect 8576 22918 8628 22924
rect 8588 22710 8616 22918
rect 8576 22704 8628 22710
rect 8576 22646 8628 22652
rect 8404 22222 8524 22250
rect 8404 22098 8432 22222
rect 8496 22166 8524 22222
rect 8668 22228 8720 22234
rect 8668 22170 8720 22176
rect 8484 22160 8536 22166
rect 8484 22102 8536 22108
rect 8220 22066 8340 22094
rect 8116 22024 8168 22030
rect 8022 21992 8078 22001
rect 7932 21956 7984 21962
rect 8116 21966 8168 21972
rect 8022 21927 8024 21936
rect 7932 21898 7984 21904
rect 8076 21927 8078 21936
rect 8024 21898 8076 21904
rect 7944 21554 7972 21898
rect 8036 21622 8064 21898
rect 8024 21616 8076 21622
rect 8024 21558 8076 21564
rect 7932 21548 7984 21554
rect 7932 21490 7984 21496
rect 7840 21140 7892 21146
rect 7840 21082 7892 21088
rect 7944 21010 7972 21490
rect 8128 21010 8156 21966
rect 8312 21468 8340 22066
rect 8392 22092 8444 22098
rect 8392 22034 8444 22040
rect 8576 21956 8628 21962
rect 8576 21898 8628 21904
rect 8392 21888 8444 21894
rect 8392 21830 8444 21836
rect 8404 21486 8432 21830
rect 8588 21593 8616 21898
rect 8574 21584 8630 21593
rect 8574 21519 8630 21528
rect 8680 21570 8708 22170
rect 8864 21690 8892 23600
rect 9404 23248 9456 23254
rect 9404 23190 9456 23196
rect 9220 23180 9272 23186
rect 9220 23122 9272 23128
rect 9232 22778 9260 23122
rect 9220 22772 9272 22778
rect 9220 22714 9272 22720
rect 9220 22568 9272 22574
rect 9220 22510 9272 22516
rect 9312 22568 9364 22574
rect 9312 22510 9364 22516
rect 9128 22160 9180 22166
rect 9128 22102 9180 22108
rect 9036 21888 9088 21894
rect 9036 21830 9088 21836
rect 8852 21684 8904 21690
rect 8852 21626 8904 21632
rect 8680 21554 8892 21570
rect 8680 21548 8904 21554
rect 8680 21542 8852 21548
rect 8220 21440 8340 21468
rect 8392 21480 8444 21486
rect 7840 21004 7892 21010
rect 7840 20946 7892 20952
rect 7932 21004 7984 21010
rect 7932 20946 7984 20952
rect 8116 21004 8168 21010
rect 8116 20946 8168 20952
rect 7656 20800 7708 20806
rect 7656 20742 7708 20748
rect 7364 20700 7740 20709
rect 7420 20698 7444 20700
rect 7500 20698 7524 20700
rect 7580 20698 7604 20700
rect 7660 20698 7684 20700
rect 7420 20646 7430 20698
rect 7674 20646 7684 20698
rect 7420 20644 7444 20646
rect 7500 20644 7524 20646
rect 7580 20644 7604 20646
rect 7660 20644 7684 20646
rect 7364 20635 7740 20644
rect 7196 20596 7248 20602
rect 7852 20584 7880 20946
rect 7196 20538 7248 20544
rect 7760 20556 7880 20584
rect 7932 20596 7984 20602
rect 7380 20392 7432 20398
rect 7380 20334 7432 20340
rect 7288 19916 7340 19922
rect 7288 19858 7340 19864
rect 7104 19712 7156 19718
rect 7104 19654 7156 19660
rect 7196 19712 7248 19718
rect 7196 19654 7248 19660
rect 7208 19242 7236 19654
rect 7196 19236 7248 19242
rect 7196 19178 7248 19184
rect 7300 18970 7328 19858
rect 7392 19825 7420 20334
rect 7656 20256 7708 20262
rect 7656 20198 7708 20204
rect 7668 19922 7696 20198
rect 7656 19916 7708 19922
rect 7656 19858 7708 19864
rect 7378 19816 7434 19825
rect 7760 19786 7788 20556
rect 7932 20538 7984 20544
rect 7944 20058 7972 20538
rect 8024 20392 8076 20398
rect 8024 20334 8076 20340
rect 7932 20052 7984 20058
rect 7932 19994 7984 20000
rect 8036 19961 8064 20334
rect 8116 20324 8168 20330
rect 8116 20266 8168 20272
rect 8022 19952 8078 19961
rect 7932 19916 7984 19922
rect 8022 19887 8078 19896
rect 7932 19858 7984 19864
rect 7944 19825 7972 19858
rect 7930 19816 7986 19825
rect 7378 19751 7434 19760
rect 7748 19780 7800 19786
rect 7930 19751 7986 19760
rect 7748 19722 7800 19728
rect 8128 19700 8156 20266
rect 8220 20097 8248 21440
rect 8392 21422 8444 21428
rect 8300 21344 8352 21350
rect 8300 21286 8352 21292
rect 8206 20088 8262 20097
rect 8206 20023 8262 20032
rect 8208 19916 8260 19922
rect 8208 19858 8260 19864
rect 7852 19672 8156 19700
rect 7364 19612 7740 19621
rect 7420 19610 7444 19612
rect 7500 19610 7524 19612
rect 7580 19610 7604 19612
rect 7660 19610 7684 19612
rect 7420 19558 7430 19610
rect 7674 19558 7684 19610
rect 7420 19556 7444 19558
rect 7500 19556 7524 19558
rect 7580 19556 7604 19558
rect 7660 19556 7684 19558
rect 7364 19547 7740 19556
rect 7288 18964 7340 18970
rect 7288 18906 7340 18912
rect 7852 18902 7880 19672
rect 8220 19378 8248 19858
rect 7932 19372 7984 19378
rect 7932 19314 7984 19320
rect 8208 19372 8260 19378
rect 8208 19314 8260 19320
rect 7840 18896 7892 18902
rect 7840 18838 7892 18844
rect 7196 18760 7248 18766
rect 7196 18702 7248 18708
rect 7010 18592 7066 18601
rect 7010 18527 7066 18536
rect 6472 18278 6592 18306
rect 7024 18306 7052 18527
rect 7208 18408 7236 18702
rect 7364 18524 7740 18533
rect 7420 18522 7444 18524
rect 7500 18522 7524 18524
rect 7580 18522 7604 18524
rect 7660 18522 7684 18524
rect 7420 18470 7430 18522
rect 7674 18470 7684 18522
rect 7420 18468 7444 18470
rect 7500 18468 7524 18470
rect 7580 18468 7604 18470
rect 7660 18468 7684 18470
rect 7364 18459 7740 18468
rect 7288 18420 7340 18426
rect 7208 18380 7288 18408
rect 7288 18362 7340 18368
rect 7944 18306 7972 19314
rect 8208 19168 8260 19174
rect 8312 19156 8340 21286
rect 8680 20942 8708 21542
rect 8852 21490 8904 21496
rect 8944 21480 8996 21486
rect 8944 21422 8996 21428
rect 8758 21312 8814 21321
rect 8758 21247 8814 21256
rect 8668 20936 8720 20942
rect 8668 20878 8720 20884
rect 8392 20868 8444 20874
rect 8392 20810 8444 20816
rect 8404 20398 8432 20810
rect 8772 20777 8800 21247
rect 8956 21185 8984 21422
rect 8942 21176 8998 21185
rect 8942 21111 8998 21120
rect 8956 20890 8984 21111
rect 9048 21049 9076 21830
rect 9140 21468 9168 22102
rect 9232 21962 9260 22510
rect 9220 21956 9272 21962
rect 9220 21898 9272 21904
rect 9324 21622 9352 22510
rect 9416 22166 9444 23190
rect 9508 22778 9536 23718
rect 9954 23600 10010 24000
rect 10506 23746 10562 24000
rect 10244 23718 10562 23746
rect 9968 22778 9996 23600
rect 10244 23322 10272 23718
rect 10506 23600 10562 23718
rect 11058 23600 11114 24000
rect 11610 23600 11666 24000
rect 12162 23746 12218 24000
rect 11808 23718 12218 23746
rect 10364 23420 10740 23429
rect 10420 23418 10444 23420
rect 10500 23418 10524 23420
rect 10580 23418 10604 23420
rect 10660 23418 10684 23420
rect 10420 23366 10430 23418
rect 10674 23366 10684 23418
rect 10420 23364 10444 23366
rect 10500 23364 10524 23366
rect 10580 23364 10604 23366
rect 10660 23364 10684 23366
rect 10364 23355 10740 23364
rect 11072 23322 11100 23600
rect 11624 23322 11652 23600
rect 11808 23322 11836 23718
rect 12162 23600 12218 23718
rect 12714 23600 12770 24000
rect 13266 23600 13322 24000
rect 17960 23724 18012 23730
rect 17960 23666 18012 23672
rect 17224 23656 17276 23662
rect 10232 23316 10284 23322
rect 10232 23258 10284 23264
rect 11060 23316 11112 23322
rect 11060 23258 11112 23264
rect 11612 23316 11664 23322
rect 11612 23258 11664 23264
rect 11796 23316 11848 23322
rect 11796 23258 11848 23264
rect 10048 23180 10100 23186
rect 10048 23122 10100 23128
rect 10784 23180 10836 23186
rect 10784 23122 10836 23128
rect 10968 23180 11020 23186
rect 10968 23122 11020 23128
rect 11244 23180 11296 23186
rect 11244 23122 11296 23128
rect 11336 23180 11388 23186
rect 11336 23122 11388 23128
rect 11796 23180 11848 23186
rect 11796 23122 11848 23128
rect 9496 22772 9548 22778
rect 9496 22714 9548 22720
rect 9956 22772 10008 22778
rect 9956 22714 10008 22720
rect 9680 22568 9732 22574
rect 10060 22545 10088 23122
rect 10140 23044 10192 23050
rect 10140 22986 10192 22992
rect 10152 22574 10180 22986
rect 10796 22681 10824 23122
rect 10782 22672 10838 22681
rect 10782 22607 10838 22616
rect 10140 22568 10192 22574
rect 9680 22510 9732 22516
rect 10046 22536 10102 22545
rect 9692 22409 9720 22510
rect 10140 22510 10192 22516
rect 10046 22471 10102 22480
rect 9678 22400 9734 22409
rect 9678 22335 9734 22344
rect 9680 22228 9732 22234
rect 9680 22170 9732 22176
rect 9404 22160 9456 22166
rect 9404 22102 9456 22108
rect 9692 22094 9720 22170
rect 10048 22160 10100 22166
rect 10048 22102 10100 22108
rect 9600 22066 9720 22094
rect 9600 22030 9628 22066
rect 9496 22024 9548 22030
rect 9402 21992 9458 22001
rect 9496 21966 9548 21972
rect 9588 22024 9640 22030
rect 9588 21966 9640 21972
rect 9680 22024 9732 22030
rect 9680 21966 9732 21972
rect 9402 21927 9458 21936
rect 9416 21894 9444 21927
rect 9404 21888 9456 21894
rect 9404 21830 9456 21836
rect 9508 21622 9536 21966
rect 9312 21616 9364 21622
rect 9312 21558 9364 21564
rect 9496 21616 9548 21622
rect 9496 21558 9548 21564
rect 9312 21480 9364 21486
rect 9140 21440 9312 21468
rect 9312 21422 9364 21428
rect 9034 21040 9090 21049
rect 9034 20975 9090 20984
rect 8956 20862 9168 20890
rect 8758 20768 8814 20777
rect 8758 20703 8814 20712
rect 8576 20596 8628 20602
rect 8576 20538 8628 20544
rect 8588 20398 8616 20538
rect 8772 20398 8800 20703
rect 8392 20392 8444 20398
rect 8392 20334 8444 20340
rect 8576 20392 8628 20398
rect 8576 20334 8628 20340
rect 8760 20392 8812 20398
rect 8760 20334 8812 20340
rect 8484 20256 8536 20262
rect 8588 20233 8616 20334
rect 8484 20198 8536 20204
rect 8574 20224 8630 20233
rect 8496 19854 8524 20198
rect 8574 20159 8630 20168
rect 8852 19984 8904 19990
rect 8680 19944 8852 19972
rect 8484 19848 8536 19854
rect 8536 19796 8616 19802
rect 8484 19790 8616 19796
rect 8496 19774 8616 19790
rect 8484 19712 8536 19718
rect 8484 19654 8536 19660
rect 8260 19128 8340 19156
rect 8208 19110 8260 19116
rect 8312 18834 8340 19128
rect 8496 18902 8524 19654
rect 8484 18896 8536 18902
rect 8484 18838 8536 18844
rect 8588 18834 8616 19774
rect 8680 19514 8708 19944
rect 8852 19926 8904 19932
rect 8852 19848 8904 19854
rect 8852 19790 8904 19796
rect 8864 19514 8892 19790
rect 9036 19780 9088 19786
rect 9036 19722 9088 19728
rect 8944 19712 8996 19718
rect 8944 19654 8996 19660
rect 8668 19508 8720 19514
rect 8668 19450 8720 19456
rect 8852 19508 8904 19514
rect 8852 19450 8904 19456
rect 8666 19272 8722 19281
rect 8666 19207 8668 19216
rect 8720 19207 8722 19216
rect 8668 19178 8720 19184
rect 8760 19168 8812 19174
rect 8760 19110 8812 19116
rect 8668 18896 8720 18902
rect 8668 18838 8720 18844
rect 8300 18828 8352 18834
rect 8300 18770 8352 18776
rect 8576 18828 8628 18834
rect 8576 18770 8628 18776
rect 8024 18692 8076 18698
rect 8024 18634 8076 18640
rect 7024 18278 7604 18306
rect 6368 18148 6420 18154
rect 6368 18090 6420 18096
rect 6276 18080 6328 18086
rect 6276 18022 6328 18028
rect 6380 17882 6408 18090
rect 6184 17876 6236 17882
rect 6184 17818 6236 17824
rect 6368 17876 6420 17882
rect 6368 17818 6420 17824
rect 6092 17740 6144 17746
rect 6092 17682 6144 17688
rect 6092 17536 6144 17542
rect 6092 17478 6144 17484
rect 6104 16998 6132 17478
rect 6196 17338 6224 17818
rect 6472 17762 6500 18278
rect 6920 18216 6972 18222
rect 7196 18216 7248 18222
rect 6972 18164 7144 18170
rect 6920 18158 7144 18164
rect 7196 18158 7248 18164
rect 7380 18216 7432 18222
rect 7380 18158 7432 18164
rect 7472 18216 7524 18222
rect 7472 18158 7524 18164
rect 6828 18148 6880 18154
rect 6932 18142 7144 18158
rect 6828 18090 6880 18096
rect 6642 17912 6698 17921
rect 6552 17876 6604 17882
rect 6642 17847 6698 17856
rect 6552 17818 6604 17824
rect 6288 17734 6500 17762
rect 6184 17332 6236 17338
rect 6184 17274 6236 17280
rect 6288 17066 6316 17734
rect 6368 17672 6420 17678
rect 6366 17640 6368 17649
rect 6564 17660 6592 17818
rect 6420 17640 6422 17649
rect 6366 17575 6422 17584
rect 6472 17632 6592 17660
rect 6368 17332 6420 17338
rect 6368 17274 6420 17280
rect 6380 17134 6408 17274
rect 6368 17128 6420 17134
rect 6368 17070 6420 17076
rect 6276 17060 6328 17066
rect 6276 17002 6328 17008
rect 6092 16992 6144 16998
rect 6092 16934 6144 16940
rect 6274 16960 6330 16969
rect 6274 16895 6330 16904
rect 6184 16040 6236 16046
rect 6184 15982 6236 15988
rect 5998 15736 6054 15745
rect 5998 15671 6054 15680
rect 5540 15632 5592 15638
rect 5446 15600 5502 15609
rect 5540 15574 5592 15580
rect 5446 15535 5502 15544
rect 5460 15502 5488 15535
rect 5448 15496 5500 15502
rect 5448 15438 5500 15444
rect 5262 14920 5318 14929
rect 5172 14884 5224 14890
rect 5262 14855 5318 14864
rect 5172 14826 5224 14832
rect 5184 14482 5212 14826
rect 5276 14521 5304 14855
rect 5460 14634 5488 15438
rect 6196 14958 6224 15982
rect 6288 15502 6316 16895
rect 6380 16697 6408 17070
rect 6366 16688 6422 16697
rect 6366 16623 6422 16632
rect 6472 16454 6500 17632
rect 6656 16794 6684 17847
rect 6840 17814 6868 18090
rect 6920 18080 6972 18086
rect 6920 18022 6972 18028
rect 6828 17808 6880 17814
rect 6828 17750 6880 17756
rect 6932 17649 6960 18022
rect 7116 17762 7144 18142
rect 7208 18086 7236 18158
rect 7196 18080 7248 18086
rect 7196 18022 7248 18028
rect 7392 17921 7420 18158
rect 7378 17912 7434 17921
rect 7378 17847 7434 17856
rect 7380 17808 7432 17814
rect 7116 17756 7380 17762
rect 7116 17750 7432 17756
rect 7116 17734 7420 17750
rect 6918 17640 6974 17649
rect 6736 17604 6788 17610
rect 7484 17626 7512 18158
rect 7576 17678 7604 18278
rect 7852 18278 7972 18306
rect 7656 18216 7708 18222
rect 7656 18158 7708 18164
rect 7668 18057 7696 18158
rect 7654 18048 7710 18057
rect 7654 17983 7710 17992
rect 7852 17882 7880 18278
rect 8036 18222 8064 18634
rect 8576 18624 8628 18630
rect 8680 18612 8708 18838
rect 8628 18584 8708 18612
rect 8576 18566 8628 18572
rect 8392 18352 8444 18358
rect 8392 18294 8444 18300
rect 7932 18216 7984 18222
rect 7932 18158 7984 18164
rect 8024 18216 8076 18222
rect 8024 18158 8076 18164
rect 7944 17882 7972 18158
rect 8024 18080 8076 18086
rect 8024 18022 8076 18028
rect 7840 17876 7892 17882
rect 7840 17818 7892 17824
rect 7932 17876 7984 17882
rect 7932 17818 7984 17824
rect 8036 17814 8064 18022
rect 8024 17808 8076 17814
rect 8024 17750 8076 17756
rect 8208 17808 8260 17814
rect 8208 17750 8260 17756
rect 8036 17678 8064 17750
rect 6918 17575 6974 17584
rect 7116 17598 7512 17626
rect 7564 17672 7616 17678
rect 7564 17614 7616 17620
rect 7932 17672 7984 17678
rect 7932 17614 7984 17620
rect 8024 17672 8076 17678
rect 8024 17614 8076 17620
rect 7840 17604 7892 17610
rect 6736 17546 6788 17552
rect 6748 16998 6776 17546
rect 7116 17338 7144 17598
rect 7840 17546 7892 17552
rect 7196 17536 7248 17542
rect 7196 17478 7248 17484
rect 7288 17536 7340 17542
rect 7288 17478 7340 17484
rect 7208 17338 7236 17478
rect 7104 17332 7156 17338
rect 7104 17274 7156 17280
rect 7196 17332 7248 17338
rect 7196 17274 7248 17280
rect 6828 17264 6880 17270
rect 6828 17206 6880 17212
rect 6736 16992 6788 16998
rect 6736 16934 6788 16940
rect 6644 16788 6696 16794
rect 6644 16730 6696 16736
rect 6460 16448 6512 16454
rect 6460 16390 6512 16396
rect 6552 16448 6604 16454
rect 6552 16390 6604 16396
rect 6564 16046 6592 16390
rect 6840 16182 6868 17206
rect 7010 17096 7066 17105
rect 7066 17040 7144 17048
rect 7010 17031 7012 17040
rect 7064 17020 7144 17040
rect 7012 17002 7064 17008
rect 7012 16652 7064 16658
rect 7012 16594 7064 16600
rect 6828 16176 6880 16182
rect 6734 16144 6790 16153
rect 6828 16118 6880 16124
rect 6734 16079 6736 16088
rect 6788 16079 6790 16088
rect 6736 16050 6788 16056
rect 6552 16040 6604 16046
rect 6552 15982 6604 15988
rect 6460 15972 6512 15978
rect 6460 15914 6512 15920
rect 6276 15496 6328 15502
rect 6276 15438 6328 15444
rect 5540 14952 5592 14958
rect 5540 14894 5592 14900
rect 6184 14952 6236 14958
rect 6184 14894 6236 14900
rect 5368 14606 5488 14634
rect 5262 14512 5318 14521
rect 5172 14476 5224 14482
rect 5262 14447 5318 14456
rect 5172 14418 5224 14424
rect 5080 14000 5132 14006
rect 5080 13942 5132 13948
rect 5080 13864 5132 13870
rect 5080 13806 5132 13812
rect 4988 13388 5040 13394
rect 4988 13330 5040 13336
rect 5000 12782 5028 13330
rect 5092 12986 5120 13806
rect 5080 12980 5132 12986
rect 5080 12922 5132 12928
rect 4988 12776 5040 12782
rect 4988 12718 5040 12724
rect 4896 12708 4948 12714
rect 4816 12668 4896 12696
rect 4160 12640 4212 12646
rect 4212 12588 4292 12594
rect 4160 12582 4292 12588
rect 4172 12566 4292 12582
rect 4080 12406 4200 12434
rect 4068 12368 4120 12374
rect 4068 12310 4120 12316
rect 4080 12102 4108 12310
rect 4172 12306 4200 12406
rect 4160 12300 4212 12306
rect 4160 12242 4212 12248
rect 4264 12170 4292 12566
rect 4364 12540 4740 12549
rect 4420 12538 4444 12540
rect 4500 12538 4524 12540
rect 4580 12538 4604 12540
rect 4660 12538 4684 12540
rect 4420 12486 4430 12538
rect 4674 12486 4684 12538
rect 4420 12484 4444 12486
rect 4500 12484 4524 12486
rect 4580 12484 4604 12486
rect 4660 12484 4684 12486
rect 4364 12475 4740 12484
rect 4344 12300 4396 12306
rect 4344 12242 4396 12248
rect 4160 12164 4212 12170
rect 4160 12106 4212 12112
rect 4252 12164 4304 12170
rect 4252 12106 4304 12112
rect 3976 12096 4028 12102
rect 3976 12038 4028 12044
rect 4068 12096 4120 12102
rect 4068 12038 4120 12044
rect 3988 11558 4016 12038
rect 3976 11552 4028 11558
rect 3976 11494 4028 11500
rect 3988 10130 4016 11494
rect 4080 10198 4108 12038
rect 4172 11218 4200 12106
rect 4250 11792 4306 11801
rect 4356 11762 4384 12242
rect 4250 11727 4252 11736
rect 4304 11727 4306 11736
rect 4344 11756 4396 11762
rect 4252 11698 4304 11704
rect 4344 11698 4396 11704
rect 4252 11552 4304 11558
rect 4252 11494 4304 11500
rect 4160 11212 4212 11218
rect 4160 11154 4212 11160
rect 4264 10588 4292 11494
rect 4364 11452 4740 11461
rect 4420 11450 4444 11452
rect 4500 11450 4524 11452
rect 4580 11450 4604 11452
rect 4660 11450 4684 11452
rect 4420 11398 4430 11450
rect 4674 11398 4684 11450
rect 4420 11396 4444 11398
rect 4500 11396 4524 11398
rect 4580 11396 4604 11398
rect 4660 11396 4684 11398
rect 4364 11387 4740 11396
rect 4344 10600 4396 10606
rect 4264 10560 4344 10588
rect 4344 10542 4396 10548
rect 4364 10364 4740 10373
rect 4420 10362 4444 10364
rect 4500 10362 4524 10364
rect 4580 10362 4604 10364
rect 4660 10362 4684 10364
rect 4420 10310 4430 10362
rect 4674 10310 4684 10362
rect 4420 10308 4444 10310
rect 4500 10308 4524 10310
rect 4580 10308 4604 10310
rect 4660 10308 4684 10310
rect 4364 10299 4740 10308
rect 4068 10192 4120 10198
rect 4068 10134 4120 10140
rect 4342 10160 4398 10169
rect 3976 10124 4028 10130
rect 4342 10095 4398 10104
rect 3976 10066 4028 10072
rect 3988 9518 4016 10066
rect 4252 9920 4304 9926
rect 4252 9862 4304 9868
rect 4264 9654 4292 9862
rect 4068 9648 4120 9654
rect 4066 9616 4068 9625
rect 4252 9648 4304 9654
rect 4120 9616 4122 9625
rect 4252 9590 4304 9596
rect 4066 9551 4122 9560
rect 3976 9512 4028 9518
rect 3976 9454 4028 9460
rect 4160 9512 4212 9518
rect 4160 9454 4212 9460
rect 4068 9444 4120 9450
rect 4068 9386 4120 9392
rect 3976 9376 4028 9382
rect 3976 9318 4028 9324
rect 3988 9217 4016 9318
rect 3974 9208 4030 9217
rect 3974 9143 4030 9152
rect 4080 9042 4108 9386
rect 4172 9110 4200 9454
rect 4264 9178 4292 9590
rect 4356 9586 4384 10095
rect 4816 9722 4844 12668
rect 4896 12650 4948 12656
rect 5000 12646 5028 12718
rect 5092 12646 5120 12922
rect 5184 12646 5212 14418
rect 4988 12640 5040 12646
rect 4988 12582 5040 12588
rect 5080 12640 5132 12646
rect 5080 12582 5132 12588
rect 5172 12640 5224 12646
rect 5172 12582 5224 12588
rect 4896 12436 4948 12442
rect 4896 12378 4948 12384
rect 4908 11694 4936 12378
rect 5000 11762 5028 12582
rect 5276 12458 5304 14447
rect 5368 13462 5396 14606
rect 5448 14544 5500 14550
rect 5448 14486 5500 14492
rect 5356 13456 5408 13462
rect 5460 13444 5488 14486
rect 5552 14385 5580 14894
rect 5908 14816 5960 14822
rect 5908 14758 5960 14764
rect 5538 14376 5594 14385
rect 5538 14311 5594 14320
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5552 13841 5580 14214
rect 5538 13832 5594 13841
rect 5538 13767 5594 13776
rect 5540 13456 5592 13462
rect 5460 13416 5540 13444
rect 5356 13398 5408 13404
rect 5540 13398 5592 13404
rect 5356 13252 5408 13258
rect 5356 13194 5408 13200
rect 5184 12430 5304 12458
rect 5080 12300 5132 12306
rect 5080 12242 5132 12248
rect 5092 11898 5120 12242
rect 5080 11892 5132 11898
rect 5080 11834 5132 11840
rect 4988 11756 5040 11762
rect 4988 11698 5040 11704
rect 4896 11688 4948 11694
rect 4896 11630 4948 11636
rect 4988 11552 5040 11558
rect 4988 11494 5040 11500
rect 5080 11552 5132 11558
rect 5080 11494 5132 11500
rect 4896 11348 4948 11354
rect 4896 11290 4948 11296
rect 4804 9716 4856 9722
rect 4804 9658 4856 9664
rect 4344 9580 4396 9586
rect 4396 9540 4844 9568
rect 4344 9522 4396 9528
rect 4364 9276 4740 9285
rect 4420 9274 4444 9276
rect 4500 9274 4524 9276
rect 4580 9274 4604 9276
rect 4660 9274 4684 9276
rect 4420 9222 4430 9274
rect 4674 9222 4684 9274
rect 4420 9220 4444 9222
rect 4500 9220 4524 9222
rect 4580 9220 4604 9222
rect 4660 9220 4684 9222
rect 4364 9211 4740 9220
rect 4252 9172 4304 9178
rect 4252 9114 4304 9120
rect 4160 9104 4212 9110
rect 4160 9046 4212 9052
rect 4816 9042 4844 9540
rect 4068 9036 4120 9042
rect 4068 8978 4120 8984
rect 4804 9036 4856 9042
rect 4804 8978 4856 8984
rect 4160 8832 4212 8838
rect 4160 8774 4212 8780
rect 4068 8356 4120 8362
rect 4068 8298 4120 8304
rect 3976 8016 4028 8022
rect 3976 7958 4028 7964
rect 3804 7772 3924 7800
rect 3700 6860 3752 6866
rect 3700 6802 3752 6808
rect 3712 6458 3740 6802
rect 3700 6452 3752 6458
rect 3700 6394 3752 6400
rect 3804 5778 3832 7772
rect 3884 7404 3936 7410
rect 3884 7346 3936 7352
rect 3792 5772 3844 5778
rect 3792 5714 3844 5720
rect 3606 5672 3662 5681
rect 3606 5607 3662 5616
rect 3608 5296 3660 5302
rect 3608 5238 3660 5244
rect 3516 5024 3568 5030
rect 3516 4966 3568 4972
rect 3528 4826 3556 4966
rect 3516 4820 3568 4826
rect 3516 4762 3568 4768
rect 3424 4072 3476 4078
rect 3424 4014 3476 4020
rect 3148 3936 3200 3942
rect 3148 3878 3200 3884
rect 3160 3602 3188 3878
rect 3148 3596 3200 3602
rect 3148 3538 3200 3544
rect 3056 3528 3108 3534
rect 3056 3470 3108 3476
rect 3148 2984 3200 2990
rect 3148 2926 3200 2932
rect 3160 2378 3188 2926
rect 3332 2576 3384 2582
rect 3332 2518 3384 2524
rect 3148 2372 3200 2378
rect 3148 2314 3200 2320
rect 3344 2106 3372 2518
rect 3436 2514 3464 4014
rect 3424 2508 3476 2514
rect 3424 2450 3476 2456
rect 3332 2100 3384 2106
rect 3332 2042 3384 2048
rect 2504 1964 2556 1970
rect 2504 1906 2556 1912
rect 3436 1902 3464 2450
rect 1952 1896 2004 1902
rect 1952 1838 2004 1844
rect 3056 1896 3108 1902
rect 3056 1838 3108 1844
rect 3424 1896 3476 1902
rect 3424 1838 3476 1844
rect 2688 1760 2740 1766
rect 2688 1702 2740 1708
rect 2780 1760 2832 1766
rect 2780 1702 2832 1708
rect 2228 1556 2280 1562
rect 2228 1498 2280 1504
rect 1860 1420 1912 1426
rect 1860 1362 1912 1368
rect 1952 1420 2004 1426
rect 1952 1362 2004 1368
rect 1768 1216 1820 1222
rect 1768 1158 1820 1164
rect 1364 1116 1740 1125
rect 1420 1114 1444 1116
rect 1500 1114 1524 1116
rect 1580 1114 1604 1116
rect 1660 1114 1684 1116
rect 1420 1062 1430 1114
rect 1674 1062 1684 1114
rect 1420 1060 1444 1062
rect 1500 1060 1524 1062
rect 1580 1060 1604 1062
rect 1660 1060 1684 1062
rect 1364 1051 1740 1060
rect 1780 814 1808 1158
rect 1964 814 1992 1362
rect 1216 808 1268 814
rect 1216 750 1268 756
rect 1768 808 1820 814
rect 1768 750 1820 756
rect 1952 808 2004 814
rect 1952 750 2004 756
rect 1124 672 1176 678
rect 1124 614 1176 620
rect 1136 400 1164 614
rect 1228 406 1256 750
rect 1492 672 1544 678
rect 1492 614 1544 620
rect 1860 672 1912 678
rect 1860 614 1912 620
rect 1216 400 1268 406
rect 1504 400 1532 614
rect 1872 400 1900 614
rect 386 0 442 400
rect 754 0 810 400
rect 1122 0 1178 400
rect 1216 342 1268 348
rect 1490 0 1546 400
rect 1858 0 1914 400
rect 1964 202 1992 750
rect 2240 400 2268 1498
rect 2700 1494 2728 1702
rect 2688 1488 2740 1494
rect 2688 1430 2740 1436
rect 2792 1426 2820 1702
rect 2780 1420 2832 1426
rect 2780 1362 2832 1368
rect 2964 1216 3016 1222
rect 2964 1158 3016 1164
rect 2596 944 2648 950
rect 2596 886 2648 892
rect 2608 400 2636 886
rect 2976 400 3004 1158
rect 3068 950 3096 1838
rect 3332 1828 3384 1834
rect 3332 1770 3384 1776
rect 3344 1426 3372 1770
rect 3332 1420 3384 1426
rect 3332 1362 3384 1368
rect 3620 1358 3648 5238
rect 3792 5228 3844 5234
rect 3792 5170 3844 5176
rect 3804 4826 3832 5170
rect 3792 4820 3844 4826
rect 3792 4762 3844 4768
rect 3698 4720 3754 4729
rect 3698 4655 3700 4664
rect 3752 4655 3754 4664
rect 3700 4626 3752 4632
rect 3896 3126 3924 7346
rect 3988 5914 4016 7958
rect 4080 7002 4108 8298
rect 4068 6996 4120 7002
rect 4068 6938 4120 6944
rect 4172 6338 4200 8774
rect 4802 8664 4858 8673
rect 4802 8599 4804 8608
rect 4856 8599 4858 8608
rect 4804 8570 4856 8576
rect 4804 8492 4856 8498
rect 4804 8434 4856 8440
rect 4364 8188 4740 8197
rect 4420 8186 4444 8188
rect 4500 8186 4524 8188
rect 4580 8186 4604 8188
rect 4660 8186 4684 8188
rect 4420 8134 4430 8186
rect 4674 8134 4684 8186
rect 4420 8132 4444 8134
rect 4500 8132 4524 8134
rect 4580 8132 4604 8134
rect 4660 8132 4684 8134
rect 4364 8123 4740 8132
rect 4816 7886 4844 8434
rect 4908 8430 4936 11290
rect 5000 11218 5028 11494
rect 4988 11212 5040 11218
rect 4988 11154 5040 11160
rect 5000 9110 5028 11154
rect 4988 9104 5040 9110
rect 4988 9046 5040 9052
rect 4896 8424 4948 8430
rect 4894 8392 4896 8401
rect 4948 8392 4950 8401
rect 4894 8327 4950 8336
rect 4896 8288 4948 8294
rect 4896 8230 4948 8236
rect 4908 8022 4936 8230
rect 4896 8016 4948 8022
rect 4896 7958 4948 7964
rect 4804 7880 4856 7886
rect 4804 7822 4856 7828
rect 4252 7336 4304 7342
rect 4252 7278 4304 7284
rect 4896 7336 4948 7342
rect 4896 7278 4948 7284
rect 4264 6866 4292 7278
rect 4804 7200 4856 7206
rect 4804 7142 4856 7148
rect 4364 7100 4740 7109
rect 4420 7098 4444 7100
rect 4500 7098 4524 7100
rect 4580 7098 4604 7100
rect 4660 7098 4684 7100
rect 4420 7046 4430 7098
rect 4674 7046 4684 7098
rect 4420 7044 4444 7046
rect 4500 7044 4524 7046
rect 4580 7044 4604 7046
rect 4660 7044 4684 7046
rect 4364 7035 4740 7044
rect 4436 6996 4488 7002
rect 4436 6938 4488 6944
rect 4448 6866 4476 6938
rect 4816 6866 4844 7142
rect 4908 6934 4936 7278
rect 4896 6928 4948 6934
rect 4896 6870 4948 6876
rect 4252 6860 4304 6866
rect 4252 6802 4304 6808
rect 4436 6860 4488 6866
rect 4436 6802 4488 6808
rect 4804 6860 4856 6866
rect 4804 6802 4856 6808
rect 4528 6656 4580 6662
rect 4528 6598 4580 6604
rect 4080 6322 4200 6338
rect 4540 6322 4568 6598
rect 4068 6316 4200 6322
rect 4120 6310 4200 6316
rect 4528 6316 4580 6322
rect 4068 6258 4120 6264
rect 4528 6258 4580 6264
rect 4364 6012 4740 6021
rect 4420 6010 4444 6012
rect 4500 6010 4524 6012
rect 4580 6010 4604 6012
rect 4660 6010 4684 6012
rect 4420 5958 4430 6010
rect 4674 5958 4684 6010
rect 4420 5956 4444 5958
rect 4500 5956 4524 5958
rect 4580 5956 4604 5958
rect 4660 5956 4684 5958
rect 4364 5947 4740 5956
rect 3976 5908 4028 5914
rect 4160 5908 4212 5914
rect 4028 5868 4108 5896
rect 3976 5850 4028 5856
rect 3976 5772 4028 5778
rect 3976 5714 4028 5720
rect 3988 5574 4016 5714
rect 3976 5568 4028 5574
rect 3976 5510 4028 5516
rect 3988 5166 4016 5510
rect 3976 5160 4028 5166
rect 3976 5102 4028 5108
rect 4080 4690 4108 5868
rect 4160 5850 4212 5856
rect 4172 4690 4200 5850
rect 4528 5772 4580 5778
rect 4528 5714 4580 5720
rect 4620 5772 4672 5778
rect 4620 5714 4672 5720
rect 4804 5772 4856 5778
rect 4804 5714 4856 5720
rect 4344 5636 4396 5642
rect 4344 5578 4396 5584
rect 4252 5568 4304 5574
rect 4252 5510 4304 5516
rect 4068 4684 4120 4690
rect 4068 4626 4120 4632
rect 4160 4684 4212 4690
rect 4160 4626 4212 4632
rect 4172 4146 4200 4626
rect 4264 4622 4292 5510
rect 4356 5137 4384 5578
rect 4540 5574 4568 5714
rect 4528 5568 4580 5574
rect 4528 5510 4580 5516
rect 4632 5370 4660 5714
rect 4620 5364 4672 5370
rect 4620 5306 4672 5312
rect 4342 5128 4398 5137
rect 4342 5063 4398 5072
rect 4364 4924 4740 4933
rect 4420 4922 4444 4924
rect 4500 4922 4524 4924
rect 4580 4922 4604 4924
rect 4660 4922 4684 4924
rect 4420 4870 4430 4922
rect 4674 4870 4684 4922
rect 4420 4868 4444 4870
rect 4500 4868 4524 4870
rect 4580 4868 4604 4870
rect 4660 4868 4684 4870
rect 4364 4859 4740 4868
rect 4816 4826 4844 5714
rect 5000 5166 5028 9046
rect 5092 7936 5120 11494
rect 5184 8566 5212 12430
rect 5264 12164 5316 12170
rect 5264 12106 5316 12112
rect 5276 11121 5304 12106
rect 5368 11898 5396 13194
rect 5448 13184 5500 13190
rect 5448 13126 5500 13132
rect 5460 12209 5488 13126
rect 5552 12714 5580 13398
rect 5540 12708 5592 12714
rect 5540 12650 5592 12656
rect 5446 12200 5502 12209
rect 5446 12135 5502 12144
rect 5356 11892 5408 11898
rect 5356 11834 5408 11840
rect 5356 11620 5408 11626
rect 5356 11562 5408 11568
rect 5262 11112 5318 11121
rect 5262 11047 5318 11056
rect 5264 10600 5316 10606
rect 5264 10542 5316 10548
rect 5276 10266 5304 10542
rect 5264 10260 5316 10266
rect 5264 10202 5316 10208
rect 5264 9376 5316 9382
rect 5264 9318 5316 9324
rect 5172 8560 5224 8566
rect 5172 8502 5224 8508
rect 5092 7908 5212 7936
rect 5080 7812 5132 7818
rect 5080 7754 5132 7760
rect 5092 5710 5120 7754
rect 5184 7478 5212 7908
rect 5172 7472 5224 7478
rect 5172 7414 5224 7420
rect 5172 7200 5224 7206
rect 5172 7142 5224 7148
rect 5184 5914 5212 7142
rect 5172 5908 5224 5914
rect 5172 5850 5224 5856
rect 5080 5704 5132 5710
rect 5080 5646 5132 5652
rect 5184 5522 5212 5850
rect 5092 5494 5212 5522
rect 4988 5160 5040 5166
rect 4988 5102 5040 5108
rect 4896 5024 4948 5030
rect 4896 4966 4948 4972
rect 4804 4820 4856 4826
rect 4804 4762 4856 4768
rect 4908 4758 4936 4966
rect 4528 4752 4580 4758
rect 4342 4720 4398 4729
rect 4528 4694 4580 4700
rect 4896 4752 4948 4758
rect 4896 4694 4948 4700
rect 4342 4655 4398 4664
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 4160 4140 4212 4146
rect 4160 4082 4212 4088
rect 4356 4078 4384 4655
rect 4540 4078 4568 4694
rect 4896 4616 4948 4622
rect 4896 4558 4948 4564
rect 4908 4078 4936 4558
rect 4988 4548 5040 4554
rect 4988 4490 5040 4496
rect 5000 4282 5028 4490
rect 4988 4276 5040 4282
rect 4988 4218 5040 4224
rect 4344 4072 4396 4078
rect 4344 4014 4396 4020
rect 4528 4072 4580 4078
rect 4528 4014 4580 4020
rect 4896 4072 4948 4078
rect 4988 4072 5040 4078
rect 4896 4014 4948 4020
rect 4986 4040 4988 4049
rect 5040 4040 5042 4049
rect 4986 3975 5042 3984
rect 4344 3936 4396 3942
rect 4264 3896 4344 3924
rect 4264 3602 4292 3896
rect 4344 3878 4396 3884
rect 4364 3836 4740 3845
rect 4420 3834 4444 3836
rect 4500 3834 4524 3836
rect 4580 3834 4604 3836
rect 4660 3834 4684 3836
rect 4420 3782 4430 3834
rect 4674 3782 4684 3834
rect 4420 3780 4444 3782
rect 4500 3780 4524 3782
rect 4580 3780 4604 3782
rect 4660 3780 4684 3782
rect 4364 3771 4740 3780
rect 4252 3596 4304 3602
rect 4252 3538 4304 3544
rect 3884 3120 3936 3126
rect 3884 3062 3936 3068
rect 4264 2990 4292 3538
rect 4620 3392 4672 3398
rect 4620 3334 4672 3340
rect 4632 3058 4660 3334
rect 4986 3088 5042 3097
rect 4620 3052 4672 3058
rect 4986 3023 4988 3032
rect 4620 2994 4672 3000
rect 5040 3023 5042 3032
rect 4988 2994 5040 3000
rect 4252 2984 4304 2990
rect 4252 2926 4304 2932
rect 4252 2848 4304 2854
rect 4252 2790 4304 2796
rect 3884 2440 3936 2446
rect 3884 2382 3936 2388
rect 3896 2038 3924 2382
rect 3976 2304 4028 2310
rect 3976 2246 4028 2252
rect 3884 2032 3936 2038
rect 3884 1974 3936 1980
rect 3988 1766 4016 2246
rect 3976 1760 4028 1766
rect 3976 1702 4028 1708
rect 4160 1760 4212 1766
rect 4160 1702 4212 1708
rect 3608 1352 3660 1358
rect 3608 1294 3660 1300
rect 3332 1012 3384 1018
rect 3332 954 3384 960
rect 3056 944 3108 950
rect 3056 886 3108 892
rect 1952 196 2004 202
rect 1952 138 2004 144
rect 2226 0 2282 400
rect 2594 0 2650 400
rect 2962 0 3018 400
rect 3068 338 3096 886
rect 3344 400 3372 954
rect 4068 944 4120 950
rect 4068 886 4120 892
rect 3424 808 3476 814
rect 3424 750 3476 756
rect 3056 332 3108 338
rect 3056 274 3108 280
rect 3330 0 3386 400
rect 3436 270 3464 750
rect 3700 672 3752 678
rect 3700 614 3752 620
rect 3712 400 3740 614
rect 4080 400 4108 886
rect 4172 814 4200 1702
rect 4264 1426 4292 2790
rect 4364 2748 4740 2757
rect 4420 2746 4444 2748
rect 4500 2746 4524 2748
rect 4580 2746 4604 2748
rect 4660 2746 4684 2748
rect 4420 2694 4430 2746
rect 4674 2694 4684 2746
rect 4420 2692 4444 2694
rect 4500 2692 4524 2694
rect 4580 2692 4604 2694
rect 4660 2692 4684 2694
rect 4364 2683 4740 2692
rect 5092 2650 5120 5494
rect 5276 5250 5304 9318
rect 5368 9081 5396 11562
rect 5552 11558 5580 12650
rect 5920 12434 5948 14758
rect 5998 14648 6054 14657
rect 6196 14618 6224 14894
rect 6288 14890 6316 15438
rect 6472 15434 6500 15914
rect 6564 15570 6592 15982
rect 6644 15700 6696 15706
rect 6644 15642 6696 15648
rect 6656 15609 6684 15642
rect 6642 15600 6698 15609
rect 6552 15564 6604 15570
rect 6642 15535 6698 15544
rect 6552 15506 6604 15512
rect 6460 15428 6512 15434
rect 6460 15370 6512 15376
rect 6368 15360 6420 15366
rect 6368 15302 6420 15308
rect 6276 14884 6328 14890
rect 6276 14826 6328 14832
rect 5998 14583 6054 14592
rect 6184 14612 6236 14618
rect 5736 12406 5948 12434
rect 5540 11552 5592 11558
rect 5540 11494 5592 11500
rect 5448 11212 5500 11218
rect 5448 11154 5500 11160
rect 5460 10810 5488 11154
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5354 9072 5410 9081
rect 5354 9007 5410 9016
rect 5356 8968 5408 8974
rect 5356 8910 5408 8916
rect 5368 8498 5396 8910
rect 5356 8492 5408 8498
rect 5356 8434 5408 8440
rect 5356 7336 5408 7342
rect 5356 7278 5408 7284
rect 5368 5846 5396 7278
rect 5460 6746 5488 10202
rect 5540 9988 5592 9994
rect 5540 9930 5592 9936
rect 5552 9518 5580 9930
rect 5632 9920 5684 9926
rect 5632 9862 5684 9868
rect 5644 9518 5672 9862
rect 5736 9674 5764 12406
rect 5908 12232 5960 12238
rect 6012 12220 6040 14583
rect 6184 14554 6236 14560
rect 6092 14476 6144 14482
rect 6092 14418 6144 14424
rect 6104 13977 6132 14418
rect 6090 13968 6146 13977
rect 6090 13903 6146 13912
rect 6184 13524 6236 13530
rect 6184 13466 6236 13472
rect 6196 13258 6224 13466
rect 6184 13252 6236 13258
rect 6184 13194 6236 13200
rect 6196 12714 6224 13194
rect 6276 12912 6328 12918
rect 6276 12854 6328 12860
rect 6184 12708 6236 12714
rect 6184 12650 6236 12656
rect 6288 12442 6316 12854
rect 6276 12436 6328 12442
rect 6276 12378 6328 12384
rect 5960 12192 6040 12220
rect 5908 12174 5960 12180
rect 5816 12164 5868 12170
rect 5816 12106 5868 12112
rect 5828 11558 5856 12106
rect 6092 11688 6144 11694
rect 6092 11630 6144 11636
rect 5816 11552 5868 11558
rect 5816 11494 5868 11500
rect 5828 10198 5856 11494
rect 5908 11212 5960 11218
rect 5908 11154 5960 11160
rect 5920 10674 5948 11154
rect 6104 11150 6132 11630
rect 6092 11144 6144 11150
rect 6380 11098 6408 15302
rect 6564 15162 6592 15506
rect 6552 15156 6604 15162
rect 6552 15098 6604 15104
rect 6460 15088 6512 15094
rect 6458 15056 6460 15065
rect 6512 15056 6514 15065
rect 6458 14991 6514 15000
rect 6564 14618 6592 15098
rect 6552 14612 6604 14618
rect 6552 14554 6604 14560
rect 6748 14550 6776 16050
rect 6920 16040 6972 16046
rect 7024 16028 7052 16594
rect 7116 16538 7144 17020
rect 7300 16794 7328 17478
rect 7364 17436 7740 17445
rect 7420 17434 7444 17436
rect 7500 17434 7524 17436
rect 7580 17434 7604 17436
rect 7660 17434 7684 17436
rect 7420 17382 7430 17434
rect 7674 17382 7684 17434
rect 7420 17380 7444 17382
rect 7500 17380 7524 17382
rect 7580 17380 7604 17382
rect 7660 17380 7684 17382
rect 7364 17371 7740 17380
rect 7852 16794 7880 17546
rect 7944 17338 7972 17614
rect 7932 17332 7984 17338
rect 7932 17274 7984 17280
rect 7288 16788 7340 16794
rect 7288 16730 7340 16736
rect 7840 16788 7892 16794
rect 7840 16730 7892 16736
rect 7472 16652 7524 16658
rect 7472 16594 7524 16600
rect 7748 16652 7800 16658
rect 7748 16594 7800 16600
rect 7484 16561 7512 16594
rect 7286 16552 7342 16561
rect 7116 16510 7236 16538
rect 7104 16448 7156 16454
rect 7104 16390 7156 16396
rect 6972 16000 7052 16028
rect 6920 15982 6972 15988
rect 7116 15570 7144 16390
rect 7208 16114 7236 16510
rect 7286 16487 7342 16496
rect 7470 16552 7526 16561
rect 7760 16522 7788 16594
rect 7470 16487 7526 16496
rect 7748 16516 7800 16522
rect 7196 16108 7248 16114
rect 7196 16050 7248 16056
rect 7300 15994 7328 16487
rect 7748 16458 7800 16464
rect 7364 16348 7740 16357
rect 7420 16346 7444 16348
rect 7500 16346 7524 16348
rect 7580 16346 7604 16348
rect 7660 16346 7684 16348
rect 7420 16294 7430 16346
rect 7674 16294 7684 16346
rect 7420 16292 7444 16294
rect 7500 16292 7524 16294
rect 7580 16292 7604 16294
rect 7660 16292 7684 16294
rect 7364 16283 7740 16292
rect 7852 16046 7880 16730
rect 8220 16250 8248 17750
rect 8404 17746 8432 18294
rect 8392 17740 8444 17746
rect 8392 17682 8444 17688
rect 8484 17740 8536 17746
rect 8484 17682 8536 17688
rect 8208 16244 8260 16250
rect 8208 16186 8260 16192
rect 8220 16046 8248 16186
rect 7840 16040 7892 16046
rect 7196 15972 7248 15978
rect 7300 15966 7420 15994
rect 7840 15982 7892 15988
rect 8208 16040 8260 16046
rect 8208 15982 8260 15988
rect 7196 15914 7248 15920
rect 7104 15564 7156 15570
rect 7104 15506 7156 15512
rect 6920 15428 6972 15434
rect 6920 15370 6972 15376
rect 6932 14958 6960 15370
rect 6920 14952 6972 14958
rect 6920 14894 6972 14900
rect 6920 14816 6972 14822
rect 6920 14758 6972 14764
rect 7012 14816 7064 14822
rect 7012 14758 7064 14764
rect 6736 14544 6788 14550
rect 6736 14486 6788 14492
rect 6828 14068 6880 14074
rect 6932 14056 6960 14758
rect 7024 14362 7052 14758
rect 7116 14482 7144 15506
rect 7208 15162 7236 15914
rect 7288 15904 7340 15910
rect 7288 15846 7340 15852
rect 7196 15156 7248 15162
rect 7196 15098 7248 15104
rect 7104 14476 7156 14482
rect 7104 14418 7156 14424
rect 7024 14334 7144 14362
rect 7012 14272 7064 14278
rect 7012 14214 7064 14220
rect 6880 14028 6960 14056
rect 6828 14010 6880 14016
rect 6932 13462 6960 14028
rect 6920 13456 6972 13462
rect 6920 13398 6972 13404
rect 6826 13288 6882 13297
rect 6826 13223 6882 13232
rect 6840 12850 6868 13223
rect 6828 12844 6880 12850
rect 6828 12786 6880 12792
rect 6920 12844 6972 12850
rect 6920 12786 6972 12792
rect 6460 12640 6512 12646
rect 6460 12582 6512 12588
rect 6736 12640 6788 12646
rect 6736 12582 6788 12588
rect 6092 11086 6144 11092
rect 6104 10962 6132 11086
rect 6012 10934 6132 10962
rect 6288 11070 6408 11098
rect 6012 10674 6040 10934
rect 6092 10736 6144 10742
rect 6092 10678 6144 10684
rect 5908 10668 5960 10674
rect 5908 10610 5960 10616
rect 6000 10668 6052 10674
rect 6000 10610 6052 10616
rect 5816 10192 5868 10198
rect 5816 10134 5868 10140
rect 5736 9646 5856 9674
rect 5540 9512 5592 9518
rect 5540 9454 5592 9460
rect 5632 9512 5684 9518
rect 5632 9454 5684 9460
rect 5552 8838 5580 9454
rect 5644 9042 5672 9454
rect 5632 9036 5684 9042
rect 5632 8978 5684 8984
rect 5630 8936 5686 8945
rect 5630 8871 5686 8880
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 5538 7032 5594 7041
rect 5538 6967 5594 6976
rect 5552 6866 5580 6967
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 5460 6718 5580 6746
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 5460 6254 5488 6598
rect 5448 6248 5500 6254
rect 5448 6190 5500 6196
rect 5356 5840 5408 5846
rect 5356 5782 5408 5788
rect 5552 5778 5580 6718
rect 5540 5772 5592 5778
rect 5540 5714 5592 5720
rect 5540 5636 5592 5642
rect 5540 5578 5592 5584
rect 5276 5222 5396 5250
rect 5368 5166 5396 5222
rect 5552 5166 5580 5578
rect 5644 5216 5672 8871
rect 5722 8664 5778 8673
rect 5722 8599 5724 8608
rect 5776 8599 5778 8608
rect 5724 8570 5776 8576
rect 5828 7954 5856 9646
rect 6104 9586 6132 10678
rect 6184 10600 6236 10606
rect 6184 10542 6236 10548
rect 6196 10198 6224 10542
rect 6184 10192 6236 10198
rect 6184 10134 6236 10140
rect 6288 9602 6316 11070
rect 6472 10554 6500 12582
rect 6748 12306 6776 12582
rect 6736 12300 6788 12306
rect 6736 12242 6788 12248
rect 6644 12096 6696 12102
rect 6644 12038 6696 12044
rect 6552 11076 6604 11082
rect 6552 11018 6604 11024
rect 6564 10810 6592 11018
rect 6552 10804 6604 10810
rect 6552 10746 6604 10752
rect 6550 10704 6606 10713
rect 6550 10639 6606 10648
rect 6564 10606 6592 10639
rect 6092 9580 6144 9586
rect 6092 9522 6144 9528
rect 6196 9574 6316 9602
rect 6380 10526 6500 10554
rect 6552 10600 6604 10606
rect 6552 10542 6604 10548
rect 6196 9110 6224 9574
rect 6380 9518 6408 10526
rect 6460 10464 6512 10470
rect 6460 10406 6512 10412
rect 6276 9512 6328 9518
rect 6276 9454 6328 9460
rect 6368 9512 6420 9518
rect 6368 9454 6420 9460
rect 6288 9178 6316 9454
rect 6276 9172 6328 9178
rect 6276 9114 6328 9120
rect 6184 9104 6236 9110
rect 6184 9046 6236 9052
rect 6274 9072 6330 9081
rect 5908 9036 5960 9042
rect 5908 8978 5960 8984
rect 5816 7948 5868 7954
rect 5816 7890 5868 7896
rect 5816 7336 5868 7342
rect 5920 7324 5948 8978
rect 6196 8514 6224 9046
rect 6274 9007 6330 9016
rect 6104 8486 6224 8514
rect 6104 8430 6132 8486
rect 6288 8430 6316 9007
rect 6380 8974 6408 9454
rect 6368 8968 6420 8974
rect 6368 8910 6420 8916
rect 6368 8492 6420 8498
rect 6368 8434 6420 8440
rect 6092 8424 6144 8430
rect 6276 8424 6328 8430
rect 6092 8366 6144 8372
rect 6196 8384 6276 8412
rect 6092 8288 6144 8294
rect 6092 8230 6144 8236
rect 6104 7410 6132 8230
rect 6092 7404 6144 7410
rect 6092 7346 6144 7352
rect 5868 7296 5948 7324
rect 5816 7278 5868 7284
rect 5724 7200 5776 7206
rect 5724 7142 5776 7148
rect 5736 6458 5764 7142
rect 5816 6996 5868 7002
rect 5816 6938 5868 6944
rect 5828 6458 5856 6938
rect 5920 6882 5948 7296
rect 6000 7336 6052 7342
rect 6000 7278 6052 7284
rect 6012 7002 6040 7278
rect 6000 6996 6052 7002
rect 6000 6938 6052 6944
rect 5920 6854 6040 6882
rect 6196 6866 6224 8384
rect 6276 8366 6328 8372
rect 6274 7984 6330 7993
rect 6380 7954 6408 8434
rect 6274 7919 6276 7928
rect 6328 7919 6330 7928
rect 6368 7948 6420 7954
rect 6276 7890 6328 7896
rect 6368 7890 6420 7896
rect 6276 7744 6328 7750
rect 6276 7686 6328 7692
rect 6288 7002 6316 7686
rect 6366 7440 6422 7449
rect 6366 7375 6422 7384
rect 6276 6996 6328 7002
rect 6276 6938 6328 6944
rect 5908 6656 5960 6662
rect 5908 6598 5960 6604
rect 5920 6458 5948 6598
rect 5724 6452 5776 6458
rect 5724 6394 5776 6400
rect 5816 6452 5868 6458
rect 5816 6394 5868 6400
rect 5908 6452 5960 6458
rect 5908 6394 5960 6400
rect 5828 5760 5856 6394
rect 6012 6254 6040 6854
rect 6184 6860 6236 6866
rect 6184 6802 6236 6808
rect 6380 6730 6408 7375
rect 6472 7041 6500 10406
rect 6564 10130 6592 10542
rect 6552 10124 6604 10130
rect 6552 10066 6604 10072
rect 6552 9512 6604 9518
rect 6552 9454 6604 9460
rect 6564 9081 6592 9454
rect 6550 9072 6606 9081
rect 6550 9007 6606 9016
rect 6552 8628 6604 8634
rect 6552 8570 6604 8576
rect 6564 8022 6592 8570
rect 6552 8016 6604 8022
rect 6552 7958 6604 7964
rect 6564 7313 6592 7958
rect 6550 7304 6606 7313
rect 6550 7239 6606 7248
rect 6552 7200 6604 7206
rect 6552 7142 6604 7148
rect 6458 7032 6514 7041
rect 6458 6967 6514 6976
rect 6458 6760 6514 6769
rect 6368 6724 6420 6730
rect 6564 6730 6592 7142
rect 6458 6695 6460 6704
rect 6368 6666 6420 6672
rect 6512 6695 6514 6704
rect 6552 6724 6604 6730
rect 6460 6666 6512 6672
rect 6552 6666 6604 6672
rect 6000 6248 6052 6254
rect 6000 6190 6052 6196
rect 6092 6248 6144 6254
rect 6092 6190 6144 6196
rect 6276 6248 6328 6254
rect 6276 6190 6328 6196
rect 6104 5846 6132 6190
rect 6288 5914 6316 6190
rect 6276 5908 6328 5914
rect 6276 5850 6328 5856
rect 6092 5840 6144 5846
rect 6092 5782 6144 5788
rect 5908 5772 5960 5778
rect 5828 5732 5908 5760
rect 5908 5714 5960 5720
rect 6380 5710 6408 6666
rect 6552 6112 6604 6118
rect 6552 6054 6604 6060
rect 6460 5772 6512 5778
rect 6460 5714 6512 5720
rect 6368 5704 6420 5710
rect 6368 5646 6420 5652
rect 6000 5636 6052 5642
rect 6000 5578 6052 5584
rect 5644 5188 5764 5216
rect 5264 5160 5316 5166
rect 5264 5102 5316 5108
rect 5356 5160 5408 5166
rect 5356 5102 5408 5108
rect 5448 5160 5500 5166
rect 5448 5102 5500 5108
rect 5540 5160 5592 5166
rect 5540 5102 5592 5108
rect 5172 5024 5224 5030
rect 5172 4966 5224 4972
rect 5184 3602 5212 4966
rect 5276 4826 5304 5102
rect 5356 5024 5408 5030
rect 5356 4966 5408 4972
rect 5264 4820 5316 4826
rect 5264 4762 5316 4768
rect 5368 4622 5396 4966
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 5264 4480 5316 4486
rect 5264 4422 5316 4428
rect 5276 4078 5304 4422
rect 5368 4282 5396 4558
rect 5356 4276 5408 4282
rect 5356 4218 5408 4224
rect 5460 4078 5488 5102
rect 5632 5092 5684 5098
rect 5632 5034 5684 5040
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 5264 4072 5316 4078
rect 5264 4014 5316 4020
rect 5448 4072 5500 4078
rect 5448 4014 5500 4020
rect 5356 4004 5408 4010
rect 5356 3946 5408 3952
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 5368 2990 5396 3946
rect 5356 2984 5408 2990
rect 5356 2926 5408 2932
rect 5552 2650 5580 4966
rect 5644 4826 5672 5034
rect 5632 4820 5684 4826
rect 5632 4762 5684 4768
rect 5736 4758 5764 5188
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 5724 4752 5776 4758
rect 5724 4694 5776 4700
rect 5920 4554 5948 5102
rect 5908 4548 5960 4554
rect 5908 4490 5960 4496
rect 6012 3126 6040 5578
rect 6368 5568 6420 5574
rect 6368 5510 6420 5516
rect 6184 5024 6236 5030
rect 6184 4966 6236 4972
rect 6196 4690 6224 4966
rect 6184 4684 6236 4690
rect 6184 4626 6236 4632
rect 6092 4140 6144 4146
rect 6092 4082 6144 4088
rect 6104 3670 6132 4082
rect 6196 3670 6224 4626
rect 6276 4072 6328 4078
rect 6276 4014 6328 4020
rect 6092 3664 6144 3670
rect 6092 3606 6144 3612
rect 6184 3664 6236 3670
rect 6184 3606 6236 3612
rect 6288 3602 6316 4014
rect 6276 3596 6328 3602
rect 6276 3538 6328 3544
rect 6000 3120 6052 3126
rect 6000 3062 6052 3068
rect 5724 2984 5776 2990
rect 5724 2926 5776 2932
rect 5736 2650 5764 2926
rect 5816 2848 5868 2854
rect 5816 2790 5868 2796
rect 5080 2644 5132 2650
rect 5080 2586 5132 2592
rect 5540 2644 5592 2650
rect 5540 2586 5592 2592
rect 5724 2644 5776 2650
rect 5724 2586 5776 2592
rect 5736 1902 5764 2586
rect 5828 2446 5856 2790
rect 6000 2508 6052 2514
rect 6000 2450 6052 2456
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 5828 2106 5856 2382
rect 5816 2100 5868 2106
rect 5816 2042 5868 2048
rect 6012 1902 6040 2450
rect 6184 2372 6236 2378
rect 6184 2314 6236 2320
rect 6196 1970 6224 2314
rect 6184 1964 6236 1970
rect 6184 1906 6236 1912
rect 4988 1896 5040 1902
rect 4988 1838 5040 1844
rect 5264 1896 5316 1902
rect 5264 1838 5316 1844
rect 5724 1896 5776 1902
rect 5724 1838 5776 1844
rect 6000 1896 6052 1902
rect 6000 1838 6052 1844
rect 4896 1760 4948 1766
rect 4896 1702 4948 1708
rect 4364 1660 4740 1669
rect 4420 1658 4444 1660
rect 4500 1658 4524 1660
rect 4580 1658 4604 1660
rect 4660 1658 4684 1660
rect 4420 1606 4430 1658
rect 4674 1606 4684 1658
rect 4420 1604 4444 1606
rect 4500 1604 4524 1606
rect 4580 1604 4604 1606
rect 4660 1604 4684 1606
rect 4364 1595 4740 1604
rect 4252 1420 4304 1426
rect 4252 1362 4304 1368
rect 4908 814 4936 1702
rect 4160 808 4212 814
rect 4528 808 4580 814
rect 4160 750 4212 756
rect 4526 776 4528 785
rect 4896 808 4948 814
rect 4580 776 4582 785
rect 4896 750 4948 756
rect 5000 746 5028 1838
rect 5172 944 5224 950
rect 5172 886 5224 892
rect 4526 711 4582 720
rect 4988 740 5040 746
rect 4988 682 5040 688
rect 4252 672 4304 678
rect 4252 614 4304 620
rect 4804 672 4856 678
rect 4804 614 4856 620
rect 4264 456 4292 614
rect 4364 572 4740 581
rect 4420 570 4444 572
rect 4500 570 4524 572
rect 4580 570 4604 572
rect 4660 570 4684 572
rect 4420 518 4430 570
rect 4674 518 4684 570
rect 4420 516 4444 518
rect 4500 516 4524 518
rect 4580 516 4604 518
rect 4660 516 4684 518
rect 4364 507 4740 516
rect 4264 428 4476 456
rect 4448 400 4476 428
rect 4816 400 4844 614
rect 3424 264 3476 270
rect 3424 206 3476 212
rect 3698 0 3754 400
rect 4066 0 4122 400
rect 4434 0 4490 400
rect 4802 0 4858 400
rect 5000 202 5028 682
rect 5184 400 5212 886
rect 5276 785 5304 1838
rect 5448 1828 5500 1834
rect 5448 1770 5500 1776
rect 5460 1601 5488 1770
rect 5446 1592 5502 1601
rect 5446 1527 5502 1536
rect 5460 1494 5488 1527
rect 5448 1488 5500 1494
rect 5448 1430 5500 1436
rect 5736 1426 5764 1838
rect 5908 1760 5960 1766
rect 5908 1702 5960 1708
rect 5724 1420 5776 1426
rect 5724 1362 5776 1368
rect 5920 898 5948 1702
rect 6000 1420 6052 1426
rect 6000 1362 6052 1368
rect 6012 1018 6040 1362
rect 6380 1290 6408 5510
rect 6472 5098 6500 5714
rect 6460 5092 6512 5098
rect 6460 5034 6512 5040
rect 6564 2650 6592 6054
rect 6656 5710 6684 12038
rect 6828 11212 6880 11218
rect 6828 11154 6880 11160
rect 6840 10606 6868 11154
rect 6932 10810 6960 12786
rect 7024 12306 7052 14214
rect 7116 13462 7144 14334
rect 7104 13456 7156 13462
rect 7104 13398 7156 13404
rect 7208 12986 7236 15098
rect 7196 12980 7248 12986
rect 7196 12922 7248 12928
rect 7208 12782 7236 12922
rect 7196 12776 7248 12782
rect 7196 12718 7248 12724
rect 7300 12434 7328 15846
rect 7392 15706 7420 15966
rect 7840 15904 7892 15910
rect 7840 15846 7892 15852
rect 8024 15904 8076 15910
rect 8024 15846 8076 15852
rect 8298 15872 8354 15881
rect 7380 15700 7432 15706
rect 7380 15642 7432 15648
rect 7378 15600 7434 15609
rect 7378 15535 7380 15544
rect 7432 15535 7434 15544
rect 7380 15506 7432 15512
rect 7364 15260 7740 15269
rect 7420 15258 7444 15260
rect 7500 15258 7524 15260
rect 7580 15258 7604 15260
rect 7660 15258 7684 15260
rect 7420 15206 7430 15258
rect 7674 15206 7684 15258
rect 7420 15204 7444 15206
rect 7500 15204 7524 15206
rect 7580 15204 7604 15206
rect 7660 15204 7684 15206
rect 7364 15195 7740 15204
rect 7852 14958 7880 15846
rect 7932 15564 7984 15570
rect 7932 15506 7984 15512
rect 7840 14952 7892 14958
rect 7840 14894 7892 14900
rect 7472 14884 7524 14890
rect 7472 14826 7524 14832
rect 7484 14482 7512 14826
rect 7472 14476 7524 14482
rect 7472 14418 7524 14424
rect 7364 14172 7740 14181
rect 7420 14170 7444 14172
rect 7500 14170 7524 14172
rect 7580 14170 7604 14172
rect 7660 14170 7684 14172
rect 7420 14118 7430 14170
rect 7674 14118 7684 14170
rect 7420 14116 7444 14118
rect 7500 14116 7524 14118
rect 7580 14116 7604 14118
rect 7660 14116 7684 14118
rect 7364 14107 7740 14116
rect 7378 13968 7434 13977
rect 7378 13903 7434 13912
rect 7392 13870 7420 13903
rect 7380 13864 7432 13870
rect 7380 13806 7432 13812
rect 7656 13864 7708 13870
rect 7656 13806 7708 13812
rect 7564 13796 7616 13802
rect 7564 13738 7616 13744
rect 7472 13728 7524 13734
rect 7472 13670 7524 13676
rect 7484 13462 7512 13670
rect 7576 13530 7604 13738
rect 7564 13524 7616 13530
rect 7564 13466 7616 13472
rect 7472 13456 7524 13462
rect 7472 13398 7524 13404
rect 7668 13326 7696 13806
rect 7852 13530 7880 14894
rect 7944 14822 7972 15506
rect 7932 14816 7984 14822
rect 7932 14758 7984 14764
rect 7932 14544 7984 14550
rect 7932 14486 7984 14492
rect 7840 13524 7892 13530
rect 7840 13466 7892 13472
rect 7656 13320 7708 13326
rect 7654 13288 7656 13297
rect 7708 13288 7710 13297
rect 7654 13223 7710 13232
rect 7364 13084 7740 13093
rect 7420 13082 7444 13084
rect 7500 13082 7524 13084
rect 7580 13082 7604 13084
rect 7660 13082 7684 13084
rect 7420 13030 7430 13082
rect 7674 13030 7684 13082
rect 7420 13028 7444 13030
rect 7500 13028 7524 13030
rect 7580 13028 7604 13030
rect 7660 13028 7684 13030
rect 7364 13019 7740 13028
rect 7840 12912 7892 12918
rect 7840 12854 7892 12860
rect 7472 12776 7524 12782
rect 7472 12718 7524 12724
rect 7484 12442 7512 12718
rect 7208 12406 7328 12434
rect 7472 12436 7524 12442
rect 7012 12300 7064 12306
rect 7012 12242 7064 12248
rect 7012 12164 7064 12170
rect 7012 12106 7064 12112
rect 7024 11354 7052 12106
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 7012 11348 7064 11354
rect 7012 11290 7064 11296
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 7024 10538 7052 11290
rect 7116 11150 7144 12038
rect 7104 11144 7156 11150
rect 7104 11086 7156 11092
rect 7012 10532 7064 10538
rect 7012 10474 7064 10480
rect 7208 10418 7236 12406
rect 7472 12378 7524 12384
rect 7484 12306 7512 12378
rect 7472 12300 7524 12306
rect 7472 12242 7524 12248
rect 7364 11996 7740 12005
rect 7420 11994 7444 11996
rect 7500 11994 7524 11996
rect 7580 11994 7604 11996
rect 7660 11994 7684 11996
rect 7420 11942 7430 11994
rect 7674 11942 7684 11994
rect 7420 11940 7444 11942
rect 7500 11940 7524 11942
rect 7580 11940 7604 11942
rect 7660 11940 7684 11942
rect 7364 11931 7740 11940
rect 7288 11688 7340 11694
rect 7288 11630 7340 11636
rect 7300 11354 7328 11630
rect 7656 11620 7708 11626
rect 7656 11562 7708 11568
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 7288 11212 7340 11218
rect 7288 11154 7340 11160
rect 7300 10810 7328 11154
rect 7668 11150 7696 11562
rect 7564 11144 7616 11150
rect 7564 11086 7616 11092
rect 7656 11144 7708 11150
rect 7852 11121 7880 12854
rect 7656 11086 7708 11092
rect 7838 11112 7894 11121
rect 7576 11014 7604 11086
rect 7838 11047 7894 11056
rect 7564 11008 7616 11014
rect 7564 10950 7616 10956
rect 7364 10908 7740 10917
rect 7420 10906 7444 10908
rect 7500 10906 7524 10908
rect 7580 10906 7604 10908
rect 7660 10906 7684 10908
rect 7420 10854 7430 10906
rect 7674 10854 7684 10906
rect 7420 10852 7444 10854
rect 7500 10852 7524 10854
rect 7580 10852 7604 10854
rect 7660 10852 7684 10854
rect 7364 10843 7740 10852
rect 7288 10804 7340 10810
rect 7288 10746 7340 10752
rect 7748 10804 7800 10810
rect 7748 10746 7800 10752
rect 6840 10390 7236 10418
rect 6734 10160 6790 10169
rect 6734 10095 6790 10104
rect 6748 8498 6776 10095
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 6840 8022 6868 10390
rect 7104 10124 7156 10130
rect 7104 10066 7156 10072
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 7012 10056 7064 10062
rect 6918 10024 6974 10033
rect 7012 9998 7064 10004
rect 6918 9959 6974 9968
rect 6932 9042 6960 9959
rect 6920 9036 6972 9042
rect 6920 8978 6972 8984
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6828 8016 6880 8022
rect 6828 7958 6880 7964
rect 6932 7954 6960 8774
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 6932 7562 6960 7890
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 6840 7534 6960 7562
rect 6748 7449 6776 7482
rect 6734 7440 6790 7449
rect 6734 7375 6790 7384
rect 6736 7336 6788 7342
rect 6736 7278 6788 7284
rect 6748 6118 6776 7278
rect 6840 7274 6868 7534
rect 6920 7472 6972 7478
rect 6920 7414 6972 7420
rect 6828 7268 6880 7274
rect 6828 7210 6880 7216
rect 6826 7168 6882 7177
rect 6826 7103 6882 7112
rect 6840 6254 6868 7103
rect 6932 6798 6960 7414
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 6736 6112 6788 6118
rect 6736 6054 6788 6060
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 6656 5166 6684 5646
rect 6644 5160 6696 5166
rect 6644 5102 6696 5108
rect 6748 4622 6776 5850
rect 7024 5710 7052 9998
rect 7116 9450 7144 10066
rect 7196 9920 7248 9926
rect 7196 9862 7248 9868
rect 7208 9586 7236 9862
rect 7300 9722 7328 10066
rect 7760 9908 7788 10746
rect 7760 9880 7794 9908
rect 7766 9874 7794 9880
rect 7766 9846 7880 9874
rect 7364 9820 7740 9829
rect 7420 9818 7444 9820
rect 7500 9818 7524 9820
rect 7580 9818 7604 9820
rect 7660 9818 7684 9820
rect 7420 9766 7430 9818
rect 7674 9766 7684 9818
rect 7420 9764 7444 9766
rect 7500 9764 7524 9766
rect 7580 9764 7604 9766
rect 7660 9764 7684 9766
rect 7364 9755 7740 9764
rect 7288 9716 7340 9722
rect 7288 9658 7340 9664
rect 7564 9716 7616 9722
rect 7852 9704 7880 9846
rect 7564 9658 7616 9664
rect 7668 9676 7880 9704
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 7300 9450 7328 9658
rect 7576 9518 7604 9658
rect 7564 9512 7616 9518
rect 7564 9454 7616 9460
rect 7104 9444 7156 9450
rect 7104 9386 7156 9392
rect 7288 9444 7340 9450
rect 7288 9386 7340 9392
rect 7668 9217 7696 9676
rect 7654 9208 7710 9217
rect 7654 9143 7710 9152
rect 7840 9172 7892 9178
rect 7840 9114 7892 9120
rect 7104 9036 7156 9042
rect 7104 8978 7156 8984
rect 7288 9036 7340 9042
rect 7288 8978 7340 8984
rect 7116 8945 7144 8978
rect 7102 8936 7158 8945
rect 7102 8871 7158 8880
rect 7196 8900 7248 8906
rect 7196 8842 7248 8848
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 7116 8498 7144 8774
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 7116 7426 7144 8434
rect 7208 7954 7236 8842
rect 7196 7948 7248 7954
rect 7196 7890 7248 7896
rect 7196 7812 7248 7818
rect 7196 7754 7248 7760
rect 7208 7546 7236 7754
rect 7196 7540 7248 7546
rect 7196 7482 7248 7488
rect 7116 7410 7236 7426
rect 7116 7404 7248 7410
rect 7116 7398 7196 7404
rect 7196 7346 7248 7352
rect 7300 7342 7328 8978
rect 7748 8968 7800 8974
rect 7748 8910 7800 8916
rect 7760 8838 7788 8910
rect 7748 8832 7800 8838
rect 7852 8809 7880 9114
rect 7748 8774 7800 8780
rect 7838 8800 7894 8809
rect 7364 8732 7740 8741
rect 7838 8735 7894 8744
rect 7420 8730 7444 8732
rect 7500 8730 7524 8732
rect 7580 8730 7604 8732
rect 7660 8730 7684 8732
rect 7420 8678 7430 8730
rect 7674 8678 7684 8730
rect 7420 8676 7444 8678
rect 7500 8676 7524 8678
rect 7580 8676 7604 8678
rect 7660 8676 7684 8678
rect 7364 8667 7740 8676
rect 7748 8424 7800 8430
rect 7852 8412 7880 8735
rect 7800 8384 7880 8412
rect 7748 8366 7800 8372
rect 7564 7948 7616 7954
rect 7564 7890 7616 7896
rect 7470 7848 7526 7857
rect 7470 7783 7526 7792
rect 7484 7750 7512 7783
rect 7576 7750 7604 7890
rect 7760 7834 7788 8366
rect 7840 7948 7892 7954
rect 7944 7936 7972 14486
rect 8036 13705 8064 15846
rect 8298 15807 8354 15816
rect 8312 15638 8340 15807
rect 8300 15632 8352 15638
rect 8300 15574 8352 15580
rect 8298 15464 8354 15473
rect 8208 15428 8260 15434
rect 8298 15399 8354 15408
rect 8208 15370 8260 15376
rect 8116 15360 8168 15366
rect 8116 15302 8168 15308
rect 8128 14600 8156 15302
rect 8220 14793 8248 15370
rect 8312 15366 8340 15399
rect 8300 15360 8352 15366
rect 8300 15302 8352 15308
rect 8206 14784 8262 14793
rect 8206 14719 8262 14728
rect 8404 14618 8432 17682
rect 8496 16794 8524 17682
rect 8680 17338 8708 18584
rect 8772 18426 8800 19110
rect 8760 18420 8812 18426
rect 8760 18362 8812 18368
rect 8760 18148 8812 18154
rect 8760 18090 8812 18096
rect 8772 17882 8800 18090
rect 8760 17876 8812 17882
rect 8760 17818 8812 17824
rect 8668 17332 8720 17338
rect 8668 17274 8720 17280
rect 8576 16992 8628 16998
rect 8576 16934 8628 16940
rect 8760 16992 8812 16998
rect 8760 16934 8812 16940
rect 8484 16788 8536 16794
rect 8484 16730 8536 16736
rect 8588 16674 8616 16934
rect 8496 16646 8616 16674
rect 8666 16688 8722 16697
rect 8496 16590 8524 16646
rect 8666 16623 8722 16632
rect 8484 16584 8536 16590
rect 8680 16538 8708 16623
rect 8484 16526 8536 16532
rect 8496 16250 8524 16526
rect 8588 16510 8708 16538
rect 8484 16244 8536 16250
rect 8484 16186 8536 16192
rect 8484 15632 8536 15638
rect 8484 15574 8536 15580
rect 8496 15162 8524 15574
rect 8484 15156 8536 15162
rect 8484 15098 8536 15104
rect 8482 14784 8538 14793
rect 8482 14719 8538 14728
rect 8392 14612 8444 14618
rect 8128 14572 8340 14600
rect 8312 14521 8340 14572
rect 8392 14554 8444 14560
rect 8298 14512 8354 14521
rect 8208 14476 8260 14482
rect 8496 14482 8524 14719
rect 8298 14447 8354 14456
rect 8484 14476 8536 14482
rect 8208 14418 8260 14424
rect 8116 14000 8168 14006
rect 8114 13968 8116 13977
rect 8168 13968 8170 13977
rect 8114 13903 8170 13912
rect 8022 13696 8078 13705
rect 8022 13631 8078 13640
rect 8024 13524 8076 13530
rect 8024 13466 8076 13472
rect 8036 10810 8064 13466
rect 8220 12434 8248 14418
rect 8312 13734 8340 14447
rect 8484 14418 8536 14424
rect 8392 14272 8444 14278
rect 8392 14214 8444 14220
rect 8300 13728 8352 13734
rect 8300 13670 8352 13676
rect 8312 13394 8340 13670
rect 8300 13388 8352 13394
rect 8300 13330 8352 13336
rect 8298 12744 8354 12753
rect 8404 12714 8432 14214
rect 8588 12753 8616 16510
rect 8772 16250 8800 16934
rect 8760 16244 8812 16250
rect 8760 16186 8812 16192
rect 8668 15904 8720 15910
rect 8668 15846 8720 15852
rect 8680 13818 8708 15846
rect 8758 15736 8814 15745
rect 8758 15671 8814 15680
rect 8772 14822 8800 15671
rect 8864 15366 8892 19450
rect 8956 18834 8984 19654
rect 9048 19174 9076 19722
rect 9140 19281 9168 20862
rect 9126 19272 9182 19281
rect 9126 19207 9182 19216
rect 9220 19236 9272 19242
rect 9220 19178 9272 19184
rect 9036 19168 9088 19174
rect 9232 19145 9260 19178
rect 9036 19110 9088 19116
rect 9218 19136 9274 19145
rect 8944 18828 8996 18834
rect 8944 18770 8996 18776
rect 8944 18080 8996 18086
rect 8944 18022 8996 18028
rect 8956 17746 8984 18022
rect 9048 17882 9076 19110
rect 9218 19071 9274 19080
rect 9324 18970 9352 21422
rect 9692 21350 9720 21966
rect 9864 21956 9916 21962
rect 9864 21898 9916 21904
rect 9876 21486 9904 21898
rect 10060 21690 10088 22102
rect 10048 21684 10100 21690
rect 10048 21626 10100 21632
rect 9864 21480 9916 21486
rect 9864 21422 9916 21428
rect 10046 21448 10102 21457
rect 10046 21383 10102 21392
rect 9680 21344 9732 21350
rect 9680 21286 9732 21292
rect 9864 21344 9916 21350
rect 9864 21286 9916 21292
rect 9588 21140 9640 21146
rect 9588 21082 9640 21088
rect 9600 20942 9628 21082
rect 9692 21078 9720 21286
rect 9772 21140 9824 21146
rect 9772 21082 9824 21088
rect 9680 21072 9732 21078
rect 9680 21014 9732 21020
rect 9784 20942 9812 21082
rect 9876 21010 9904 21286
rect 10060 21010 10088 21383
rect 9864 21004 9916 21010
rect 9864 20946 9916 20952
rect 10048 21004 10100 21010
rect 10048 20946 10100 20952
rect 9588 20936 9640 20942
rect 9772 20936 9824 20942
rect 9640 20884 9720 20890
rect 9588 20878 9720 20884
rect 9772 20878 9824 20884
rect 9862 20904 9918 20913
rect 9600 20862 9720 20878
rect 9496 20800 9548 20806
rect 9496 20742 9548 20748
rect 9586 20768 9642 20777
rect 9508 20398 9536 20742
rect 9586 20703 9642 20712
rect 9496 20392 9548 20398
rect 9496 20334 9548 20340
rect 9404 19780 9456 19786
rect 9404 19722 9456 19728
rect 9416 19378 9444 19722
rect 9600 19378 9628 20703
rect 9692 19718 9720 20862
rect 9784 20602 9812 20878
rect 9862 20839 9918 20848
rect 9772 20596 9824 20602
rect 9772 20538 9824 20544
rect 9876 20398 9904 20839
rect 9954 20632 10010 20641
rect 9954 20567 10010 20576
rect 9968 20398 9996 20567
rect 9864 20392 9916 20398
rect 9864 20334 9916 20340
rect 9956 20392 10008 20398
rect 9956 20334 10008 20340
rect 9772 20256 9824 20262
rect 9772 20198 9824 20204
rect 9784 20058 9812 20198
rect 9772 20052 9824 20058
rect 9772 19994 9824 20000
rect 9784 19854 9812 19994
rect 9876 19922 9904 20334
rect 10152 20058 10180 22510
rect 10232 22432 10284 22438
rect 10232 22374 10284 22380
rect 10244 20602 10272 22374
rect 10364 22332 10740 22341
rect 10420 22330 10444 22332
rect 10500 22330 10524 22332
rect 10580 22330 10604 22332
rect 10660 22330 10684 22332
rect 10420 22278 10430 22330
rect 10674 22278 10684 22330
rect 10420 22276 10444 22278
rect 10500 22276 10524 22278
rect 10580 22276 10604 22278
rect 10660 22276 10684 22278
rect 10364 22267 10740 22276
rect 10980 22234 11008 23122
rect 11256 22778 11284 23122
rect 11244 22772 11296 22778
rect 11244 22714 11296 22720
rect 11244 22432 11296 22438
rect 11244 22374 11296 22380
rect 10968 22228 11020 22234
rect 10968 22170 11020 22176
rect 11256 22166 11284 22374
rect 11244 22160 11296 22166
rect 11244 22102 11296 22108
rect 10324 22092 10376 22098
rect 10324 22034 10376 22040
rect 10784 22092 10836 22098
rect 10784 22034 10836 22040
rect 10336 21486 10364 22034
rect 10796 21486 10824 22034
rect 11150 21584 11206 21593
rect 11150 21519 11206 21528
rect 10324 21480 10376 21486
rect 10324 21422 10376 21428
rect 10784 21480 10836 21486
rect 10784 21422 10836 21428
rect 10784 21344 10836 21350
rect 10784 21286 10836 21292
rect 10364 21244 10740 21253
rect 10420 21242 10444 21244
rect 10500 21242 10524 21244
rect 10580 21242 10604 21244
rect 10660 21242 10684 21244
rect 10420 21190 10430 21242
rect 10674 21190 10684 21242
rect 10420 21188 10444 21190
rect 10500 21188 10524 21190
rect 10580 21188 10604 21190
rect 10660 21188 10684 21190
rect 10364 21179 10740 21188
rect 10796 21078 10824 21286
rect 10784 21072 10836 21078
rect 10784 21014 10836 21020
rect 10692 21004 10744 21010
rect 10692 20946 10744 20952
rect 10324 20936 10376 20942
rect 10324 20878 10376 20884
rect 10232 20596 10284 20602
rect 10232 20538 10284 20544
rect 10336 20398 10364 20878
rect 10704 20602 10732 20946
rect 11060 20936 11112 20942
rect 11060 20878 11112 20884
rect 10692 20596 10744 20602
rect 10744 20556 10824 20584
rect 10692 20538 10744 20544
rect 10324 20392 10376 20398
rect 10324 20334 10376 20340
rect 10416 20392 10468 20398
rect 10416 20334 10468 20340
rect 10428 20244 10456 20334
rect 10244 20216 10456 20244
rect 10140 20052 10192 20058
rect 10140 19994 10192 20000
rect 9864 19916 9916 19922
rect 9864 19858 9916 19864
rect 9772 19848 9824 19854
rect 9772 19790 9824 19796
rect 9680 19712 9732 19718
rect 9680 19654 9732 19660
rect 9678 19544 9734 19553
rect 9784 19514 9812 19790
rect 9678 19479 9734 19488
rect 9772 19508 9824 19514
rect 9692 19378 9720 19479
rect 9772 19450 9824 19456
rect 9404 19372 9456 19378
rect 9404 19314 9456 19320
rect 9588 19372 9640 19378
rect 9588 19314 9640 19320
rect 9680 19372 9732 19378
rect 9680 19314 9732 19320
rect 9312 18964 9364 18970
rect 9312 18906 9364 18912
rect 9220 18828 9272 18834
rect 9220 18770 9272 18776
rect 9128 18080 9180 18086
rect 9232 18057 9260 18770
rect 9416 18766 9444 19314
rect 9864 19304 9916 19310
rect 9864 19246 9916 19252
rect 9956 19304 10008 19310
rect 9956 19246 10008 19252
rect 10048 19304 10100 19310
rect 10048 19246 10100 19252
rect 9876 19174 9904 19246
rect 9864 19168 9916 19174
rect 9862 19136 9864 19145
rect 9916 19136 9918 19145
rect 9862 19071 9918 19080
rect 9968 18834 9996 19246
rect 10060 18970 10088 19246
rect 10152 19242 10180 19994
rect 10140 19236 10192 19242
rect 10140 19178 10192 19184
rect 10048 18964 10100 18970
rect 10048 18906 10100 18912
rect 10152 18902 10180 19178
rect 10140 18896 10192 18902
rect 10140 18838 10192 18844
rect 9956 18828 10008 18834
rect 9956 18770 10008 18776
rect 9404 18760 9456 18766
rect 9404 18702 9456 18708
rect 9312 18624 9364 18630
rect 9312 18566 9364 18572
rect 9404 18624 9456 18630
rect 9404 18566 9456 18572
rect 9324 18329 9352 18566
rect 9310 18320 9366 18329
rect 9310 18255 9366 18264
rect 9310 18184 9366 18193
rect 9310 18119 9366 18128
rect 9128 18022 9180 18028
rect 9218 18048 9274 18057
rect 9036 17876 9088 17882
rect 9036 17818 9088 17824
rect 8944 17740 8996 17746
rect 8944 17682 8996 17688
rect 9140 17066 9168 18022
rect 9218 17983 9274 17992
rect 9324 17882 9352 18119
rect 9312 17876 9364 17882
rect 9312 17818 9364 17824
rect 9310 17776 9366 17785
rect 9310 17711 9366 17720
rect 9324 17202 9352 17711
rect 9312 17196 9364 17202
rect 9312 17138 9364 17144
rect 9128 17060 9180 17066
rect 9128 17002 9180 17008
rect 9036 16788 9088 16794
rect 9036 16730 9088 16736
rect 8944 16720 8996 16726
rect 8942 16688 8944 16697
rect 8996 16688 8998 16697
rect 8942 16623 8998 16632
rect 9048 16046 9076 16730
rect 9036 16040 9088 16046
rect 9036 15982 9088 15988
rect 9048 15570 9076 15982
rect 9140 15978 9168 17002
rect 9312 16992 9364 16998
rect 9312 16934 9364 16940
rect 9324 16658 9352 16934
rect 9312 16652 9364 16658
rect 9312 16594 9364 16600
rect 9128 15972 9180 15978
rect 9128 15914 9180 15920
rect 9036 15564 9088 15570
rect 9036 15506 9088 15512
rect 8852 15360 8904 15366
rect 8852 15302 8904 15308
rect 8942 15328 8998 15337
rect 8942 15263 8998 15272
rect 8850 14920 8906 14929
rect 8850 14855 8906 14864
rect 8760 14816 8812 14822
rect 8760 14758 8812 14764
rect 8864 14482 8892 14855
rect 8760 14476 8812 14482
rect 8760 14418 8812 14424
rect 8852 14476 8904 14482
rect 8852 14418 8904 14424
rect 8772 13938 8800 14418
rect 8760 13932 8812 13938
rect 8760 13874 8812 13880
rect 8956 13870 8984 15263
rect 9140 14890 9168 15914
rect 9416 15910 9444 18566
rect 9680 18352 9732 18358
rect 10244 18329 10272 20216
rect 10364 20156 10740 20165
rect 10420 20154 10444 20156
rect 10500 20154 10524 20156
rect 10580 20154 10604 20156
rect 10660 20154 10684 20156
rect 10420 20102 10430 20154
rect 10674 20102 10684 20154
rect 10420 20100 10444 20102
rect 10500 20100 10524 20102
rect 10580 20100 10604 20102
rect 10660 20100 10684 20102
rect 10364 20091 10740 20100
rect 10416 20052 10468 20058
rect 10416 19994 10468 20000
rect 10428 19718 10456 19994
rect 10416 19712 10468 19718
rect 10416 19654 10468 19660
rect 10506 19680 10562 19689
rect 10428 19514 10456 19654
rect 10506 19615 10562 19624
rect 10416 19508 10468 19514
rect 10416 19450 10468 19456
rect 10520 19378 10548 19615
rect 10796 19446 10824 20556
rect 11072 20262 11100 20878
rect 11060 20256 11112 20262
rect 10966 20224 11022 20233
rect 11060 20198 11112 20204
rect 10966 20159 11022 20168
rect 10876 19984 10928 19990
rect 10876 19926 10928 19932
rect 10784 19440 10836 19446
rect 10784 19382 10836 19388
rect 10508 19372 10560 19378
rect 10508 19314 10560 19320
rect 10364 19068 10740 19077
rect 10420 19066 10444 19068
rect 10500 19066 10524 19068
rect 10580 19066 10604 19068
rect 10660 19066 10684 19068
rect 10420 19014 10430 19066
rect 10674 19014 10684 19066
rect 10420 19012 10444 19014
rect 10500 19012 10524 19014
rect 10580 19012 10604 19014
rect 10660 19012 10684 19014
rect 10364 19003 10740 19012
rect 10508 18828 10560 18834
rect 10508 18770 10560 18776
rect 10416 18624 10468 18630
rect 10416 18566 10468 18572
rect 9680 18294 9732 18300
rect 10230 18320 10286 18329
rect 9496 18216 9548 18222
rect 9496 18158 9548 18164
rect 9508 17218 9536 18158
rect 9588 18148 9640 18154
rect 9588 18090 9640 18096
rect 9600 17338 9628 18090
rect 9692 17746 9720 18294
rect 10230 18255 10286 18264
rect 10428 18222 10456 18566
rect 10520 18426 10548 18770
rect 10508 18420 10560 18426
rect 10508 18362 10560 18368
rect 10416 18216 10468 18222
rect 10416 18158 10468 18164
rect 10140 18148 10192 18154
rect 10140 18090 10192 18096
rect 9772 18080 9824 18086
rect 9772 18022 9824 18028
rect 9680 17740 9732 17746
rect 9680 17682 9732 17688
rect 9588 17332 9640 17338
rect 9588 17274 9640 17280
rect 9784 17270 9812 18022
rect 9772 17264 9824 17270
rect 9508 17190 9628 17218
rect 9772 17206 9824 17212
rect 9600 17134 9628 17190
rect 9588 17128 9640 17134
rect 9588 17070 9640 17076
rect 9600 16998 9628 17070
rect 9956 17060 10008 17066
rect 9956 17002 10008 17008
rect 9588 16992 9640 16998
rect 9588 16934 9640 16940
rect 9404 15904 9456 15910
rect 9404 15846 9456 15852
rect 9494 15872 9550 15881
rect 9494 15807 9550 15816
rect 9508 15706 9536 15807
rect 9496 15700 9548 15706
rect 9496 15642 9548 15648
rect 9600 15638 9628 16934
rect 9968 16794 9996 17002
rect 9956 16788 10008 16794
rect 9956 16730 10008 16736
rect 10152 16590 10180 18090
rect 10364 17980 10740 17989
rect 10420 17978 10444 17980
rect 10500 17978 10524 17980
rect 10580 17978 10604 17980
rect 10660 17978 10684 17980
rect 10420 17926 10430 17978
rect 10674 17926 10684 17978
rect 10420 17924 10444 17926
rect 10500 17924 10524 17926
rect 10580 17924 10604 17926
rect 10660 17924 10684 17926
rect 10364 17915 10740 17924
rect 10796 17066 10824 19382
rect 10888 17202 10916 19926
rect 10980 19922 11008 20159
rect 10968 19916 11020 19922
rect 10968 19858 11020 19864
rect 11164 19174 11192 21519
rect 11244 21004 11296 21010
rect 11244 20946 11296 20952
rect 11256 20398 11284 20946
rect 11244 20392 11296 20398
rect 11244 20334 11296 20340
rect 11152 19168 11204 19174
rect 11152 19110 11204 19116
rect 10968 18828 11020 18834
rect 10968 18770 11020 18776
rect 11060 18828 11112 18834
rect 11060 18770 11112 18776
rect 10980 17746 11008 18770
rect 11072 18154 11100 18770
rect 11348 18408 11376 23122
rect 11520 22568 11572 22574
rect 11520 22510 11572 22516
rect 11532 22234 11560 22510
rect 11520 22228 11572 22234
rect 11520 22170 11572 22176
rect 11428 22092 11480 22098
rect 11428 22034 11480 22040
rect 11440 21486 11468 22034
rect 11428 21480 11480 21486
rect 11428 21422 11480 21428
rect 11520 21480 11572 21486
rect 11520 21422 11572 21428
rect 11428 21344 11480 21350
rect 11428 21286 11480 21292
rect 11440 20602 11468 21286
rect 11532 20913 11560 21422
rect 11704 21344 11756 21350
rect 11704 21286 11756 21292
rect 11716 21146 11744 21286
rect 11704 21140 11756 21146
rect 11704 21082 11756 21088
rect 11808 21078 11836 23122
rect 12624 22568 12676 22574
rect 12624 22510 12676 22516
rect 11980 22432 12032 22438
rect 11980 22374 12032 22380
rect 12256 22432 12308 22438
rect 12256 22374 12308 22380
rect 11992 21554 12020 22374
rect 12268 22166 12296 22374
rect 12256 22160 12308 22166
rect 12256 22102 12308 22108
rect 12532 22092 12584 22098
rect 12532 22034 12584 22040
rect 12544 21894 12572 22034
rect 12636 21894 12664 22510
rect 12728 21962 12756 23600
rect 13176 22976 13228 22982
rect 13176 22918 13228 22924
rect 13188 22574 13216 22918
rect 13176 22568 13228 22574
rect 13176 22510 13228 22516
rect 13174 21992 13230 22001
rect 12716 21956 12768 21962
rect 13280 21962 13308 23600
rect 17224 23598 17276 23604
rect 16364 23420 16740 23429
rect 16420 23418 16444 23420
rect 16500 23418 16524 23420
rect 16580 23418 16604 23420
rect 16660 23418 16684 23420
rect 16420 23366 16430 23418
rect 16674 23366 16684 23418
rect 16420 23364 16444 23366
rect 16500 23364 16524 23366
rect 16580 23364 16604 23366
rect 16660 23364 16684 23366
rect 16364 23355 16740 23364
rect 15844 23316 15896 23322
rect 15844 23258 15896 23264
rect 14832 23180 14884 23186
rect 14832 23122 14884 23128
rect 15660 23180 15712 23186
rect 15660 23122 15712 23128
rect 13820 23112 13872 23118
rect 13820 23054 13872 23060
rect 13364 22876 13740 22885
rect 13420 22874 13444 22876
rect 13500 22874 13524 22876
rect 13580 22874 13604 22876
rect 13660 22874 13684 22876
rect 13420 22822 13430 22874
rect 13674 22822 13684 22874
rect 13420 22820 13444 22822
rect 13500 22820 13524 22822
rect 13580 22820 13604 22822
rect 13660 22820 13684 22822
rect 13364 22811 13740 22820
rect 13832 22710 13860 23054
rect 14464 22976 14516 22982
rect 14464 22918 14516 22924
rect 13820 22704 13872 22710
rect 13820 22646 13872 22652
rect 14372 22704 14424 22710
rect 14372 22646 14424 22652
rect 13452 22568 13504 22574
rect 13452 22510 13504 22516
rect 13464 22166 13492 22510
rect 13636 22500 13688 22506
rect 13636 22442 13688 22448
rect 13648 22166 13676 22442
rect 14280 22432 14332 22438
rect 14280 22374 14332 22380
rect 13452 22160 13504 22166
rect 13452 22102 13504 22108
rect 13636 22160 13688 22166
rect 13636 22102 13688 22108
rect 13728 22092 13780 22098
rect 13728 22034 13780 22040
rect 14188 22092 14240 22098
rect 14188 22034 14240 22040
rect 13174 21927 13230 21936
rect 13268 21956 13320 21962
rect 12716 21898 12768 21904
rect 12072 21888 12124 21894
rect 12532 21888 12584 21894
rect 12072 21830 12124 21836
rect 12530 21856 12532 21865
rect 12624 21888 12676 21894
rect 12584 21856 12586 21865
rect 11980 21548 12032 21554
rect 11980 21490 12032 21496
rect 11980 21412 12032 21418
rect 11980 21354 12032 21360
rect 11796 21072 11848 21078
rect 11796 21014 11848 21020
rect 11518 20904 11574 20913
rect 11518 20839 11574 20848
rect 11428 20596 11480 20602
rect 11428 20538 11480 20544
rect 11440 20505 11468 20538
rect 11532 20534 11560 20839
rect 11520 20528 11572 20534
rect 11426 20496 11482 20505
rect 11520 20470 11572 20476
rect 11808 20466 11836 21014
rect 11992 21010 12020 21354
rect 12084 21010 12112 21830
rect 12624 21830 12676 21836
rect 12530 21791 12586 21800
rect 12636 21486 12664 21830
rect 13188 21486 13216 21927
rect 13268 21898 13320 21904
rect 13740 21876 13768 22034
rect 13740 21865 13860 21876
rect 13740 21856 13874 21865
rect 13740 21848 13818 21856
rect 13364 21788 13740 21797
rect 13818 21791 13874 21800
rect 13420 21786 13444 21788
rect 13500 21786 13524 21788
rect 13580 21786 13604 21788
rect 13660 21786 13684 21788
rect 13420 21734 13430 21786
rect 13674 21734 13684 21786
rect 13420 21732 13444 21734
rect 13500 21732 13524 21734
rect 13580 21732 13604 21734
rect 13660 21732 13684 21734
rect 13364 21723 13740 21732
rect 14200 21690 14228 22034
rect 14292 22030 14320 22374
rect 14384 22166 14412 22646
rect 14476 22574 14504 22918
rect 14464 22568 14516 22574
rect 14464 22510 14516 22516
rect 14556 22500 14608 22506
rect 14556 22442 14608 22448
rect 14372 22160 14424 22166
rect 14372 22102 14424 22108
rect 14280 22024 14332 22030
rect 14280 21966 14332 21972
rect 14188 21684 14240 21690
rect 14188 21626 14240 21632
rect 12624 21480 12676 21486
rect 12624 21422 12676 21428
rect 13176 21480 13228 21486
rect 14188 21480 14240 21486
rect 13176 21422 13228 21428
rect 13910 21448 13966 21457
rect 14188 21422 14240 21428
rect 14280 21480 14332 21486
rect 14280 21422 14332 21428
rect 14372 21480 14424 21486
rect 14372 21422 14424 21428
rect 14464 21480 14516 21486
rect 14464 21422 14516 21428
rect 13910 21383 13966 21392
rect 14096 21412 14148 21418
rect 13924 21350 13952 21383
rect 14096 21354 14148 21360
rect 12716 21344 12768 21350
rect 12716 21286 12768 21292
rect 12808 21344 12860 21350
rect 12808 21286 12860 21292
rect 13912 21344 13964 21350
rect 13912 21286 13964 21292
rect 12164 21140 12216 21146
rect 12164 21082 12216 21088
rect 11980 21004 12032 21010
rect 11980 20946 12032 20952
rect 12072 21004 12124 21010
rect 12072 20946 12124 20952
rect 12072 20868 12124 20874
rect 12072 20810 12124 20816
rect 11426 20431 11482 20440
rect 11796 20460 11848 20466
rect 11848 20420 11928 20448
rect 11796 20402 11848 20408
rect 11520 20392 11572 20398
rect 11520 20334 11572 20340
rect 11428 20256 11480 20262
rect 11428 20198 11480 20204
rect 11440 20058 11468 20198
rect 11532 20058 11560 20334
rect 11428 20052 11480 20058
rect 11428 19994 11480 20000
rect 11520 20052 11572 20058
rect 11520 19994 11572 20000
rect 11796 20052 11848 20058
rect 11796 19994 11848 20000
rect 11808 19378 11836 19994
rect 11900 19854 11928 20420
rect 12084 20330 12112 20810
rect 12176 20806 12204 21082
rect 12622 20904 12678 20913
rect 12622 20839 12678 20848
rect 12164 20800 12216 20806
rect 12532 20800 12584 20806
rect 12164 20742 12216 20748
rect 12530 20768 12532 20777
rect 12584 20768 12586 20777
rect 12530 20703 12586 20712
rect 12072 20324 12124 20330
rect 12072 20266 12124 20272
rect 12636 20262 12664 20839
rect 12728 20584 12756 21286
rect 12820 20777 12848 21286
rect 14108 21078 14136 21354
rect 14096 21072 14148 21078
rect 14096 21014 14148 21020
rect 13268 21004 13320 21010
rect 13268 20946 13320 20952
rect 13820 21004 13872 21010
rect 13820 20946 13872 20952
rect 12806 20768 12862 20777
rect 12806 20703 12862 20712
rect 13280 20602 13308 20946
rect 13364 20700 13740 20709
rect 13420 20698 13444 20700
rect 13500 20698 13524 20700
rect 13580 20698 13604 20700
rect 13660 20698 13684 20700
rect 13420 20646 13430 20698
rect 13674 20646 13684 20698
rect 13420 20644 13444 20646
rect 13500 20644 13524 20646
rect 13580 20644 13604 20646
rect 13660 20644 13684 20646
rect 13364 20635 13740 20644
rect 12808 20596 12860 20602
rect 12728 20556 12808 20584
rect 12808 20538 12860 20544
rect 13268 20596 13320 20602
rect 13268 20538 13320 20544
rect 13832 20466 13860 20946
rect 14200 20942 14228 21422
rect 14188 20936 14240 20942
rect 14188 20878 14240 20884
rect 14096 20868 14148 20874
rect 14096 20810 14148 20816
rect 13820 20460 13872 20466
rect 13820 20402 13872 20408
rect 14108 20398 14136 20810
rect 14096 20392 14148 20398
rect 14096 20334 14148 20340
rect 14292 20330 14320 21422
rect 14384 20806 14412 21422
rect 14372 20800 14424 20806
rect 14372 20742 14424 20748
rect 14476 20602 14504 21422
rect 14568 20602 14596 22442
rect 14844 22166 14872 23122
rect 15016 22704 15068 22710
rect 15016 22646 15068 22652
rect 15476 22704 15528 22710
rect 15476 22646 15528 22652
rect 15028 22166 15056 22646
rect 15200 22568 15252 22574
rect 15200 22510 15252 22516
rect 15108 22432 15160 22438
rect 15108 22374 15160 22380
rect 14832 22160 14884 22166
rect 14832 22102 14884 22108
rect 15016 22160 15068 22166
rect 15120 22137 15148 22374
rect 15016 22102 15068 22108
rect 15106 22128 15162 22137
rect 15106 22063 15162 22072
rect 15016 21888 15068 21894
rect 15016 21830 15068 21836
rect 14740 21480 14792 21486
rect 14740 21422 14792 21428
rect 14752 21162 14780 21422
rect 14660 21134 14780 21162
rect 14464 20596 14516 20602
rect 14464 20538 14516 20544
rect 14556 20596 14608 20602
rect 14556 20538 14608 20544
rect 14280 20324 14332 20330
rect 14280 20266 14332 20272
rect 12624 20256 12676 20262
rect 12624 20198 12676 20204
rect 13084 20052 13136 20058
rect 13084 19994 13136 20000
rect 14372 20052 14424 20058
rect 14372 19994 14424 20000
rect 12072 19916 12124 19922
rect 11992 19876 12072 19904
rect 11888 19848 11940 19854
rect 11888 19790 11940 19796
rect 11888 19440 11940 19446
rect 11888 19382 11940 19388
rect 11796 19372 11848 19378
rect 11796 19314 11848 19320
rect 11808 19242 11836 19314
rect 11900 19242 11928 19382
rect 11796 19236 11848 19242
rect 11796 19178 11848 19184
rect 11888 19236 11940 19242
rect 11888 19178 11940 19184
rect 11808 18698 11836 19178
rect 11992 19174 12020 19876
rect 12072 19858 12124 19864
rect 12532 19916 12584 19922
rect 12532 19858 12584 19864
rect 12072 19712 12124 19718
rect 12072 19654 12124 19660
rect 12084 19242 12112 19654
rect 12072 19236 12124 19242
rect 12072 19178 12124 19184
rect 11980 19168 12032 19174
rect 11980 19110 12032 19116
rect 12440 19168 12492 19174
rect 12440 19110 12492 19116
rect 11992 18834 12020 19110
rect 12452 18834 12480 19110
rect 12544 18970 12572 19858
rect 12808 19508 12860 19514
rect 12808 19450 12860 19456
rect 12532 18964 12584 18970
rect 12532 18906 12584 18912
rect 11980 18828 12032 18834
rect 11980 18770 12032 18776
rect 12072 18828 12124 18834
rect 12072 18770 12124 18776
rect 12348 18828 12400 18834
rect 12348 18770 12400 18776
rect 12440 18828 12492 18834
rect 12440 18770 12492 18776
rect 12532 18828 12584 18834
rect 12532 18770 12584 18776
rect 11520 18692 11572 18698
rect 11520 18634 11572 18640
rect 11796 18692 11848 18698
rect 11796 18634 11848 18640
rect 11256 18380 11376 18408
rect 11060 18148 11112 18154
rect 11112 18108 11192 18136
rect 11060 18090 11112 18096
rect 10968 17740 11020 17746
rect 10968 17682 11020 17688
rect 11060 17740 11112 17746
rect 11060 17682 11112 17688
rect 11072 17338 11100 17682
rect 11060 17332 11112 17338
rect 11060 17274 11112 17280
rect 10876 17196 10928 17202
rect 10876 17138 10928 17144
rect 10784 17060 10836 17066
rect 10784 17002 10836 17008
rect 10364 16892 10740 16901
rect 10420 16890 10444 16892
rect 10500 16890 10524 16892
rect 10580 16890 10604 16892
rect 10660 16890 10684 16892
rect 10420 16838 10430 16890
rect 10674 16838 10684 16890
rect 10420 16836 10444 16838
rect 10500 16836 10524 16838
rect 10580 16836 10604 16838
rect 10660 16836 10684 16838
rect 10364 16827 10740 16836
rect 10598 16688 10654 16697
rect 10598 16623 10600 16632
rect 10652 16623 10654 16632
rect 10784 16652 10836 16658
rect 10600 16594 10652 16600
rect 10784 16594 10836 16600
rect 10140 16584 10192 16590
rect 10140 16526 10192 16532
rect 9680 16448 9732 16454
rect 9680 16390 9732 16396
rect 10416 16448 10468 16454
rect 10416 16390 10468 16396
rect 9692 16250 9720 16390
rect 9680 16244 9732 16250
rect 9680 16186 9732 16192
rect 9956 16244 10008 16250
rect 9956 16186 10008 16192
rect 9772 16176 9824 16182
rect 9772 16118 9824 16124
rect 9680 16040 9732 16046
rect 9680 15982 9732 15988
rect 9588 15632 9640 15638
rect 9588 15574 9640 15580
rect 9692 15570 9720 15982
rect 9784 15570 9812 16118
rect 9968 15892 9996 16186
rect 10428 16114 10456 16390
rect 10612 16250 10640 16594
rect 10692 16584 10744 16590
rect 10692 16526 10744 16532
rect 10600 16244 10652 16250
rect 10600 16186 10652 16192
rect 10704 16130 10732 16526
rect 10796 16250 10824 16594
rect 10968 16448 11020 16454
rect 10968 16390 11020 16396
rect 10784 16244 10836 16250
rect 10784 16186 10836 16192
rect 10416 16108 10468 16114
rect 10704 16102 10824 16130
rect 10416 16050 10468 16056
rect 10048 16040 10100 16046
rect 10048 15982 10100 15988
rect 10232 16040 10284 16046
rect 10232 15982 10284 15988
rect 9876 15864 9996 15892
rect 9680 15564 9732 15570
rect 9680 15506 9732 15512
rect 9772 15564 9824 15570
rect 9772 15506 9824 15512
rect 9220 15496 9272 15502
rect 9220 15438 9272 15444
rect 9312 15496 9364 15502
rect 9312 15438 9364 15444
rect 9404 15496 9456 15502
rect 9456 15444 9536 15450
rect 9404 15438 9536 15444
rect 9232 15162 9260 15438
rect 9220 15156 9272 15162
rect 9220 15098 9272 15104
rect 9324 15026 9352 15438
rect 9416 15422 9536 15438
rect 9404 15360 9456 15366
rect 9404 15302 9456 15308
rect 9312 15020 9364 15026
rect 9312 14962 9364 14968
rect 9128 14884 9180 14890
rect 9128 14826 9180 14832
rect 9036 14816 9088 14822
rect 9036 14758 9088 14764
rect 9048 14521 9076 14758
rect 9034 14512 9090 14521
rect 9034 14447 9090 14456
rect 8944 13864 8996 13870
rect 8680 13790 8800 13818
rect 8996 13824 9076 13852
rect 8944 13806 8996 13812
rect 8668 13728 8720 13734
rect 8668 13670 8720 13676
rect 8680 13530 8708 13670
rect 8668 13524 8720 13530
rect 8668 13466 8720 13472
rect 8772 12986 8800 13790
rect 8942 13560 8998 13569
rect 8942 13495 8998 13504
rect 8760 12980 8812 12986
rect 8760 12922 8812 12928
rect 8668 12776 8720 12782
rect 8574 12744 8630 12753
rect 8298 12679 8354 12688
rect 8392 12708 8444 12714
rect 8312 12646 8340 12679
rect 8668 12718 8720 12724
rect 8574 12679 8630 12688
rect 8392 12650 8444 12656
rect 8300 12640 8352 12646
rect 8300 12582 8352 12588
rect 8128 12406 8248 12434
rect 8680 12434 8708 12718
rect 8852 12640 8904 12646
rect 8852 12582 8904 12588
rect 8680 12406 8800 12434
rect 8024 10804 8076 10810
rect 8024 10746 8076 10752
rect 8024 9920 8076 9926
rect 8024 9862 8076 9868
rect 8036 9518 8064 9862
rect 8024 9512 8076 9518
rect 8024 9454 8076 9460
rect 7892 7908 7972 7936
rect 7840 7890 7892 7896
rect 7760 7806 7880 7834
rect 7472 7744 7524 7750
rect 7472 7686 7524 7692
rect 7564 7744 7616 7750
rect 7564 7686 7616 7692
rect 7364 7644 7740 7653
rect 7420 7642 7444 7644
rect 7500 7642 7524 7644
rect 7580 7642 7604 7644
rect 7660 7642 7684 7644
rect 7420 7590 7430 7642
rect 7674 7590 7684 7642
rect 7420 7588 7444 7590
rect 7500 7588 7524 7590
rect 7580 7588 7604 7590
rect 7660 7588 7684 7590
rect 7364 7579 7740 7588
rect 7852 7528 7880 7806
rect 7932 7812 7984 7818
rect 7932 7754 7984 7760
rect 7668 7500 7880 7528
rect 7668 7342 7696 7500
rect 7748 7404 7800 7410
rect 7800 7364 7880 7392
rect 7748 7346 7800 7352
rect 7288 7336 7340 7342
rect 7288 7278 7340 7284
rect 7656 7336 7708 7342
rect 7656 7278 7708 7284
rect 7104 7268 7156 7274
rect 7104 7210 7156 7216
rect 7116 6254 7144 7210
rect 7196 7200 7248 7206
rect 7196 7142 7248 7148
rect 7472 7200 7524 7206
rect 7472 7142 7524 7148
rect 7208 6866 7236 7142
rect 7484 6934 7512 7142
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 7472 6928 7524 6934
rect 7472 6870 7524 6876
rect 7196 6860 7248 6866
rect 7248 6820 7328 6848
rect 7196 6802 7248 6808
rect 7196 6656 7248 6662
rect 7196 6598 7248 6604
rect 7208 6497 7236 6598
rect 7194 6488 7250 6497
rect 7194 6423 7250 6432
rect 7208 6254 7236 6423
rect 7104 6248 7156 6254
rect 7104 6190 7156 6196
rect 7196 6248 7248 6254
rect 7196 6190 7248 6196
rect 7196 5840 7248 5846
rect 7196 5782 7248 5788
rect 7012 5704 7064 5710
rect 7012 5646 7064 5652
rect 6920 5568 6972 5574
rect 6920 5510 6972 5516
rect 6828 5296 6880 5302
rect 6828 5238 6880 5244
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 6840 3942 6868 5238
rect 6932 5166 6960 5510
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 7012 5160 7064 5166
rect 7012 5102 7064 5108
rect 6920 5024 6972 5030
rect 6920 4966 6972 4972
rect 6932 4706 6960 4966
rect 7024 4826 7052 5102
rect 7208 5098 7236 5782
rect 7196 5092 7248 5098
rect 7196 5034 7248 5040
rect 7012 4820 7064 4826
rect 7012 4762 7064 4768
rect 7196 4752 7248 4758
rect 6932 4678 7052 4706
rect 7196 4694 7248 4700
rect 7024 4622 7052 4678
rect 7012 4616 7064 4622
rect 7012 4558 7064 4564
rect 7024 4282 7052 4558
rect 7012 4276 7064 4282
rect 7012 4218 7064 4224
rect 7104 4208 7156 4214
rect 7104 4150 7156 4156
rect 7116 4078 7144 4150
rect 7104 4072 7156 4078
rect 7104 4014 7156 4020
rect 6828 3936 6880 3942
rect 6828 3878 6880 3884
rect 7208 3194 7236 4694
rect 7300 3602 7328 6820
rect 7760 6662 7788 6938
rect 7748 6656 7800 6662
rect 7748 6598 7800 6604
rect 7364 6556 7740 6565
rect 7420 6554 7444 6556
rect 7500 6554 7524 6556
rect 7580 6554 7604 6556
rect 7660 6554 7684 6556
rect 7420 6502 7430 6554
rect 7674 6502 7684 6554
rect 7420 6500 7444 6502
rect 7500 6500 7524 6502
rect 7580 6500 7604 6502
rect 7660 6500 7684 6502
rect 7364 6491 7740 6500
rect 7852 6390 7880 7364
rect 7840 6384 7892 6390
rect 7840 6326 7892 6332
rect 7748 6248 7800 6254
rect 7748 6190 7800 6196
rect 7840 6248 7892 6254
rect 7840 6190 7892 6196
rect 7380 6180 7432 6186
rect 7380 6122 7432 6128
rect 7392 5642 7420 6122
rect 7760 6089 7788 6190
rect 7746 6080 7802 6089
rect 7746 6015 7802 6024
rect 7760 5914 7788 6015
rect 7748 5908 7800 5914
rect 7748 5850 7800 5856
rect 7380 5636 7432 5642
rect 7380 5578 7432 5584
rect 7364 5468 7740 5477
rect 7420 5466 7444 5468
rect 7500 5466 7524 5468
rect 7580 5466 7604 5468
rect 7660 5466 7684 5468
rect 7420 5414 7430 5466
rect 7674 5414 7684 5466
rect 7420 5412 7444 5414
rect 7500 5412 7524 5414
rect 7580 5412 7604 5414
rect 7660 5412 7684 5414
rect 7364 5403 7740 5412
rect 7852 5250 7880 6190
rect 7668 5222 7880 5250
rect 7668 5166 7696 5222
rect 7656 5160 7708 5166
rect 7944 5114 7972 7754
rect 7656 5102 7708 5108
rect 7668 4758 7696 5102
rect 7852 5086 7972 5114
rect 7656 4752 7708 4758
rect 7656 4694 7708 4700
rect 7852 4622 7880 5086
rect 7932 5024 7984 5030
rect 7932 4966 7984 4972
rect 7840 4616 7892 4622
rect 7840 4558 7892 4564
rect 7840 4480 7892 4486
rect 7840 4422 7892 4428
rect 7364 4380 7740 4389
rect 7420 4378 7444 4380
rect 7500 4378 7524 4380
rect 7580 4378 7604 4380
rect 7660 4378 7684 4380
rect 7420 4326 7430 4378
rect 7674 4326 7684 4378
rect 7420 4324 7444 4326
rect 7500 4324 7524 4326
rect 7580 4324 7604 4326
rect 7660 4324 7684 4326
rect 7364 4315 7740 4324
rect 7852 4282 7880 4422
rect 7656 4276 7708 4282
rect 7656 4218 7708 4224
rect 7840 4276 7892 4282
rect 7840 4218 7892 4224
rect 7668 4162 7696 4218
rect 7668 4134 7788 4162
rect 7656 4072 7708 4078
rect 7484 4032 7656 4060
rect 7484 3942 7512 4032
rect 7656 4014 7708 4020
rect 7760 3942 7788 4134
rect 7472 3936 7524 3942
rect 7472 3878 7524 3884
rect 7748 3936 7800 3942
rect 7748 3878 7800 3884
rect 7944 3738 7972 4966
rect 8036 4282 8064 9454
rect 8128 9178 8156 12406
rect 8484 12368 8536 12374
rect 8484 12310 8536 12316
rect 8392 12300 8444 12306
rect 8392 12242 8444 12248
rect 8404 12209 8432 12242
rect 8390 12200 8446 12209
rect 8390 12135 8446 12144
rect 8496 11694 8524 12310
rect 8576 12300 8628 12306
rect 8576 12242 8628 12248
rect 8588 12102 8616 12242
rect 8772 12186 8800 12406
rect 8864 12306 8892 12582
rect 8852 12300 8904 12306
rect 8852 12242 8904 12248
rect 8772 12158 8892 12186
rect 8864 12102 8892 12158
rect 8576 12096 8628 12102
rect 8576 12038 8628 12044
rect 8760 12096 8812 12102
rect 8760 12038 8812 12044
rect 8852 12096 8904 12102
rect 8852 12038 8904 12044
rect 8484 11688 8536 11694
rect 8484 11630 8536 11636
rect 8298 11248 8354 11257
rect 8588 11218 8616 12038
rect 8772 11830 8800 12038
rect 8760 11824 8812 11830
rect 8680 11784 8760 11812
rect 8680 11218 8708 11784
rect 8760 11766 8812 11772
rect 8864 11762 8892 12038
rect 8852 11756 8904 11762
rect 8852 11698 8904 11704
rect 8760 11688 8812 11694
rect 8760 11630 8812 11636
rect 8772 11354 8800 11630
rect 8760 11348 8812 11354
rect 8760 11290 8812 11296
rect 8298 11183 8354 11192
rect 8576 11212 8628 11218
rect 8312 10742 8340 11183
rect 8576 11154 8628 11160
rect 8668 11212 8720 11218
rect 8668 11154 8720 11160
rect 8392 11144 8444 11150
rect 8392 11086 8444 11092
rect 8300 10736 8352 10742
rect 8206 10704 8262 10713
rect 8300 10678 8352 10684
rect 8206 10639 8262 10648
rect 8220 10554 8248 10639
rect 8220 10526 8340 10554
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 8220 10130 8248 10406
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 8206 10024 8262 10033
rect 8312 10010 8340 10526
rect 8404 10198 8432 11086
rect 8668 11076 8720 11082
rect 8668 11018 8720 11024
rect 8484 11008 8536 11014
rect 8484 10950 8536 10956
rect 8496 10266 8524 10950
rect 8680 10606 8708 11018
rect 8668 10600 8720 10606
rect 8668 10542 8720 10548
rect 8758 10568 8814 10577
rect 8758 10503 8814 10512
rect 8484 10260 8536 10266
rect 8772 10248 8800 10503
rect 8484 10202 8536 10208
rect 8680 10220 8800 10248
rect 8392 10192 8444 10198
rect 8392 10134 8444 10140
rect 8262 9982 8340 10010
rect 8206 9959 8262 9968
rect 8220 9586 8248 9959
rect 8496 9738 8524 10202
rect 8576 9920 8628 9926
rect 8576 9862 8628 9868
rect 8312 9722 8524 9738
rect 8300 9716 8524 9722
rect 8352 9710 8524 9716
rect 8300 9658 8352 9664
rect 8392 9648 8444 9654
rect 8392 9590 8444 9596
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 8208 9376 8260 9382
rect 8208 9318 8260 9324
rect 8116 9172 8168 9178
rect 8116 9114 8168 9120
rect 8116 8968 8168 8974
rect 8114 8936 8116 8945
rect 8168 8936 8170 8945
rect 8114 8871 8170 8880
rect 8128 7274 8156 8871
rect 8220 7834 8248 9318
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 8312 9042 8340 9114
rect 8300 9036 8352 9042
rect 8300 8978 8352 8984
rect 8312 8430 8340 8978
rect 8404 8498 8432 9590
rect 8484 9580 8536 9586
rect 8484 9522 8536 9528
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8300 8424 8352 8430
rect 8300 8366 8352 8372
rect 8390 7984 8446 7993
rect 8390 7919 8446 7928
rect 8220 7806 8340 7834
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 8116 7268 8168 7274
rect 8116 7210 8168 7216
rect 8116 6860 8168 6866
rect 8116 6802 8168 6808
rect 8128 6225 8156 6802
rect 8114 6216 8170 6225
rect 8114 6151 8170 6160
rect 8128 5846 8156 6151
rect 8116 5840 8168 5846
rect 8116 5782 8168 5788
rect 8220 5778 8248 7686
rect 8312 6390 8340 7806
rect 8404 7546 8432 7919
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 8390 7440 8446 7449
rect 8390 7375 8446 7384
rect 8404 7342 8432 7375
rect 8392 7336 8444 7342
rect 8392 7278 8444 7284
rect 8404 6662 8432 7278
rect 8392 6656 8444 6662
rect 8496 6633 8524 9522
rect 8588 9518 8616 9862
rect 8680 9586 8708 10220
rect 8760 10124 8812 10130
rect 8760 10066 8812 10072
rect 8772 9722 8800 10066
rect 8760 9716 8812 9722
rect 8760 9658 8812 9664
rect 8852 9716 8904 9722
rect 8852 9658 8904 9664
rect 8668 9580 8720 9586
rect 8668 9522 8720 9528
rect 8576 9512 8628 9518
rect 8576 9454 8628 9460
rect 8668 9444 8720 9450
rect 8668 9386 8720 9392
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 8588 8430 8616 8774
rect 8680 8537 8708 9386
rect 8760 9376 8812 9382
rect 8760 9318 8812 9324
rect 8666 8528 8722 8537
rect 8666 8463 8722 8472
rect 8576 8424 8628 8430
rect 8576 8366 8628 8372
rect 8680 6780 8708 8463
rect 8772 6798 8800 9318
rect 8864 8090 8892 9658
rect 8956 9586 8984 13495
rect 9048 13326 9076 13824
rect 9036 13320 9088 13326
rect 9036 13262 9088 13268
rect 9036 12164 9088 12170
rect 9036 12106 9088 12112
rect 9048 10305 9076 12106
rect 9140 10849 9168 14826
rect 9218 14784 9274 14793
rect 9218 14719 9274 14728
rect 9232 14618 9260 14719
rect 9220 14612 9272 14618
rect 9220 14554 9272 14560
rect 9324 14550 9352 14962
rect 9312 14544 9364 14550
rect 9312 14486 9364 14492
rect 9416 14482 9444 15302
rect 9220 14476 9272 14482
rect 9220 14418 9272 14424
rect 9404 14476 9456 14482
rect 9404 14418 9456 14424
rect 9232 13734 9260 14418
rect 9404 13864 9456 13870
rect 9404 13806 9456 13812
rect 9312 13796 9364 13802
rect 9312 13738 9364 13744
rect 9220 13728 9272 13734
rect 9220 13670 9272 13676
rect 9324 13462 9352 13738
rect 9312 13456 9364 13462
rect 9312 13398 9364 13404
rect 9220 13388 9272 13394
rect 9220 13330 9272 13336
rect 9232 12986 9260 13330
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 9220 12232 9272 12238
rect 9218 12200 9220 12209
rect 9272 12200 9274 12209
rect 9218 12135 9274 12144
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9126 10840 9182 10849
rect 9126 10775 9182 10784
rect 9034 10296 9090 10305
rect 9034 10231 9090 10240
rect 9036 10124 9088 10130
rect 9036 10066 9088 10072
rect 9220 10124 9272 10130
rect 9220 10066 9272 10072
rect 8944 9580 8996 9586
rect 8944 9522 8996 9528
rect 9048 9450 9076 10066
rect 9232 10033 9260 10066
rect 9218 10024 9274 10033
rect 9218 9959 9274 9968
rect 9128 9920 9180 9926
rect 9128 9862 9180 9868
rect 9140 9761 9168 9862
rect 9126 9752 9182 9761
rect 9126 9687 9182 9696
rect 9324 9625 9352 11290
rect 9416 10606 9444 13806
rect 9508 13705 9536 15422
rect 9588 15428 9640 15434
rect 9588 15370 9640 15376
rect 9600 14657 9628 15370
rect 9586 14648 9642 14657
rect 9586 14583 9642 14592
rect 9770 14512 9826 14521
rect 9588 14476 9640 14482
rect 9588 14418 9640 14424
rect 9680 14476 9732 14482
rect 9770 14447 9826 14456
rect 9680 14418 9732 14424
rect 9494 13696 9550 13705
rect 9494 13631 9550 13640
rect 9496 13388 9548 13394
rect 9600 13376 9628 14418
rect 9692 13530 9720 14418
rect 9784 14278 9812 14447
rect 9772 14272 9824 14278
rect 9772 14214 9824 14220
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 9784 13802 9812 14010
rect 9772 13796 9824 13802
rect 9772 13738 9824 13744
rect 9680 13524 9732 13530
rect 9680 13466 9732 13472
rect 9680 13388 9732 13394
rect 9600 13348 9680 13376
rect 9496 13330 9548 13336
rect 9680 13330 9732 13336
rect 9404 10600 9456 10606
rect 9404 10542 9456 10548
rect 9404 10124 9456 10130
rect 9404 10066 9456 10072
rect 9416 9926 9444 10066
rect 9404 9920 9456 9926
rect 9404 9862 9456 9868
rect 9416 9722 9444 9862
rect 9404 9716 9456 9722
rect 9404 9658 9456 9664
rect 9310 9616 9366 9625
rect 9310 9551 9366 9560
rect 9404 9580 9456 9586
rect 9036 9444 9088 9450
rect 9036 9386 9088 9392
rect 8944 8900 8996 8906
rect 8944 8842 8996 8848
rect 8956 8634 8984 8842
rect 8944 8628 8996 8634
rect 8944 8570 8996 8576
rect 8956 8498 8984 8570
rect 8944 8492 8996 8498
rect 8944 8434 8996 8440
rect 8944 8288 8996 8294
rect 8944 8230 8996 8236
rect 8852 8084 8904 8090
rect 8852 8026 8904 8032
rect 8864 6934 8892 8026
rect 8956 7993 8984 8230
rect 9048 8090 9076 9386
rect 9324 8922 9352 9551
rect 9404 9522 9456 9528
rect 9140 8894 9352 8922
rect 9036 8084 9088 8090
rect 9036 8026 9088 8032
rect 8942 7984 8998 7993
rect 9140 7936 9168 8894
rect 9416 8566 9444 9522
rect 9508 9500 9536 13330
rect 9772 13252 9824 13258
rect 9772 13194 9824 13200
rect 9784 13025 9812 13194
rect 9770 13016 9826 13025
rect 9770 12951 9826 12960
rect 9770 12880 9826 12889
rect 9770 12815 9826 12824
rect 9680 12776 9732 12782
rect 9680 12718 9732 12724
rect 9692 12442 9720 12718
rect 9784 12646 9812 12815
rect 9772 12640 9824 12646
rect 9772 12582 9824 12588
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9588 11552 9640 11558
rect 9588 11494 9640 11500
rect 9600 9926 9628 11494
rect 9692 11218 9720 12378
rect 9772 12096 9824 12102
rect 9772 12038 9824 12044
rect 9784 11898 9812 12038
rect 9876 11898 9904 15864
rect 9956 15632 10008 15638
rect 9956 15574 10008 15580
rect 9968 14414 9996 15574
rect 10060 15570 10088 15982
rect 10140 15972 10192 15978
rect 10140 15914 10192 15920
rect 10048 15564 10100 15570
rect 10048 15506 10100 15512
rect 10152 15502 10180 15914
rect 10140 15496 10192 15502
rect 10140 15438 10192 15444
rect 10244 15434 10272 15982
rect 10364 15804 10740 15813
rect 10420 15802 10444 15804
rect 10500 15802 10524 15804
rect 10580 15802 10604 15804
rect 10660 15802 10684 15804
rect 10420 15750 10430 15802
rect 10674 15750 10684 15802
rect 10420 15748 10444 15750
rect 10500 15748 10524 15750
rect 10580 15748 10604 15750
rect 10660 15748 10684 15750
rect 10364 15739 10740 15748
rect 10324 15564 10376 15570
rect 10324 15506 10376 15512
rect 10232 15428 10284 15434
rect 10232 15370 10284 15376
rect 10336 15162 10364 15506
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 10692 15496 10744 15502
rect 10692 15438 10744 15444
rect 10324 15156 10376 15162
rect 10324 15098 10376 15104
rect 10232 15088 10284 15094
rect 10046 15056 10102 15065
rect 10232 15030 10284 15036
rect 10046 14991 10102 15000
rect 10060 14618 10088 14991
rect 10140 14952 10192 14958
rect 10140 14894 10192 14900
rect 10152 14657 10180 14894
rect 10138 14648 10194 14657
rect 10048 14612 10100 14618
rect 10138 14583 10194 14592
rect 10048 14554 10100 14560
rect 10048 14476 10100 14482
rect 10048 14418 10100 14424
rect 9956 14408 10008 14414
rect 9956 14350 10008 14356
rect 9956 14272 10008 14278
rect 9956 14214 10008 14220
rect 9772 11892 9824 11898
rect 9772 11834 9824 11840
rect 9864 11892 9916 11898
rect 9864 11834 9916 11840
rect 9876 11694 9904 11834
rect 9864 11688 9916 11694
rect 9864 11630 9916 11636
rect 9680 11212 9732 11218
rect 9680 11154 9732 11160
rect 9968 10554 9996 14214
rect 10060 13734 10088 14418
rect 10138 14376 10194 14385
rect 10138 14311 10140 14320
rect 10192 14311 10194 14320
rect 10244 14328 10272 15030
rect 10428 14822 10456 15438
rect 10598 15056 10654 15065
rect 10704 15026 10732 15438
rect 10598 14991 10654 15000
rect 10692 15020 10744 15026
rect 10612 14958 10640 14991
rect 10692 14962 10744 14968
rect 10600 14952 10652 14958
rect 10600 14894 10652 14900
rect 10416 14816 10468 14822
rect 10416 14758 10468 14764
rect 10364 14716 10740 14725
rect 10420 14714 10444 14716
rect 10500 14714 10524 14716
rect 10580 14714 10604 14716
rect 10660 14714 10684 14716
rect 10420 14662 10430 14714
rect 10674 14662 10684 14714
rect 10420 14660 10444 14662
rect 10500 14660 10524 14662
rect 10580 14660 10604 14662
rect 10660 14660 10684 14662
rect 10364 14651 10740 14660
rect 10600 14544 10652 14550
rect 10600 14486 10652 14492
rect 10416 14408 10468 14414
rect 10416 14350 10468 14356
rect 10324 14340 10376 14346
rect 10140 14282 10192 14288
rect 10244 14300 10324 14328
rect 10138 14104 10194 14113
rect 10138 14039 10194 14048
rect 10048 13728 10100 13734
rect 10048 13670 10100 13676
rect 10152 13462 10180 14039
rect 10244 13870 10272 14300
rect 10324 14282 10376 14288
rect 10428 14074 10456 14350
rect 10508 14272 10560 14278
rect 10508 14214 10560 14220
rect 10416 14068 10468 14074
rect 10416 14010 10468 14016
rect 10232 13864 10284 13870
rect 10232 13806 10284 13812
rect 10322 13832 10378 13841
rect 10322 13767 10378 13776
rect 10336 13734 10364 13767
rect 10520 13734 10548 14214
rect 10612 13802 10640 14486
rect 10796 14278 10824 16102
rect 10980 15570 11008 16390
rect 10968 15564 11020 15570
rect 10968 15506 11020 15512
rect 10876 15428 10928 15434
rect 10876 15370 10928 15376
rect 10784 14272 10836 14278
rect 10690 14240 10746 14249
rect 10784 14214 10836 14220
rect 10690 14175 10746 14184
rect 10704 14006 10732 14175
rect 10692 14000 10744 14006
rect 10692 13942 10744 13948
rect 10600 13796 10652 13802
rect 10600 13738 10652 13744
rect 10232 13728 10284 13734
rect 10232 13670 10284 13676
rect 10324 13728 10376 13734
rect 10324 13670 10376 13676
rect 10508 13728 10560 13734
rect 10508 13670 10560 13676
rect 10244 13530 10272 13670
rect 10364 13628 10740 13637
rect 10420 13626 10444 13628
rect 10500 13626 10524 13628
rect 10580 13626 10604 13628
rect 10660 13626 10684 13628
rect 10420 13574 10430 13626
rect 10674 13574 10684 13626
rect 10420 13572 10444 13574
rect 10500 13572 10524 13574
rect 10580 13572 10604 13574
rect 10660 13572 10684 13574
rect 10364 13563 10740 13572
rect 10232 13524 10284 13530
rect 10888 13512 10916 15370
rect 10966 15192 11022 15201
rect 10966 15127 11022 15136
rect 10980 14958 11008 15127
rect 10968 14952 11020 14958
rect 10968 14894 11020 14900
rect 11060 14952 11112 14958
rect 11060 14894 11112 14900
rect 10968 14816 11020 14822
rect 10968 14758 11020 14764
rect 10980 14482 11008 14758
rect 11072 14618 11100 14894
rect 11060 14612 11112 14618
rect 11060 14554 11112 14560
rect 10968 14476 11020 14482
rect 10968 14418 11020 14424
rect 10232 13466 10284 13472
rect 10796 13484 10916 13512
rect 10140 13456 10192 13462
rect 10140 13398 10192 13404
rect 10140 13184 10192 13190
rect 10140 13126 10192 13132
rect 10048 12912 10100 12918
rect 10048 12854 10100 12860
rect 9876 10526 9996 10554
rect 9876 10010 9904 10526
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 9968 10130 9996 10406
rect 9956 10124 10008 10130
rect 9956 10066 10008 10072
rect 9876 9982 9996 10010
rect 9588 9920 9640 9926
rect 9588 9862 9640 9868
rect 9862 9752 9918 9761
rect 9862 9687 9918 9696
rect 9680 9512 9732 9518
rect 9508 9489 9680 9500
rect 9494 9480 9680 9489
rect 9550 9472 9680 9480
rect 9680 9454 9732 9460
rect 9494 9415 9550 9424
rect 9772 9036 9824 9042
rect 9772 8978 9824 8984
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 9586 8664 9642 8673
rect 9496 8628 9548 8634
rect 9586 8599 9588 8608
rect 9496 8570 9548 8576
rect 9640 8599 9642 8608
rect 9588 8570 9640 8576
rect 9404 8560 9456 8566
rect 9404 8502 9456 8508
rect 9220 8356 9272 8362
rect 9220 8298 9272 8304
rect 9232 8090 9260 8298
rect 9310 8256 9366 8265
rect 9310 8191 9366 8200
rect 9220 8084 9272 8090
rect 9220 8026 9272 8032
rect 8942 7919 8998 7928
rect 9048 7908 9168 7936
rect 9220 7948 9272 7954
rect 8944 7880 8996 7886
rect 8944 7822 8996 7828
rect 8852 6928 8904 6934
rect 8852 6870 8904 6876
rect 8588 6752 8708 6780
rect 8760 6792 8812 6798
rect 8392 6598 8444 6604
rect 8482 6624 8538 6633
rect 8300 6384 8352 6390
rect 8300 6326 8352 6332
rect 8404 6254 8432 6598
rect 8482 6559 8538 6568
rect 8588 6254 8616 6752
rect 8956 6780 8984 7822
rect 9048 6866 9076 7908
rect 9220 7890 9272 7896
rect 9126 7848 9182 7857
rect 9126 7783 9128 7792
rect 9180 7783 9182 7792
rect 9128 7754 9180 7760
rect 9140 7478 9168 7754
rect 9128 7472 9180 7478
rect 9128 7414 9180 7420
rect 9232 7342 9260 7890
rect 9220 7336 9272 7342
rect 9220 7278 9272 7284
rect 9128 7200 9180 7206
rect 9128 7142 9180 7148
rect 9036 6860 9088 6866
rect 9036 6802 9088 6808
rect 8760 6734 8812 6740
rect 8864 6752 8984 6780
rect 8668 6656 8720 6662
rect 8864 6644 8892 6752
rect 8668 6598 8720 6604
rect 8772 6616 8892 6644
rect 9034 6624 9090 6633
rect 8680 6254 8708 6598
rect 8392 6248 8444 6254
rect 8392 6190 8444 6196
rect 8576 6248 8628 6254
rect 8576 6190 8628 6196
rect 8668 6248 8720 6254
rect 8668 6190 8720 6196
rect 8392 6112 8444 6118
rect 8392 6054 8444 6060
rect 8208 5772 8260 5778
rect 8208 5714 8260 5720
rect 8116 5704 8168 5710
rect 8114 5672 8116 5681
rect 8168 5672 8170 5681
rect 8114 5607 8170 5616
rect 8114 5536 8170 5545
rect 8114 5471 8170 5480
rect 8128 5098 8156 5471
rect 8116 5092 8168 5098
rect 8116 5034 8168 5040
rect 8404 4690 8432 6054
rect 8484 5772 8536 5778
rect 8484 5714 8536 5720
rect 8496 5370 8524 5714
rect 8668 5704 8720 5710
rect 8668 5646 8720 5652
rect 8576 5568 8628 5574
rect 8576 5510 8628 5516
rect 8484 5364 8536 5370
rect 8484 5306 8536 5312
rect 8588 5234 8616 5510
rect 8576 5228 8628 5234
rect 8576 5170 8628 5176
rect 8392 4684 8444 4690
rect 8392 4626 8444 4632
rect 8576 4684 8628 4690
rect 8680 4672 8708 5646
rect 8772 5166 8800 6616
rect 9034 6559 9090 6568
rect 8852 6452 8904 6458
rect 8852 6394 8904 6400
rect 8864 6254 8892 6394
rect 9048 6254 9076 6559
rect 8852 6248 8904 6254
rect 8852 6190 8904 6196
rect 9036 6248 9088 6254
rect 9036 6190 9088 6196
rect 8852 5908 8904 5914
rect 8852 5850 8904 5856
rect 8864 5658 8892 5850
rect 8864 5630 9076 5658
rect 8852 5568 8904 5574
rect 8852 5510 8904 5516
rect 8944 5568 8996 5574
rect 8944 5510 8996 5516
rect 8760 5160 8812 5166
rect 8760 5102 8812 5108
rect 8628 4644 8708 4672
rect 8576 4626 8628 4632
rect 8116 4616 8168 4622
rect 8116 4558 8168 4564
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 8024 4276 8076 4282
rect 8024 4218 8076 4224
rect 8022 4176 8078 4185
rect 8128 4146 8156 4558
rect 8022 4111 8078 4120
rect 8116 4140 8168 4146
rect 7932 3732 7984 3738
rect 7932 3674 7984 3680
rect 7840 3664 7892 3670
rect 7840 3606 7892 3612
rect 7288 3596 7340 3602
rect 7288 3538 7340 3544
rect 6736 3188 6788 3194
rect 6736 3130 6788 3136
rect 7196 3188 7248 3194
rect 7196 3130 7248 3136
rect 6552 2644 6604 2650
rect 6552 2586 6604 2592
rect 6748 2514 6776 3130
rect 6828 3052 6880 3058
rect 6828 2994 6880 3000
rect 6840 2582 6868 2994
rect 7300 2990 7328 3538
rect 7364 3292 7740 3301
rect 7420 3290 7444 3292
rect 7500 3290 7524 3292
rect 7580 3290 7604 3292
rect 7660 3290 7684 3292
rect 7420 3238 7430 3290
rect 7674 3238 7684 3290
rect 7420 3236 7444 3238
rect 7500 3236 7524 3238
rect 7580 3236 7604 3238
rect 7660 3236 7684 3238
rect 7364 3227 7740 3236
rect 7746 3088 7802 3097
rect 7852 3074 7880 3606
rect 7802 3046 7880 3074
rect 7746 3023 7802 3032
rect 7288 2984 7340 2990
rect 7288 2926 7340 2932
rect 7472 2984 7524 2990
rect 7472 2926 7524 2932
rect 7288 2848 7340 2854
rect 7288 2790 7340 2796
rect 6828 2576 6880 2582
rect 6828 2518 6880 2524
rect 6736 2508 6788 2514
rect 6736 2450 6788 2456
rect 6644 2032 6696 2038
rect 6642 2000 6644 2009
rect 6696 2000 6698 2009
rect 6748 1970 6776 2450
rect 7012 2440 7064 2446
rect 7012 2382 7064 2388
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 6642 1935 6698 1944
rect 6736 1964 6788 1970
rect 6656 1562 6684 1935
rect 6736 1906 6788 1912
rect 7024 1902 7052 2382
rect 7116 1902 7144 2382
rect 7300 2106 7328 2790
rect 7484 2650 7512 2926
rect 7472 2644 7524 2650
rect 7472 2586 7524 2592
rect 7760 2514 7788 3023
rect 7748 2508 7800 2514
rect 7748 2450 7800 2456
rect 7840 2304 7892 2310
rect 7840 2246 7892 2252
rect 7364 2204 7740 2213
rect 7420 2202 7444 2204
rect 7500 2202 7524 2204
rect 7580 2202 7604 2204
rect 7660 2202 7684 2204
rect 7420 2150 7430 2202
rect 7674 2150 7684 2202
rect 7420 2148 7444 2150
rect 7500 2148 7524 2150
rect 7580 2148 7604 2150
rect 7660 2148 7684 2150
rect 7364 2139 7740 2148
rect 7288 2100 7340 2106
rect 7288 2042 7340 2048
rect 7012 1896 7064 1902
rect 7012 1838 7064 1844
rect 7104 1896 7156 1902
rect 7104 1838 7156 1844
rect 6644 1556 6696 1562
rect 6644 1498 6696 1504
rect 6734 1456 6790 1465
rect 6734 1391 6736 1400
rect 6788 1391 6790 1400
rect 6736 1362 6788 1368
rect 6368 1284 6420 1290
rect 6368 1226 6420 1232
rect 6184 1216 6236 1222
rect 6184 1158 6236 1164
rect 6000 1012 6052 1018
rect 6000 954 6052 960
rect 6092 1012 6144 1018
rect 6092 954 6144 960
rect 6104 898 6132 954
rect 5920 870 6132 898
rect 5920 814 5948 870
rect 6196 814 6224 1158
rect 5908 808 5960 814
rect 5262 776 5318 785
rect 5908 750 5960 756
rect 6184 808 6236 814
rect 6184 750 6236 756
rect 6748 746 6776 1362
rect 7116 1358 7144 1838
rect 7852 1426 7880 2246
rect 7932 1760 7984 1766
rect 7932 1702 7984 1708
rect 7944 1426 7972 1702
rect 7840 1420 7892 1426
rect 7840 1362 7892 1368
rect 7932 1420 7984 1426
rect 7932 1362 7984 1368
rect 6828 1352 6880 1358
rect 6828 1294 6880 1300
rect 7104 1352 7156 1358
rect 7104 1294 7156 1300
rect 6840 1018 6868 1294
rect 7364 1116 7740 1125
rect 7420 1114 7444 1116
rect 7500 1114 7524 1116
rect 7580 1114 7604 1116
rect 7660 1114 7684 1116
rect 7420 1062 7430 1114
rect 7674 1062 7684 1114
rect 7420 1060 7444 1062
rect 7500 1060 7524 1062
rect 7580 1060 7604 1062
rect 7660 1060 7684 1062
rect 7364 1051 7740 1060
rect 7852 1018 7880 1362
rect 6828 1012 6880 1018
rect 6828 954 6880 960
rect 7840 1012 7892 1018
rect 7840 954 7892 960
rect 7104 944 7156 950
rect 7102 912 7104 921
rect 7156 912 7158 921
rect 7944 882 7972 1362
rect 8036 1290 8064 4111
rect 8116 4082 8168 4088
rect 8312 3602 8340 4558
rect 8392 4548 8444 4554
rect 8392 4490 8444 4496
rect 8404 4282 8432 4490
rect 8392 4276 8444 4282
rect 8392 4218 8444 4224
rect 8588 4078 8616 4626
rect 8668 4480 8720 4486
rect 8668 4422 8720 4428
rect 8576 4072 8628 4078
rect 8576 4014 8628 4020
rect 8300 3596 8352 3602
rect 8300 3538 8352 3544
rect 8300 3392 8352 3398
rect 8300 3334 8352 3340
rect 8312 3058 8340 3334
rect 8680 3194 8708 4422
rect 8864 3738 8892 5510
rect 8956 5302 8984 5510
rect 8944 5296 8996 5302
rect 8944 5238 8996 5244
rect 8944 4480 8996 4486
rect 8944 4422 8996 4428
rect 8956 4146 8984 4422
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 8944 4004 8996 4010
rect 8944 3946 8996 3952
rect 8852 3732 8904 3738
rect 8852 3674 8904 3680
rect 8956 3602 8984 3946
rect 9048 3641 9076 5630
rect 9140 5234 9168 7142
rect 9324 6984 9352 8191
rect 9416 7954 9444 8502
rect 9508 8412 9536 8570
rect 9692 8430 9720 8774
rect 9588 8424 9640 8430
rect 9508 8384 9588 8412
rect 9588 8366 9640 8372
rect 9680 8424 9732 8430
rect 9784 8401 9812 8978
rect 9876 8566 9904 9687
rect 9864 8560 9916 8566
rect 9864 8502 9916 8508
rect 9680 8366 9732 8372
rect 9770 8392 9826 8401
rect 9770 8327 9826 8336
rect 9496 8288 9548 8294
rect 9548 8248 9674 8276
rect 9496 8230 9548 8236
rect 9646 8072 9674 8248
rect 9508 8044 9674 8072
rect 9404 7948 9456 7954
rect 9404 7890 9456 7896
rect 9508 7886 9536 8044
rect 9586 7984 9642 7993
rect 9784 7954 9812 8327
rect 9864 8288 9916 8294
rect 9864 8230 9916 8236
rect 9586 7919 9642 7928
rect 9772 7948 9824 7954
rect 9496 7880 9548 7886
rect 9496 7822 9548 7828
rect 9600 7818 9628 7919
rect 9772 7890 9824 7896
rect 9588 7812 9640 7818
rect 9588 7754 9640 7760
rect 9404 7744 9456 7750
rect 9404 7686 9456 7692
rect 9680 7744 9732 7750
rect 9680 7686 9732 7692
rect 9232 6956 9352 6984
rect 9232 6458 9260 6956
rect 9312 6860 9364 6866
rect 9312 6802 9364 6808
rect 9220 6452 9272 6458
rect 9220 6394 9272 6400
rect 9218 6352 9274 6361
rect 9324 6322 9352 6802
rect 9218 6287 9274 6296
rect 9312 6316 9364 6322
rect 9232 6254 9260 6287
rect 9312 6258 9364 6264
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 9128 5228 9180 5234
rect 9128 5170 9180 5176
rect 9140 4146 9168 5170
rect 9220 5160 9272 5166
rect 9220 5102 9272 5108
rect 9232 4826 9260 5102
rect 9324 5098 9352 6258
rect 9416 5778 9444 7686
rect 9692 7410 9720 7686
rect 9680 7404 9732 7410
rect 9680 7346 9732 7352
rect 9772 7404 9824 7410
rect 9772 7346 9824 7352
rect 9678 7304 9734 7313
rect 9678 7239 9734 7248
rect 9588 6860 9640 6866
rect 9588 6802 9640 6808
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9404 5772 9456 5778
rect 9404 5714 9456 5720
rect 9312 5092 9364 5098
rect 9312 5034 9364 5040
rect 9220 4820 9272 4826
rect 9220 4762 9272 4768
rect 9416 4214 9444 5714
rect 9404 4208 9456 4214
rect 9404 4150 9456 4156
rect 9128 4140 9180 4146
rect 9128 4082 9180 4088
rect 9312 4072 9364 4078
rect 9312 4014 9364 4020
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 9034 3632 9090 3641
rect 8760 3596 8812 3602
rect 8760 3538 8812 3544
rect 8944 3596 8996 3602
rect 9034 3567 9090 3576
rect 8944 3538 8996 3544
rect 8772 3482 8800 3538
rect 8772 3454 8892 3482
rect 8864 3398 8892 3454
rect 8760 3392 8812 3398
rect 8760 3334 8812 3340
rect 8852 3392 8904 3398
rect 8852 3334 8904 3340
rect 8668 3188 8720 3194
rect 8668 3130 8720 3136
rect 8300 3052 8352 3058
rect 8300 2994 8352 3000
rect 8484 2848 8536 2854
rect 8484 2790 8536 2796
rect 8496 2514 8524 2790
rect 8772 2514 8800 3334
rect 9232 3126 9260 3878
rect 9324 3618 9352 4014
rect 9324 3602 9444 3618
rect 9508 3602 9536 6598
rect 9600 6458 9628 6802
rect 9588 6452 9640 6458
rect 9588 6394 9640 6400
rect 9586 6352 9642 6361
rect 9586 6287 9642 6296
rect 9600 6254 9628 6287
rect 9588 6248 9640 6254
rect 9588 6190 9640 6196
rect 9692 4434 9720 7239
rect 9784 6866 9812 7346
rect 9876 7002 9904 8230
rect 9864 6996 9916 7002
rect 9864 6938 9916 6944
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9772 5636 9824 5642
rect 9772 5578 9824 5584
rect 9784 5030 9812 5578
rect 9772 5024 9824 5030
rect 9772 4966 9824 4972
rect 9784 4758 9812 4966
rect 9772 4752 9824 4758
rect 9772 4694 9824 4700
rect 9772 4480 9824 4486
rect 9692 4428 9772 4434
rect 9692 4422 9824 4428
rect 9692 4406 9812 4422
rect 9680 4276 9732 4282
rect 9680 4218 9732 4224
rect 9588 4208 9640 4214
rect 9588 4150 9640 4156
rect 9600 4010 9628 4150
rect 9692 4078 9720 4218
rect 9772 4208 9824 4214
rect 9772 4150 9824 4156
rect 9680 4072 9732 4078
rect 9680 4014 9732 4020
rect 9588 4004 9640 4010
rect 9588 3946 9640 3952
rect 9680 3936 9732 3942
rect 9680 3878 9732 3884
rect 9588 3732 9640 3738
rect 9588 3674 9640 3680
rect 9312 3596 9444 3602
rect 9364 3590 9444 3596
rect 9312 3538 9364 3544
rect 9312 3460 9364 3466
rect 9312 3402 9364 3408
rect 9220 3120 9272 3126
rect 9220 3062 9272 3068
rect 9324 3058 9352 3402
rect 9416 3194 9444 3590
rect 9496 3596 9548 3602
rect 9496 3538 9548 3544
rect 9496 3460 9548 3466
rect 9496 3402 9548 3408
rect 9404 3188 9456 3194
rect 9404 3130 9456 3136
rect 9312 3052 9364 3058
rect 9312 2994 9364 3000
rect 9128 2848 9180 2854
rect 9128 2790 9180 2796
rect 9140 2582 9168 2790
rect 9128 2576 9180 2582
rect 9128 2518 9180 2524
rect 9508 2514 9536 3402
rect 9600 3126 9628 3674
rect 9692 3670 9720 3878
rect 9784 3670 9812 4150
rect 9680 3664 9732 3670
rect 9680 3606 9732 3612
rect 9772 3664 9824 3670
rect 9772 3606 9824 3612
rect 9588 3120 9640 3126
rect 9588 3062 9640 3068
rect 9588 2984 9640 2990
rect 9586 2952 9588 2961
rect 9640 2952 9642 2961
rect 9586 2887 9642 2896
rect 9692 2582 9720 3606
rect 9772 3528 9824 3534
rect 9876 3516 9904 6938
rect 9968 5953 9996 9982
rect 10060 9897 10088 12854
rect 10152 11354 10180 13126
rect 10244 12782 10272 13466
rect 10508 13388 10560 13394
rect 10508 13330 10560 13336
rect 10520 12918 10548 13330
rect 10508 12912 10560 12918
rect 10508 12854 10560 12860
rect 10520 12782 10548 12854
rect 10232 12776 10284 12782
rect 10232 12718 10284 12724
rect 10508 12776 10560 12782
rect 10508 12718 10560 12724
rect 10364 12540 10740 12549
rect 10420 12538 10444 12540
rect 10500 12538 10524 12540
rect 10580 12538 10604 12540
rect 10660 12538 10684 12540
rect 10420 12486 10430 12538
rect 10674 12486 10684 12538
rect 10420 12484 10444 12486
rect 10500 12484 10524 12486
rect 10580 12484 10604 12486
rect 10660 12484 10684 12486
rect 10364 12475 10740 12484
rect 10796 12170 10824 13484
rect 10980 13444 11008 14418
rect 11060 14272 11112 14278
rect 11060 14214 11112 14220
rect 11072 14113 11100 14214
rect 11058 14104 11114 14113
rect 11058 14039 11114 14048
rect 10888 13416 11008 13444
rect 10888 12170 10916 13416
rect 11060 13388 11112 13394
rect 11060 13330 11112 13336
rect 10968 13320 11020 13326
rect 10968 13262 11020 13268
rect 10980 12986 11008 13262
rect 10968 12980 11020 12986
rect 10968 12922 11020 12928
rect 11072 12374 11100 13330
rect 11164 12434 11192 18108
rect 11256 17241 11284 18380
rect 11428 18352 11480 18358
rect 11428 18294 11480 18300
rect 11336 18284 11388 18290
rect 11336 18226 11388 18232
rect 11242 17232 11298 17241
rect 11242 17167 11298 17176
rect 11348 17066 11376 18226
rect 11440 17338 11468 18294
rect 11532 18193 11560 18634
rect 11704 18420 11756 18426
rect 11756 18380 11928 18408
rect 11704 18362 11756 18368
rect 11704 18216 11756 18222
rect 11518 18184 11574 18193
rect 11704 18158 11756 18164
rect 11518 18119 11574 18128
rect 11532 18086 11560 18119
rect 11520 18080 11572 18086
rect 11520 18022 11572 18028
rect 11716 17338 11744 18158
rect 11428 17332 11480 17338
rect 11428 17274 11480 17280
rect 11704 17332 11756 17338
rect 11704 17274 11756 17280
rect 11336 17060 11388 17066
rect 11256 17020 11336 17048
rect 11256 14090 11284 17020
rect 11336 17002 11388 17008
rect 11334 16688 11390 16697
rect 11334 16623 11336 16632
rect 11388 16623 11390 16632
rect 11336 16594 11388 16600
rect 11336 15904 11388 15910
rect 11336 15846 11388 15852
rect 11348 15502 11376 15846
rect 11336 15496 11388 15502
rect 11336 15438 11388 15444
rect 11440 14940 11468 17274
rect 11702 16688 11758 16697
rect 11702 16623 11758 16632
rect 11520 16448 11572 16454
rect 11520 16390 11572 16396
rect 11612 16448 11664 16454
rect 11612 16390 11664 16396
rect 11348 14912 11468 14940
rect 11348 14278 11376 14912
rect 11336 14272 11388 14278
rect 11336 14214 11388 14220
rect 11256 14062 11468 14090
rect 11244 14000 11296 14006
rect 11244 13942 11296 13948
rect 11256 13394 11284 13942
rect 11336 13796 11388 13802
rect 11336 13738 11388 13744
rect 11348 13530 11376 13738
rect 11336 13524 11388 13530
rect 11336 13466 11388 13472
rect 11244 13388 11296 13394
rect 11244 13330 11296 13336
rect 11336 12844 11388 12850
rect 11336 12786 11388 12792
rect 11164 12406 11284 12434
rect 11060 12368 11112 12374
rect 11060 12310 11112 12316
rect 10784 12164 10836 12170
rect 10784 12106 10836 12112
rect 10876 12164 10928 12170
rect 10876 12106 10928 12112
rect 10874 11928 10930 11937
rect 10874 11863 10930 11872
rect 10364 11452 10740 11461
rect 10420 11450 10444 11452
rect 10500 11450 10524 11452
rect 10580 11450 10604 11452
rect 10660 11450 10684 11452
rect 10420 11398 10430 11450
rect 10674 11398 10684 11450
rect 10420 11396 10444 11398
rect 10500 11396 10524 11398
rect 10580 11396 10604 11398
rect 10660 11396 10684 11398
rect 10364 11387 10740 11396
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 10784 11008 10836 11014
rect 10784 10950 10836 10956
rect 10232 10804 10284 10810
rect 10232 10746 10284 10752
rect 10140 10736 10192 10742
rect 10140 10678 10192 10684
rect 10152 10130 10180 10678
rect 10244 10606 10272 10746
rect 10232 10600 10284 10606
rect 10232 10542 10284 10548
rect 10324 10600 10376 10606
rect 10324 10542 10376 10548
rect 10336 10452 10364 10542
rect 10244 10424 10364 10452
rect 10140 10124 10192 10130
rect 10140 10066 10192 10072
rect 10140 9988 10192 9994
rect 10244 9976 10272 10424
rect 10364 10364 10740 10373
rect 10420 10362 10444 10364
rect 10500 10362 10524 10364
rect 10580 10362 10604 10364
rect 10660 10362 10684 10364
rect 10420 10310 10430 10362
rect 10674 10310 10684 10362
rect 10420 10308 10444 10310
rect 10500 10308 10524 10310
rect 10580 10308 10604 10310
rect 10660 10308 10684 10310
rect 10364 10299 10740 10308
rect 10508 10124 10560 10130
rect 10508 10066 10560 10072
rect 10192 9948 10272 9976
rect 10140 9930 10192 9936
rect 10046 9888 10102 9897
rect 10046 9823 10102 9832
rect 10152 9674 10180 9930
rect 10520 9926 10548 10066
rect 10508 9920 10560 9926
rect 10508 9862 10560 9868
rect 10060 9646 10180 9674
rect 10796 9654 10824 10950
rect 10888 10742 10916 11863
rect 11152 11688 11204 11694
rect 11152 11630 11204 11636
rect 10968 11552 11020 11558
rect 10968 11494 11020 11500
rect 11060 11552 11112 11558
rect 11060 11494 11112 11500
rect 10876 10736 10928 10742
rect 10876 10678 10928 10684
rect 10876 10600 10928 10606
rect 10876 10542 10928 10548
rect 10888 10470 10916 10542
rect 10876 10464 10928 10470
rect 10876 10406 10928 10412
rect 10980 10198 11008 11494
rect 11072 11218 11100 11494
rect 11164 11218 11192 11630
rect 11060 11212 11112 11218
rect 11060 11154 11112 11160
rect 11152 11212 11204 11218
rect 11152 11154 11204 11160
rect 11152 10532 11204 10538
rect 11152 10474 11204 10480
rect 11164 10266 11192 10474
rect 11152 10260 11204 10266
rect 11152 10202 11204 10208
rect 10968 10192 11020 10198
rect 10968 10134 11020 10140
rect 11058 9752 11114 9761
rect 11058 9687 11114 9696
rect 10784 9648 10836 9654
rect 10060 9450 10088 9646
rect 10784 9590 10836 9596
rect 10692 9512 10744 9518
rect 10322 9480 10378 9489
rect 10048 9444 10100 9450
rect 10048 9386 10100 9392
rect 10244 9438 10322 9466
rect 10796 9500 10824 9590
rect 11072 9518 11100 9687
rect 10744 9472 10824 9500
rect 10876 9512 10928 9518
rect 10692 9454 10744 9460
rect 11060 9512 11112 9518
rect 10928 9472 11008 9500
rect 10876 9454 10928 9460
rect 10048 8560 10100 8566
rect 10048 8502 10100 8508
rect 10060 7342 10088 8502
rect 10244 7936 10272 9438
rect 10322 9415 10324 9424
rect 10376 9415 10378 9424
rect 10324 9386 10376 9392
rect 10874 9344 10930 9353
rect 10364 9276 10740 9285
rect 10874 9279 10930 9288
rect 10420 9274 10444 9276
rect 10500 9274 10524 9276
rect 10580 9274 10604 9276
rect 10660 9274 10684 9276
rect 10420 9222 10430 9274
rect 10674 9222 10684 9274
rect 10420 9220 10444 9222
rect 10500 9220 10524 9222
rect 10580 9220 10604 9222
rect 10660 9220 10684 9222
rect 10364 9211 10740 9220
rect 10416 8968 10468 8974
rect 10416 8910 10468 8916
rect 10428 8430 10456 8910
rect 10888 8906 10916 9279
rect 10876 8900 10928 8906
rect 10876 8842 10928 8848
rect 10324 8424 10376 8430
rect 10322 8392 10324 8401
rect 10416 8424 10468 8430
rect 10376 8392 10378 8401
rect 10416 8366 10468 8372
rect 10876 8424 10928 8430
rect 10876 8366 10928 8372
rect 10322 8327 10378 8336
rect 10364 8188 10740 8197
rect 10420 8186 10444 8188
rect 10500 8186 10524 8188
rect 10580 8186 10604 8188
rect 10660 8186 10684 8188
rect 10420 8134 10430 8186
rect 10674 8134 10684 8186
rect 10420 8132 10444 8134
rect 10500 8132 10524 8134
rect 10580 8132 10604 8134
rect 10660 8132 10684 8134
rect 10364 8123 10740 8132
rect 10508 8084 10560 8090
rect 10508 8026 10560 8032
rect 10520 7954 10548 8026
rect 10782 7984 10838 7993
rect 10324 7948 10376 7954
rect 10244 7908 10324 7936
rect 10048 7336 10100 7342
rect 10048 7278 10100 7284
rect 10060 6089 10088 7278
rect 10140 7268 10192 7274
rect 10140 7210 10192 7216
rect 10046 6080 10102 6089
rect 10046 6015 10102 6024
rect 9954 5944 10010 5953
rect 9954 5879 10010 5888
rect 9956 5772 10008 5778
rect 9956 5714 10008 5720
rect 9968 5370 9996 5714
rect 10152 5574 10180 7210
rect 10244 7002 10272 7908
rect 10324 7890 10376 7896
rect 10508 7948 10560 7954
rect 10782 7919 10838 7928
rect 10508 7890 10560 7896
rect 10520 7546 10548 7890
rect 10508 7540 10560 7546
rect 10508 7482 10560 7488
rect 10364 7100 10740 7109
rect 10420 7098 10444 7100
rect 10500 7098 10524 7100
rect 10580 7098 10604 7100
rect 10660 7098 10684 7100
rect 10420 7046 10430 7098
rect 10674 7046 10684 7098
rect 10420 7044 10444 7046
rect 10500 7044 10524 7046
rect 10580 7044 10604 7046
rect 10660 7044 10684 7046
rect 10364 7035 10740 7044
rect 10232 6996 10284 7002
rect 10232 6938 10284 6944
rect 10414 6896 10470 6905
rect 10324 6860 10376 6866
rect 10414 6831 10416 6840
rect 10324 6802 10376 6808
rect 10468 6831 10470 6840
rect 10692 6860 10744 6866
rect 10416 6802 10468 6808
rect 10796 6848 10824 7919
rect 10888 7886 10916 8366
rect 10876 7880 10928 7886
rect 10876 7822 10928 7828
rect 10876 7540 10928 7546
rect 10876 7482 10928 7488
rect 10744 6820 10824 6848
rect 10692 6802 10744 6808
rect 10232 6656 10284 6662
rect 10232 6598 10284 6604
rect 10140 5568 10192 5574
rect 10046 5536 10102 5545
rect 10140 5510 10192 5516
rect 10046 5471 10102 5480
rect 9956 5364 10008 5370
rect 9956 5306 10008 5312
rect 10060 5234 10088 5471
rect 10138 5400 10194 5409
rect 10138 5335 10194 5344
rect 10152 5302 10180 5335
rect 10140 5296 10192 5302
rect 10140 5238 10192 5244
rect 10048 5228 10100 5234
rect 10048 5170 10100 5176
rect 10140 5092 10192 5098
rect 10140 5034 10192 5040
rect 10152 4826 10180 5034
rect 10140 4820 10192 4826
rect 10140 4762 10192 4768
rect 10244 4622 10272 6598
rect 10336 6458 10364 6802
rect 10324 6452 10376 6458
rect 10324 6394 10376 6400
rect 10428 6186 10456 6802
rect 10508 6792 10560 6798
rect 10508 6734 10560 6740
rect 10520 6633 10548 6734
rect 10506 6624 10562 6633
rect 10506 6559 10562 6568
rect 10888 6361 10916 7482
rect 10980 7410 11008 9472
rect 11060 9454 11112 9460
rect 11152 9512 11204 9518
rect 11152 9454 11204 9460
rect 11060 9376 11112 9382
rect 11060 9318 11112 9324
rect 11072 9042 11100 9318
rect 11164 9217 11192 9454
rect 11150 9208 11206 9217
rect 11150 9143 11206 9152
rect 11152 9104 11204 9110
rect 11152 9046 11204 9052
rect 11060 9036 11112 9042
rect 11060 8978 11112 8984
rect 11164 8634 11192 9046
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 11060 8560 11112 8566
rect 11060 8502 11112 8508
rect 11072 7886 11100 8502
rect 11060 7880 11112 7886
rect 11060 7822 11112 7828
rect 11152 7812 11204 7818
rect 11152 7754 11204 7760
rect 11060 7744 11112 7750
rect 11060 7686 11112 7692
rect 10968 7404 11020 7410
rect 10968 7346 11020 7352
rect 10874 6352 10930 6361
rect 10874 6287 10930 6296
rect 10416 6180 10468 6186
rect 10416 6122 10468 6128
rect 10364 6012 10740 6021
rect 10420 6010 10444 6012
rect 10500 6010 10524 6012
rect 10580 6010 10604 6012
rect 10660 6010 10684 6012
rect 10420 5958 10430 6010
rect 10674 5958 10684 6010
rect 10420 5956 10444 5958
rect 10500 5956 10524 5958
rect 10580 5956 10604 5958
rect 10660 5956 10684 5958
rect 10364 5947 10740 5956
rect 10416 5772 10468 5778
rect 10416 5714 10468 5720
rect 10428 5370 10456 5714
rect 10968 5636 11020 5642
rect 10968 5578 11020 5584
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 10416 5364 10468 5370
rect 10416 5306 10468 5312
rect 10364 4924 10740 4933
rect 10420 4922 10444 4924
rect 10500 4922 10524 4924
rect 10580 4922 10604 4924
rect 10660 4922 10684 4924
rect 10420 4870 10430 4922
rect 10674 4870 10684 4922
rect 10420 4868 10444 4870
rect 10500 4868 10524 4870
rect 10580 4868 10604 4870
rect 10660 4868 10684 4870
rect 10364 4859 10740 4868
rect 9956 4616 10008 4622
rect 9956 4558 10008 4564
rect 10232 4616 10284 4622
rect 10232 4558 10284 4564
rect 9824 3488 9904 3516
rect 9772 3470 9824 3476
rect 9968 3398 9996 4558
rect 10692 4072 10744 4078
rect 10046 4040 10102 4049
rect 10690 4040 10692 4049
rect 10744 4040 10746 4049
rect 10046 3975 10102 3984
rect 10232 4004 10284 4010
rect 10060 3482 10088 3975
rect 10796 4010 10824 5510
rect 10690 3975 10746 3984
rect 10784 4004 10836 4010
rect 10232 3946 10284 3952
rect 10784 3946 10836 3952
rect 10140 3936 10192 3942
rect 10140 3878 10192 3884
rect 10152 3602 10180 3878
rect 10244 3738 10272 3946
rect 10364 3836 10740 3845
rect 10420 3834 10444 3836
rect 10500 3834 10524 3836
rect 10580 3834 10604 3836
rect 10660 3834 10684 3836
rect 10420 3782 10430 3834
rect 10674 3782 10684 3834
rect 10420 3780 10444 3782
rect 10500 3780 10524 3782
rect 10580 3780 10604 3782
rect 10660 3780 10684 3782
rect 10364 3771 10740 3780
rect 10232 3732 10284 3738
rect 10232 3674 10284 3680
rect 10506 3632 10562 3641
rect 10140 3596 10192 3602
rect 10980 3602 11008 5578
rect 11072 5234 11100 7686
rect 11164 6866 11192 7754
rect 11256 6866 11284 12406
rect 11348 12345 11376 12786
rect 11440 12646 11468 14062
rect 11428 12640 11480 12646
rect 11428 12582 11480 12588
rect 11428 12436 11480 12442
rect 11428 12378 11480 12384
rect 11334 12336 11390 12345
rect 11334 12271 11390 12280
rect 11440 12220 11468 12378
rect 11348 12192 11468 12220
rect 11348 11694 11376 12192
rect 11428 12096 11480 12102
rect 11428 12038 11480 12044
rect 11440 11762 11468 12038
rect 11532 11762 11560 16390
rect 11624 15337 11652 16390
rect 11610 15328 11666 15337
rect 11610 15263 11666 15272
rect 11610 15192 11666 15201
rect 11610 15127 11666 15136
rect 11624 14414 11652 15127
rect 11716 14482 11744 16623
rect 11796 16040 11848 16046
rect 11796 15982 11848 15988
rect 11808 15706 11836 15982
rect 11796 15700 11848 15706
rect 11796 15642 11848 15648
rect 11796 15496 11848 15502
rect 11796 15438 11848 15444
rect 11808 15026 11836 15438
rect 11796 15020 11848 15026
rect 11796 14962 11848 14968
rect 11704 14476 11756 14482
rect 11704 14418 11756 14424
rect 11796 14476 11848 14482
rect 11796 14418 11848 14424
rect 11612 14408 11664 14414
rect 11612 14350 11664 14356
rect 11624 13852 11652 14350
rect 11808 14006 11836 14418
rect 11796 14000 11848 14006
rect 11796 13942 11848 13948
rect 11704 13864 11756 13870
rect 11624 13824 11704 13852
rect 11704 13806 11756 13812
rect 11704 13728 11756 13734
rect 11704 13670 11756 13676
rect 11716 13462 11744 13670
rect 11808 13462 11836 13942
rect 11704 13456 11756 13462
rect 11704 13398 11756 13404
rect 11796 13456 11848 13462
rect 11796 13398 11848 13404
rect 11900 13308 11928 18380
rect 11992 17728 12020 18770
rect 12084 18698 12112 18770
rect 12072 18692 12124 18698
rect 12072 18634 12124 18640
rect 12360 18426 12388 18770
rect 12348 18420 12400 18426
rect 12348 18362 12400 18368
rect 11992 17700 12112 17728
rect 11980 17604 12032 17610
rect 11980 17546 12032 17552
rect 11992 16658 12020 17546
rect 11980 16652 12032 16658
rect 11980 16594 12032 16600
rect 11980 16448 12032 16454
rect 11980 16390 12032 16396
rect 11992 15910 12020 16390
rect 11980 15904 12032 15910
rect 11980 15846 12032 15852
rect 12084 15722 12112 17700
rect 12348 17536 12400 17542
rect 12348 17478 12400 17484
rect 12440 17536 12492 17542
rect 12440 17478 12492 17484
rect 12360 16794 12388 17478
rect 12452 17202 12480 17478
rect 12440 17196 12492 17202
rect 12440 17138 12492 17144
rect 12348 16788 12400 16794
rect 12348 16730 12400 16736
rect 12256 16720 12308 16726
rect 12256 16662 12308 16668
rect 12164 16652 12216 16658
rect 12164 16594 12216 16600
rect 12176 16454 12204 16594
rect 12164 16448 12216 16454
rect 12164 16390 12216 16396
rect 11716 13280 11928 13308
rect 11992 15694 12112 15722
rect 11612 13184 11664 13190
rect 11612 13126 11664 13132
rect 11624 12306 11652 13126
rect 11612 12300 11664 12306
rect 11612 12242 11664 12248
rect 11428 11756 11480 11762
rect 11428 11698 11480 11704
rect 11520 11756 11572 11762
rect 11520 11698 11572 11704
rect 11336 11688 11388 11694
rect 11336 11630 11388 11636
rect 11348 10606 11376 11630
rect 11440 11286 11468 11698
rect 11428 11280 11480 11286
rect 11428 11222 11480 11228
rect 11532 11218 11560 11698
rect 11520 11212 11572 11218
rect 11520 11154 11572 11160
rect 11518 11112 11574 11121
rect 11518 11047 11520 11056
rect 11572 11047 11574 11056
rect 11520 11018 11572 11024
rect 11610 10976 11666 10985
rect 11610 10911 11666 10920
rect 11624 10674 11652 10911
rect 11612 10668 11664 10674
rect 11612 10610 11664 10616
rect 11336 10600 11388 10606
rect 11336 10542 11388 10548
rect 11428 10600 11480 10606
rect 11428 10542 11480 10548
rect 11440 10198 11468 10542
rect 11428 10192 11480 10198
rect 11428 10134 11480 10140
rect 11716 10130 11744 13280
rect 11992 13138 12020 15694
rect 12176 15638 12204 16390
rect 12268 16250 12296 16662
rect 12348 16652 12400 16658
rect 12348 16594 12400 16600
rect 12256 16244 12308 16250
rect 12256 16186 12308 16192
rect 12268 16114 12296 16186
rect 12256 16108 12308 16114
rect 12256 16050 12308 16056
rect 12360 16046 12388 16594
rect 12348 16040 12400 16046
rect 12348 15982 12400 15988
rect 12256 15972 12308 15978
rect 12256 15914 12308 15920
rect 12164 15632 12216 15638
rect 12070 15600 12126 15609
rect 12164 15574 12216 15580
rect 12070 15535 12126 15544
rect 12084 14958 12112 15535
rect 12268 15434 12296 15914
rect 12438 15872 12494 15881
rect 12438 15807 12494 15816
rect 12452 15570 12480 15807
rect 12440 15564 12492 15570
rect 12440 15506 12492 15512
rect 12256 15428 12308 15434
rect 12256 15370 12308 15376
rect 12164 15156 12216 15162
rect 12164 15098 12216 15104
rect 12440 15156 12492 15162
rect 12440 15098 12492 15104
rect 12176 15065 12204 15098
rect 12162 15056 12218 15065
rect 12162 14991 12218 15000
rect 12072 14952 12124 14958
rect 12070 14920 12072 14929
rect 12124 14920 12126 14929
rect 12070 14855 12126 14864
rect 12070 14648 12126 14657
rect 12070 14583 12126 14592
rect 12084 14414 12112 14583
rect 12072 14408 12124 14414
rect 12176 14385 12204 14991
rect 12256 14612 12308 14618
rect 12256 14554 12308 14560
rect 12072 14350 12124 14356
rect 12162 14376 12218 14385
rect 12162 14311 12218 14320
rect 12268 13841 12296 14554
rect 12348 14476 12400 14482
rect 12348 14418 12400 14424
rect 12360 14074 12388 14418
rect 12452 14414 12480 15098
rect 12440 14408 12492 14414
rect 12440 14350 12492 14356
rect 12348 14068 12400 14074
rect 12348 14010 12400 14016
rect 12254 13832 12310 13841
rect 12072 13796 12124 13802
rect 12254 13767 12310 13776
rect 12072 13738 12124 13744
rect 11900 13110 12020 13138
rect 11794 12336 11850 12345
rect 11794 12271 11796 12280
rect 11848 12271 11850 12280
rect 11796 12242 11848 12248
rect 11794 12064 11850 12073
rect 11794 11999 11850 12008
rect 11808 11694 11836 11999
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 11794 11384 11850 11393
rect 11794 11319 11850 11328
rect 11704 10124 11756 10130
rect 11808 10112 11836 11319
rect 11900 10266 11928 13110
rect 11980 12980 12032 12986
rect 11980 12922 12032 12928
rect 11992 10742 12020 12922
rect 12084 12782 12112 13738
rect 12256 13728 12308 13734
rect 12176 13688 12256 13716
rect 12072 12776 12124 12782
rect 12072 12718 12124 12724
rect 12084 12374 12112 12718
rect 12072 12368 12124 12374
rect 12072 12310 12124 12316
rect 12072 12164 12124 12170
rect 12072 12106 12124 12112
rect 12084 11354 12112 12106
rect 12176 11898 12204 13688
rect 12256 13670 12308 13676
rect 12452 13546 12480 14350
rect 12268 13518 12480 13546
rect 12268 13394 12296 13518
rect 12348 13456 12400 13462
rect 12348 13398 12400 13404
rect 12256 13388 12308 13394
rect 12256 13330 12308 13336
rect 12360 13308 12388 13398
rect 12360 13280 12480 13308
rect 12256 13252 12308 13258
rect 12256 13194 12308 13200
rect 12268 12866 12296 13194
rect 12346 12880 12402 12889
rect 12268 12838 12346 12866
rect 12346 12815 12402 12824
rect 12360 12782 12388 12815
rect 12348 12776 12400 12782
rect 12348 12718 12400 12724
rect 12452 12646 12480 13280
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 12346 12472 12402 12481
rect 12346 12407 12402 12416
rect 12256 12232 12308 12238
rect 12256 12174 12308 12180
rect 12164 11892 12216 11898
rect 12164 11834 12216 11840
rect 12072 11348 12124 11354
rect 12072 11290 12124 11296
rect 12072 11212 12124 11218
rect 12072 11154 12124 11160
rect 12084 10985 12112 11154
rect 12164 11076 12216 11082
rect 12164 11018 12216 11024
rect 12070 10976 12126 10985
rect 12070 10911 12126 10920
rect 11980 10736 12032 10742
rect 11980 10678 12032 10684
rect 12084 10674 12112 10911
rect 12072 10668 12124 10674
rect 12072 10610 12124 10616
rect 11980 10600 12032 10606
rect 12176 10554 12204 11018
rect 12268 10606 12296 12174
rect 12360 11626 12388 12407
rect 12452 11830 12480 12582
rect 12440 11824 12492 11830
rect 12440 11766 12492 11772
rect 12544 11642 12572 18770
rect 12820 18630 12848 19450
rect 12900 19168 12952 19174
rect 12900 19110 12952 19116
rect 12912 18970 12940 19110
rect 12900 18964 12952 18970
rect 12900 18906 12952 18912
rect 12808 18624 12860 18630
rect 12808 18566 12860 18572
rect 12992 18080 13044 18086
rect 12992 18022 13044 18028
rect 12714 17776 12770 17785
rect 13004 17746 13032 18022
rect 12714 17711 12716 17720
rect 12768 17711 12770 17720
rect 12900 17740 12952 17746
rect 12716 17682 12768 17688
rect 12900 17682 12952 17688
rect 12992 17740 13044 17746
rect 12992 17682 13044 17688
rect 12624 17536 12676 17542
rect 12624 17478 12676 17484
rect 12636 15162 12664 17478
rect 12728 17066 12756 17682
rect 12808 17672 12860 17678
rect 12808 17614 12860 17620
rect 12716 17060 12768 17066
rect 12716 17002 12768 17008
rect 12820 16697 12848 17614
rect 12806 16688 12862 16697
rect 12806 16623 12862 16632
rect 12912 16522 12940 17682
rect 13004 17542 13032 17682
rect 12992 17536 13044 17542
rect 12992 17478 13044 17484
rect 13096 17066 13124 19994
rect 13820 19916 13872 19922
rect 13820 19858 13872 19864
rect 13364 19612 13740 19621
rect 13420 19610 13444 19612
rect 13500 19610 13524 19612
rect 13580 19610 13604 19612
rect 13660 19610 13684 19612
rect 13420 19558 13430 19610
rect 13674 19558 13684 19610
rect 13420 19556 13444 19558
rect 13500 19556 13524 19558
rect 13580 19556 13604 19558
rect 13660 19556 13684 19558
rect 13364 19547 13740 19556
rect 13832 19514 13860 19858
rect 14384 19514 14412 19994
rect 13820 19508 13872 19514
rect 13820 19450 13872 19456
rect 14372 19508 14424 19514
rect 14372 19450 14424 19456
rect 14004 19304 14056 19310
rect 14004 19246 14056 19252
rect 14016 18970 14044 19246
rect 14372 19168 14424 19174
rect 14372 19110 14424 19116
rect 14384 18970 14412 19110
rect 13452 18964 13504 18970
rect 13452 18906 13504 18912
rect 14004 18964 14056 18970
rect 14004 18906 14056 18912
rect 14372 18964 14424 18970
rect 14372 18906 14424 18912
rect 13464 18834 13492 18906
rect 13176 18828 13228 18834
rect 13176 18770 13228 18776
rect 13452 18828 13504 18834
rect 13452 18770 13504 18776
rect 13912 18828 13964 18834
rect 13912 18770 13964 18776
rect 14372 18828 14424 18834
rect 14372 18770 14424 18776
rect 13188 18630 13216 18770
rect 13820 18760 13872 18766
rect 13266 18728 13322 18737
rect 13820 18702 13872 18708
rect 13266 18663 13322 18672
rect 13176 18624 13228 18630
rect 13176 18566 13228 18572
rect 13176 17808 13228 17814
rect 13176 17750 13228 17756
rect 13188 17202 13216 17750
rect 13176 17196 13228 17202
rect 13176 17138 13228 17144
rect 13280 17134 13308 18663
rect 13364 18524 13740 18533
rect 13420 18522 13444 18524
rect 13500 18522 13524 18524
rect 13580 18522 13604 18524
rect 13660 18522 13684 18524
rect 13420 18470 13430 18522
rect 13674 18470 13684 18522
rect 13420 18468 13444 18470
rect 13500 18468 13524 18470
rect 13580 18468 13604 18470
rect 13660 18468 13684 18470
rect 13364 18459 13740 18468
rect 13832 18154 13860 18702
rect 13924 18154 13952 18770
rect 14188 18420 14240 18426
rect 14188 18362 14240 18368
rect 14200 18222 14228 18362
rect 14188 18216 14240 18222
rect 14188 18158 14240 18164
rect 13820 18148 13872 18154
rect 13820 18090 13872 18096
rect 13912 18148 13964 18154
rect 13912 18090 13964 18096
rect 14384 18086 14412 18770
rect 14372 18080 14424 18086
rect 14370 18048 14372 18057
rect 14424 18048 14426 18057
rect 14370 17983 14426 17992
rect 13820 17876 13872 17882
rect 13820 17818 13872 17824
rect 13364 17436 13740 17445
rect 13420 17434 13444 17436
rect 13500 17434 13524 17436
rect 13580 17434 13604 17436
rect 13660 17434 13684 17436
rect 13420 17382 13430 17434
rect 13674 17382 13684 17434
rect 13420 17380 13444 17382
rect 13500 17380 13524 17382
rect 13580 17380 13604 17382
rect 13660 17380 13684 17382
rect 13364 17371 13740 17380
rect 13832 17338 13860 17818
rect 14464 17808 14516 17814
rect 14464 17750 14516 17756
rect 14188 17740 14240 17746
rect 14188 17682 14240 17688
rect 14200 17626 14228 17682
rect 13924 17610 14228 17626
rect 13912 17604 14228 17610
rect 13964 17598 14228 17604
rect 14476 17592 14504 17750
rect 14556 17604 14608 17610
rect 14476 17564 14556 17592
rect 13912 17546 13964 17552
rect 14556 17546 14608 17552
rect 13924 17338 13952 17546
rect 14280 17536 14332 17542
rect 14280 17478 14332 17484
rect 13820 17332 13872 17338
rect 13820 17274 13872 17280
rect 13912 17332 13964 17338
rect 13912 17274 13964 17280
rect 13268 17128 13320 17134
rect 13268 17070 13320 17076
rect 13912 17128 13964 17134
rect 13912 17070 13964 17076
rect 12992 17060 13044 17066
rect 12992 17002 13044 17008
rect 13084 17060 13136 17066
rect 13084 17002 13136 17008
rect 13636 17060 13688 17066
rect 13636 17002 13688 17008
rect 13004 16658 13032 17002
rect 13082 16688 13138 16697
rect 12992 16652 13044 16658
rect 13082 16623 13138 16632
rect 13188 16646 13400 16674
rect 13648 16658 13676 17002
rect 13728 16788 13780 16794
rect 13728 16730 13780 16736
rect 12992 16594 13044 16600
rect 12808 16516 12860 16522
rect 12808 16458 12860 16464
rect 12900 16516 12952 16522
rect 12900 16458 12952 16464
rect 12992 16516 13044 16522
rect 12992 16458 13044 16464
rect 12716 16448 12768 16454
rect 12716 16390 12768 16396
rect 12728 16114 12756 16390
rect 12716 16108 12768 16114
rect 12716 16050 12768 16056
rect 12716 15360 12768 15366
rect 12716 15302 12768 15308
rect 12624 15156 12676 15162
rect 12624 15098 12676 15104
rect 12728 15094 12756 15302
rect 12716 15088 12768 15094
rect 12716 15030 12768 15036
rect 12820 14906 12848 16458
rect 12912 15201 12940 16458
rect 13004 16114 13032 16458
rect 13096 16454 13124 16623
rect 13084 16448 13136 16454
rect 13084 16390 13136 16396
rect 12992 16108 13044 16114
rect 12992 16050 13044 16056
rect 13084 16108 13136 16114
rect 13084 16050 13136 16056
rect 12992 15360 13044 15366
rect 12992 15302 13044 15308
rect 12898 15192 12954 15201
rect 12898 15127 12954 15136
rect 12900 15088 12952 15094
rect 12900 15030 12952 15036
rect 12912 14958 12940 15030
rect 13004 14958 13032 15302
rect 12728 14878 12848 14906
rect 12900 14952 12952 14958
rect 12900 14894 12952 14900
rect 12992 14952 13044 14958
rect 12992 14894 13044 14900
rect 12728 14657 12756 14878
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 12900 14816 12952 14822
rect 12900 14758 12952 14764
rect 12714 14648 12770 14657
rect 12820 14618 12848 14758
rect 12714 14583 12770 14592
rect 12808 14612 12860 14618
rect 12808 14554 12860 14560
rect 12716 14544 12768 14550
rect 12716 14486 12768 14492
rect 12624 14476 12676 14482
rect 12624 14418 12676 14424
rect 12636 14385 12664 14418
rect 12622 14376 12678 14385
rect 12622 14311 12678 14320
rect 12624 14272 12676 14278
rect 12624 14214 12676 14220
rect 12636 13161 12664 14214
rect 12728 13569 12756 14486
rect 12820 14482 12848 14554
rect 12808 14476 12860 14482
rect 12808 14418 12860 14424
rect 12912 14362 12940 14758
rect 12820 14334 12940 14362
rect 12820 14074 12848 14334
rect 12808 14068 12860 14074
rect 12808 14010 12860 14016
rect 13004 13938 13032 14894
rect 12992 13932 13044 13938
rect 12992 13874 13044 13880
rect 12808 13864 12860 13870
rect 12860 13824 12940 13852
rect 12808 13806 12860 13812
rect 12714 13560 12770 13569
rect 12714 13495 12770 13504
rect 12806 13424 12862 13433
rect 12716 13388 12768 13394
rect 12806 13359 12862 13368
rect 12716 13330 12768 13336
rect 12622 13152 12678 13161
rect 12622 13087 12678 13096
rect 12624 12912 12676 12918
rect 12622 12880 12624 12889
rect 12676 12880 12678 12889
rect 12622 12815 12678 12824
rect 12728 12374 12756 13330
rect 12820 13326 12848 13359
rect 12808 13320 12860 13326
rect 12808 13262 12860 13268
rect 12820 12782 12848 13262
rect 12808 12776 12860 12782
rect 12808 12718 12860 12724
rect 12716 12368 12768 12374
rect 12716 12310 12768 12316
rect 12624 12164 12676 12170
rect 12624 12106 12676 12112
rect 12636 11937 12664 12106
rect 12622 11928 12678 11937
rect 12622 11863 12678 11872
rect 12912 11830 12940 13824
rect 12992 13184 13044 13190
rect 12992 13126 13044 13132
rect 12900 11824 12952 11830
rect 12900 11766 12952 11772
rect 12348 11620 12400 11626
rect 12348 11562 12400 11568
rect 12452 11614 12572 11642
rect 12622 11656 12678 11665
rect 12360 11286 12388 11562
rect 12348 11280 12400 11286
rect 12348 11222 12400 11228
rect 12256 10600 12308 10606
rect 12032 10548 12204 10554
rect 11980 10542 12204 10548
rect 11992 10526 12204 10542
rect 12072 10464 12124 10470
rect 12072 10406 12124 10412
rect 11888 10260 11940 10266
rect 11888 10202 11940 10208
rect 11888 10124 11940 10130
rect 11808 10084 11888 10112
rect 11704 10066 11756 10072
rect 11888 10066 11940 10072
rect 11716 9926 11744 10066
rect 11980 9988 12032 9994
rect 11980 9930 12032 9936
rect 11704 9920 11756 9926
rect 11756 9880 11928 9908
rect 11704 9862 11756 9868
rect 11900 9674 11928 9880
rect 11716 9646 11928 9674
rect 11612 9580 11664 9586
rect 11532 9540 11612 9568
rect 11336 9512 11388 9518
rect 11336 9454 11388 9460
rect 11428 9512 11480 9518
rect 11428 9454 11480 9460
rect 11348 9178 11376 9454
rect 11440 9178 11468 9454
rect 11532 9217 11560 9540
rect 11612 9522 11664 9528
rect 11716 9466 11744 9646
rect 11992 9602 12020 9930
rect 12084 9926 12112 10406
rect 12072 9920 12124 9926
rect 12072 9862 12124 9868
rect 12084 9722 12112 9862
rect 12072 9716 12124 9722
rect 12072 9658 12124 9664
rect 11992 9574 12112 9602
rect 11716 9438 11836 9466
rect 11704 9376 11756 9382
rect 11624 9336 11704 9364
rect 11518 9208 11574 9217
rect 11336 9172 11388 9178
rect 11336 9114 11388 9120
rect 11428 9172 11480 9178
rect 11518 9143 11574 9152
rect 11428 9114 11480 9120
rect 11336 8900 11388 8906
rect 11336 8842 11388 8848
rect 11348 8498 11376 8842
rect 11336 8492 11388 8498
rect 11336 8434 11388 8440
rect 11348 7886 11376 8434
rect 11624 8401 11652 9336
rect 11704 9318 11756 9324
rect 11702 9208 11758 9217
rect 11702 9143 11758 9152
rect 11716 8838 11744 9143
rect 11704 8832 11756 8838
rect 11704 8774 11756 8780
rect 11808 8514 11836 9438
rect 11980 8832 12032 8838
rect 11980 8774 12032 8780
rect 11808 8486 11928 8514
rect 11900 8430 11928 8486
rect 11704 8424 11756 8430
rect 11610 8392 11666 8401
rect 11704 8366 11756 8372
rect 11796 8424 11848 8430
rect 11796 8366 11848 8372
rect 11888 8424 11940 8430
rect 11888 8366 11940 8372
rect 11610 8327 11666 8336
rect 11520 8288 11572 8294
rect 11520 8230 11572 8236
rect 11336 7880 11388 7886
rect 11336 7822 11388 7828
rect 11532 7410 11560 8230
rect 11624 7546 11652 8327
rect 11716 8090 11744 8366
rect 11808 8294 11836 8366
rect 11796 8288 11848 8294
rect 11796 8230 11848 8236
rect 11704 8084 11756 8090
rect 11704 8026 11756 8032
rect 11808 8022 11836 8230
rect 11796 8016 11848 8022
rect 11796 7958 11848 7964
rect 11900 7954 11928 8366
rect 11888 7948 11940 7954
rect 11888 7890 11940 7896
rect 11704 7880 11756 7886
rect 11704 7822 11756 7828
rect 11612 7540 11664 7546
rect 11612 7482 11664 7488
rect 11520 7404 11572 7410
rect 11520 7346 11572 7352
rect 11612 7404 11664 7410
rect 11612 7346 11664 7352
rect 11624 7290 11652 7346
rect 11440 7262 11652 7290
rect 11716 7274 11744 7822
rect 11796 7744 11848 7750
rect 11796 7686 11848 7692
rect 11808 7342 11836 7686
rect 11796 7336 11848 7342
rect 11796 7278 11848 7284
rect 11704 7268 11756 7274
rect 11152 6860 11204 6866
rect 11152 6802 11204 6808
rect 11244 6860 11296 6866
rect 11244 6802 11296 6808
rect 11152 6656 11204 6662
rect 11152 6598 11204 6604
rect 11060 5228 11112 5234
rect 11060 5170 11112 5176
rect 11072 4434 11100 5170
rect 11164 4554 11192 6598
rect 11256 6458 11284 6802
rect 11440 6798 11468 7262
rect 11704 7210 11756 7216
rect 11796 7200 11848 7206
rect 11796 7142 11848 7148
rect 11888 7200 11940 7206
rect 11888 7142 11940 7148
rect 11702 7032 11758 7041
rect 11612 6996 11664 7002
rect 11702 6967 11704 6976
rect 11612 6938 11664 6944
rect 11756 6967 11758 6976
rect 11704 6938 11756 6944
rect 11624 6866 11652 6938
rect 11612 6860 11664 6866
rect 11612 6802 11664 6808
rect 11428 6792 11480 6798
rect 11428 6734 11480 6740
rect 11704 6792 11756 6798
rect 11704 6734 11756 6740
rect 11520 6724 11572 6730
rect 11520 6666 11572 6672
rect 11244 6452 11296 6458
rect 11244 6394 11296 6400
rect 11336 6384 11388 6390
rect 11336 6326 11388 6332
rect 11244 6180 11296 6186
rect 11244 6122 11296 6128
rect 11256 5642 11284 6122
rect 11348 5778 11376 6326
rect 11532 6202 11560 6666
rect 11716 6633 11744 6734
rect 11702 6624 11758 6633
rect 11702 6559 11758 6568
rect 11440 6174 11560 6202
rect 11440 6118 11468 6174
rect 11428 6112 11480 6118
rect 11428 6054 11480 6060
rect 11520 6112 11572 6118
rect 11520 6054 11572 6060
rect 11532 5778 11560 6054
rect 11336 5772 11388 5778
rect 11336 5714 11388 5720
rect 11428 5772 11480 5778
rect 11428 5714 11480 5720
rect 11520 5772 11572 5778
rect 11520 5714 11572 5720
rect 11244 5636 11296 5642
rect 11244 5578 11296 5584
rect 11334 5264 11390 5273
rect 11334 5199 11390 5208
rect 11348 5166 11376 5199
rect 11244 5160 11296 5166
rect 11244 5102 11296 5108
rect 11336 5160 11388 5166
rect 11336 5102 11388 5108
rect 11256 4622 11284 5102
rect 11334 4720 11390 4729
rect 11334 4655 11390 4664
rect 11244 4616 11296 4622
rect 11244 4558 11296 4564
rect 11152 4548 11204 4554
rect 11152 4490 11204 4496
rect 11072 4406 11284 4434
rect 11060 4208 11112 4214
rect 11060 4150 11112 4156
rect 10506 3567 10508 3576
rect 10140 3538 10192 3544
rect 10560 3567 10562 3576
rect 10968 3596 11020 3602
rect 10508 3538 10560 3544
rect 10968 3538 11020 3544
rect 10600 3528 10652 3534
rect 10230 3496 10286 3505
rect 10060 3454 10180 3482
rect 9956 3392 10008 3398
rect 9956 3334 10008 3340
rect 10048 3392 10100 3398
rect 10048 3334 10100 3340
rect 9588 2576 9640 2582
rect 9588 2518 9640 2524
rect 9680 2576 9732 2582
rect 9680 2518 9732 2524
rect 8484 2508 8536 2514
rect 8484 2450 8536 2456
rect 8760 2508 8812 2514
rect 8760 2450 8812 2456
rect 9496 2508 9548 2514
rect 9496 2450 9548 2456
rect 8944 2440 8996 2446
rect 8298 2408 8354 2417
rect 8944 2382 8996 2388
rect 8298 2343 8300 2352
rect 8352 2343 8354 2352
rect 8300 2314 8352 2320
rect 8116 2304 8168 2310
rect 8116 2246 8168 2252
rect 8128 1426 8156 2246
rect 8312 1562 8340 2314
rect 8760 2304 8812 2310
rect 8760 2246 8812 2252
rect 8772 2106 8800 2246
rect 8956 2106 8984 2382
rect 9128 2304 9180 2310
rect 9128 2246 9180 2252
rect 9404 2304 9456 2310
rect 9404 2246 9456 2252
rect 9600 2258 9628 2518
rect 10060 2514 10088 3334
rect 10152 2990 10180 3454
rect 10600 3470 10652 3476
rect 10692 3528 10744 3534
rect 10692 3470 10744 3476
rect 10784 3528 10836 3534
rect 10784 3470 10836 3476
rect 10230 3431 10286 3440
rect 10244 3058 10272 3431
rect 10324 3392 10376 3398
rect 10612 3369 10640 3470
rect 10324 3334 10376 3340
rect 10598 3360 10654 3369
rect 10232 3052 10284 3058
rect 10232 2994 10284 3000
rect 10140 2984 10192 2990
rect 10140 2926 10192 2932
rect 10336 2836 10364 3334
rect 10598 3295 10654 3304
rect 10704 3194 10732 3470
rect 10796 3194 10824 3470
rect 10692 3188 10744 3194
rect 10692 3130 10744 3136
rect 10784 3188 10836 3194
rect 10784 3130 10836 3136
rect 11072 2990 11100 4150
rect 11256 4078 11284 4406
rect 11348 4146 11376 4655
rect 11440 4214 11468 5714
rect 11612 5636 11664 5642
rect 11612 5578 11664 5584
rect 11520 5364 11572 5370
rect 11520 5306 11572 5312
rect 11532 4690 11560 5306
rect 11520 4684 11572 4690
rect 11520 4626 11572 4632
rect 11428 4208 11480 4214
rect 11428 4150 11480 4156
rect 11336 4140 11388 4146
rect 11336 4082 11388 4088
rect 11244 4072 11296 4078
rect 11244 4014 11296 4020
rect 11336 3936 11388 3942
rect 11336 3878 11388 3884
rect 11348 3602 11376 3878
rect 11336 3596 11388 3602
rect 11336 3538 11388 3544
rect 11428 3528 11480 3534
rect 11428 3470 11480 3476
rect 11334 3088 11390 3097
rect 11440 3074 11468 3470
rect 11518 3360 11574 3369
rect 11518 3295 11574 3304
rect 11532 3194 11560 3295
rect 11520 3188 11572 3194
rect 11520 3130 11572 3136
rect 11390 3046 11468 3074
rect 11334 3023 11390 3032
rect 11348 2990 11376 3023
rect 11532 2990 11560 3130
rect 11624 2990 11652 5578
rect 11704 5568 11756 5574
rect 11704 5510 11756 5516
rect 10784 2984 10836 2990
rect 10784 2926 10836 2932
rect 11060 2984 11112 2990
rect 11060 2926 11112 2932
rect 11244 2984 11296 2990
rect 11244 2926 11296 2932
rect 11336 2984 11388 2990
rect 11336 2926 11388 2932
rect 11520 2984 11572 2990
rect 11520 2926 11572 2932
rect 11612 2984 11664 2990
rect 11612 2926 11664 2932
rect 10244 2808 10364 2836
rect 10048 2508 10100 2514
rect 10244 2496 10272 2808
rect 10796 2802 10824 2926
rect 10966 2816 11022 2825
rect 10796 2774 10966 2802
rect 10364 2748 10740 2757
rect 10966 2751 11022 2760
rect 10420 2746 10444 2748
rect 10500 2746 10524 2748
rect 10580 2746 10604 2748
rect 10660 2746 10684 2748
rect 10420 2694 10430 2746
rect 10674 2694 10684 2746
rect 10420 2692 10444 2694
rect 10500 2692 10524 2694
rect 10580 2692 10604 2694
rect 10660 2692 10684 2694
rect 10364 2683 10740 2692
rect 10784 2644 10836 2650
rect 10784 2586 10836 2592
rect 10416 2508 10468 2514
rect 10244 2468 10364 2496
rect 10048 2450 10100 2456
rect 10230 2408 10286 2417
rect 9772 2372 9824 2378
rect 10230 2343 10286 2352
rect 9772 2314 9824 2320
rect 9678 2272 9734 2281
rect 8760 2100 8812 2106
rect 8760 2042 8812 2048
rect 8944 2100 8996 2106
rect 8944 2042 8996 2048
rect 9140 1902 9168 2246
rect 8484 1896 8536 1902
rect 8484 1838 8536 1844
rect 9128 1896 9180 1902
rect 9128 1838 9180 1844
rect 9312 1896 9364 1902
rect 9312 1838 9364 1844
rect 8300 1556 8352 1562
rect 8300 1498 8352 1504
rect 8496 1426 8524 1838
rect 8668 1828 8720 1834
rect 8668 1770 8720 1776
rect 9036 1828 9088 1834
rect 9036 1770 9088 1776
rect 8576 1488 8628 1494
rect 8680 1476 8708 1770
rect 8852 1760 8904 1766
rect 8852 1702 8904 1708
rect 8628 1448 8708 1476
rect 8576 1430 8628 1436
rect 8116 1420 8168 1426
rect 8116 1362 8168 1368
rect 8484 1420 8536 1426
rect 8484 1362 8536 1368
rect 8024 1284 8076 1290
rect 8024 1226 8076 1232
rect 7102 847 7158 856
rect 7932 876 7984 882
rect 7116 814 7144 847
rect 7932 818 7984 824
rect 7104 808 7156 814
rect 7104 750 7156 756
rect 7196 808 7248 814
rect 7196 750 7248 756
rect 7840 808 7892 814
rect 8036 762 8064 1226
rect 8496 1222 8524 1362
rect 8484 1216 8536 1222
rect 8484 1158 8536 1164
rect 8496 1018 8524 1158
rect 8484 1012 8536 1018
rect 8484 954 8536 960
rect 8864 814 8892 1702
rect 8942 1456 8998 1465
rect 9048 1442 9076 1770
rect 9140 1494 9168 1838
rect 9220 1760 9272 1766
rect 9220 1702 9272 1708
rect 8998 1414 9076 1442
rect 9128 1488 9180 1494
rect 9128 1430 9180 1436
rect 8942 1391 8944 1400
rect 8996 1391 8998 1400
rect 8944 1362 8996 1368
rect 9128 1352 9180 1358
rect 9128 1294 9180 1300
rect 7892 756 8064 762
rect 7840 750 8064 756
rect 8116 808 8168 814
rect 8116 750 8168 756
rect 8852 808 8904 814
rect 8852 750 8904 756
rect 5262 711 5318 720
rect 5540 740 5592 746
rect 5540 682 5592 688
rect 6736 740 6788 746
rect 6736 682 6788 688
rect 5552 400 5580 682
rect 5816 672 5868 678
rect 5868 632 5948 660
rect 5816 614 5868 620
rect 5920 400 5948 632
rect 7208 474 7236 750
rect 7852 734 8064 750
rect 7748 672 7800 678
rect 7748 614 7800 620
rect 7196 468 7248 474
rect 7196 410 7248 416
rect 7760 406 7788 614
rect 7748 400 7800 406
rect 4988 196 5040 202
rect 4988 138 5040 144
rect 5170 0 5226 400
rect 5538 0 5594 400
rect 5906 0 5962 400
rect 7748 342 7800 348
rect 8128 338 8156 750
rect 9140 746 9168 1294
rect 9128 740 9180 746
rect 9128 682 9180 688
rect 8116 332 8168 338
rect 8116 274 8168 280
rect 9140 134 9168 682
rect 9232 400 9260 1702
rect 9324 1562 9352 1838
rect 9312 1556 9364 1562
rect 9312 1498 9364 1504
rect 9416 1426 9444 2246
rect 9600 2230 9678 2258
rect 9678 2207 9734 2216
rect 9588 1760 9640 1766
rect 9508 1720 9588 1748
rect 9404 1420 9456 1426
rect 9404 1362 9456 1368
rect 9508 1358 9536 1720
rect 9784 1748 9812 2314
rect 9954 2136 10010 2145
rect 9954 2071 10010 2080
rect 9862 2000 9918 2009
rect 9862 1935 9918 1944
rect 9876 1902 9904 1935
rect 9968 1902 9996 2071
rect 10048 2032 10100 2038
rect 10048 1974 10100 1980
rect 9864 1896 9916 1902
rect 9864 1838 9916 1844
rect 9956 1896 10008 1902
rect 10060 1873 10088 1974
rect 10244 1902 10272 2343
rect 10336 1902 10364 2468
rect 10416 2450 10468 2456
rect 10428 2106 10456 2450
rect 10416 2100 10468 2106
rect 10416 2042 10468 2048
rect 10232 1896 10284 1902
rect 9956 1838 10008 1844
rect 10046 1864 10102 1873
rect 10232 1838 10284 1844
rect 10324 1896 10376 1902
rect 10324 1838 10376 1844
rect 10046 1799 10102 1808
rect 10796 1766 10824 2586
rect 11256 2564 11284 2926
rect 11520 2848 11572 2854
rect 11520 2790 11572 2796
rect 11610 2816 11666 2825
rect 11334 2680 11390 2689
rect 11532 2650 11560 2790
rect 11610 2751 11666 2760
rect 11716 2774 11744 5510
rect 11808 5166 11836 7142
rect 11900 6934 11928 7142
rect 11888 6928 11940 6934
rect 11888 6870 11940 6876
rect 11992 6118 12020 8774
rect 11980 6112 12032 6118
rect 11980 6054 12032 6060
rect 12084 5778 12112 9574
rect 12176 9042 12204 10526
rect 12254 10568 12256 10577
rect 12308 10568 12310 10577
rect 12452 10554 12480 11614
rect 12622 11591 12678 11600
rect 12530 11520 12586 11529
rect 12530 11455 12586 11464
rect 12544 10674 12572 11455
rect 12636 11014 12664 11591
rect 12808 11552 12860 11558
rect 12912 11540 12940 11766
rect 13004 11694 13032 13126
rect 13096 11762 13124 16050
rect 13188 14618 13216 16646
rect 13268 16584 13320 16590
rect 13268 16526 13320 16532
rect 13280 15094 13308 16526
rect 13372 16454 13400 16646
rect 13636 16652 13688 16658
rect 13636 16594 13688 16600
rect 13740 16590 13768 16730
rect 13728 16584 13780 16590
rect 13728 16526 13780 16532
rect 13360 16448 13412 16454
rect 13360 16390 13412 16396
rect 13364 16348 13740 16357
rect 13420 16346 13444 16348
rect 13500 16346 13524 16348
rect 13580 16346 13604 16348
rect 13660 16346 13684 16348
rect 13420 16294 13430 16346
rect 13674 16294 13684 16346
rect 13420 16292 13444 16294
rect 13500 16292 13524 16294
rect 13580 16292 13604 16294
rect 13660 16292 13684 16294
rect 13364 16283 13740 16292
rect 13544 16040 13596 16046
rect 13544 15982 13596 15988
rect 13556 15706 13584 15982
rect 13820 15972 13872 15978
rect 13820 15914 13872 15920
rect 13832 15706 13860 15914
rect 13544 15700 13596 15706
rect 13544 15642 13596 15648
rect 13820 15700 13872 15706
rect 13820 15642 13872 15648
rect 13820 15564 13872 15570
rect 13820 15506 13872 15512
rect 13364 15260 13740 15269
rect 13420 15258 13444 15260
rect 13500 15258 13524 15260
rect 13580 15258 13604 15260
rect 13660 15258 13684 15260
rect 13420 15206 13430 15258
rect 13674 15206 13684 15258
rect 13420 15204 13444 15206
rect 13500 15204 13524 15206
rect 13580 15204 13604 15206
rect 13660 15204 13684 15206
rect 13364 15195 13740 15204
rect 13268 15088 13320 15094
rect 13268 15030 13320 15036
rect 13728 15088 13780 15094
rect 13728 15030 13780 15036
rect 13740 14890 13768 15030
rect 13832 15026 13860 15506
rect 13924 15502 13952 17070
rect 14004 17060 14056 17066
rect 14004 17002 14056 17008
rect 14016 16658 14044 17002
rect 14004 16652 14056 16658
rect 14004 16594 14056 16600
rect 13912 15496 13964 15502
rect 13912 15438 13964 15444
rect 14096 15428 14148 15434
rect 14096 15370 14148 15376
rect 13820 15020 13872 15026
rect 13820 14962 13872 14968
rect 14004 14952 14056 14958
rect 14004 14894 14056 14900
rect 13728 14884 13780 14890
rect 13728 14826 13780 14832
rect 13912 14884 13964 14890
rect 13912 14826 13964 14832
rect 13268 14816 13320 14822
rect 13268 14758 13320 14764
rect 13176 14612 13228 14618
rect 13176 14554 13228 14560
rect 13280 14482 13308 14758
rect 13636 14612 13688 14618
rect 13636 14554 13688 14560
rect 13268 14476 13320 14482
rect 13268 14418 13320 14424
rect 13176 14408 13228 14414
rect 13176 14350 13228 14356
rect 13188 11801 13216 14350
rect 13648 14260 13676 14554
rect 13648 14232 13860 14260
rect 13364 14172 13740 14181
rect 13420 14170 13444 14172
rect 13500 14170 13524 14172
rect 13580 14170 13604 14172
rect 13660 14170 13684 14172
rect 13420 14118 13430 14170
rect 13674 14118 13684 14170
rect 13420 14116 13444 14118
rect 13500 14116 13524 14118
rect 13580 14116 13604 14118
rect 13660 14116 13684 14118
rect 13364 14107 13740 14116
rect 13360 14068 13412 14074
rect 13360 14010 13412 14016
rect 13268 13864 13320 13870
rect 13266 13832 13268 13841
rect 13320 13832 13322 13841
rect 13266 13767 13322 13776
rect 13372 13326 13400 14010
rect 13832 13870 13860 14232
rect 13924 13870 13952 14826
rect 14016 14482 14044 14894
rect 14108 14822 14136 15370
rect 14096 14816 14148 14822
rect 14096 14758 14148 14764
rect 14188 14816 14240 14822
rect 14188 14758 14240 14764
rect 14094 14512 14150 14521
rect 14004 14476 14056 14482
rect 14200 14482 14228 14758
rect 14094 14447 14150 14456
rect 14188 14476 14240 14482
rect 14004 14418 14056 14424
rect 13820 13864 13872 13870
rect 13740 13824 13820 13852
rect 13360 13320 13412 13326
rect 13360 13262 13412 13268
rect 13740 13258 13768 13824
rect 13820 13806 13872 13812
rect 13912 13864 13964 13870
rect 13912 13806 13964 13812
rect 14108 13462 14136 14447
rect 14188 14418 14240 14424
rect 14096 13456 14148 13462
rect 14096 13398 14148 13404
rect 13728 13252 13780 13258
rect 13728 13194 13780 13200
rect 13364 13084 13740 13093
rect 13420 13082 13444 13084
rect 13500 13082 13524 13084
rect 13580 13082 13604 13084
rect 13660 13082 13684 13084
rect 13420 13030 13430 13082
rect 13674 13030 13684 13082
rect 13420 13028 13444 13030
rect 13500 13028 13524 13030
rect 13580 13028 13604 13030
rect 13660 13028 13684 13030
rect 13364 13019 13740 13028
rect 13910 12880 13966 12889
rect 13910 12815 13966 12824
rect 13268 12232 13320 12238
rect 13268 12174 13320 12180
rect 13174 11792 13230 11801
rect 13084 11756 13136 11762
rect 13174 11727 13230 11736
rect 13084 11698 13136 11704
rect 13280 11694 13308 12174
rect 13820 12096 13872 12102
rect 13820 12038 13872 12044
rect 13364 11996 13740 12005
rect 13420 11994 13444 11996
rect 13500 11994 13524 11996
rect 13580 11994 13604 11996
rect 13660 11994 13684 11996
rect 13420 11942 13430 11994
rect 13674 11942 13684 11994
rect 13420 11940 13444 11942
rect 13500 11940 13524 11942
rect 13580 11940 13604 11942
rect 13660 11940 13684 11942
rect 13364 11931 13740 11940
rect 13728 11824 13780 11830
rect 13728 11766 13780 11772
rect 12992 11688 13044 11694
rect 12992 11630 13044 11636
rect 13268 11688 13320 11694
rect 13268 11630 13320 11636
rect 13542 11656 13598 11665
rect 13084 11620 13136 11626
rect 13542 11591 13598 11600
rect 13084 11562 13136 11568
rect 12912 11512 13032 11540
rect 12808 11494 12860 11500
rect 12714 11248 12770 11257
rect 12714 11183 12770 11192
rect 12624 11008 12676 11014
rect 12624 10950 12676 10956
rect 12532 10668 12584 10674
rect 12532 10610 12584 10616
rect 12624 10600 12676 10606
rect 12452 10526 12572 10554
rect 12728 10588 12756 11183
rect 12820 11121 12848 11494
rect 12806 11112 12862 11121
rect 12806 11047 12862 11056
rect 12808 11008 12860 11014
rect 12806 10976 12808 10985
rect 12860 10976 12862 10985
rect 12806 10911 12862 10920
rect 12900 10668 12952 10674
rect 12900 10610 12952 10616
rect 12676 10560 12756 10588
rect 12624 10542 12676 10548
rect 12254 10503 12310 10512
rect 12440 10464 12492 10470
rect 12254 10432 12310 10441
rect 12440 10406 12492 10412
rect 12254 10367 12310 10376
rect 12268 10180 12296 10367
rect 12348 10192 12400 10198
rect 12268 10152 12348 10180
rect 12348 10134 12400 10140
rect 12256 9580 12308 9586
rect 12256 9522 12308 9528
rect 12164 9036 12216 9042
rect 12164 8978 12216 8984
rect 12268 8838 12296 9522
rect 12256 8832 12308 8838
rect 12256 8774 12308 8780
rect 12348 8832 12400 8838
rect 12348 8774 12400 8780
rect 12164 8628 12216 8634
rect 12164 8570 12216 8576
rect 12176 8022 12204 8570
rect 12360 8566 12388 8774
rect 12348 8560 12400 8566
rect 12348 8502 12400 8508
rect 12452 8514 12480 10406
rect 12544 9926 12572 10526
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 12532 9920 12584 9926
rect 12532 9862 12584 9868
rect 12544 9761 12572 9862
rect 12530 9752 12586 9761
rect 12530 9687 12586 9696
rect 12530 9480 12586 9489
rect 12530 9415 12586 9424
rect 12544 9178 12572 9415
rect 12532 9172 12584 9178
rect 12532 9114 12584 9120
rect 12636 8566 12664 10202
rect 12728 9722 12756 10406
rect 12912 10266 12940 10610
rect 13004 10606 13032 11512
rect 13096 11286 13124 11562
rect 13556 11286 13584 11591
rect 13740 11540 13768 11766
rect 13832 11694 13860 12038
rect 13820 11688 13872 11694
rect 13820 11630 13872 11636
rect 13740 11512 13860 11540
rect 13084 11280 13136 11286
rect 13544 11280 13596 11286
rect 13084 11222 13136 11228
rect 13174 11248 13230 11257
rect 13096 11121 13124 11222
rect 13544 11222 13596 11228
rect 13360 11212 13412 11218
rect 13174 11183 13176 11192
rect 13228 11183 13230 11192
rect 13176 11154 13228 11160
rect 13280 11172 13360 11200
rect 13082 11112 13138 11121
rect 13082 11047 13138 11056
rect 13176 11076 13228 11082
rect 13176 11018 13228 11024
rect 13082 10840 13138 10849
rect 13082 10775 13138 10784
rect 12992 10600 13044 10606
rect 12992 10542 13044 10548
rect 13096 10266 13124 10775
rect 12900 10260 12952 10266
rect 12900 10202 12952 10208
rect 13084 10260 13136 10266
rect 13084 10202 13136 10208
rect 12900 10056 12952 10062
rect 12952 10016 13032 10044
rect 12900 9998 12952 10004
rect 12808 9920 12860 9926
rect 12808 9862 12860 9868
rect 12716 9716 12768 9722
rect 12716 9658 12768 9664
rect 12716 9512 12768 9518
rect 12716 9454 12768 9460
rect 12624 8560 12676 8566
rect 12452 8486 12572 8514
rect 12624 8502 12676 8508
rect 12440 8424 12492 8430
rect 12440 8366 12492 8372
rect 12452 8090 12480 8366
rect 12440 8084 12492 8090
rect 12440 8026 12492 8032
rect 12164 8016 12216 8022
rect 12164 7958 12216 7964
rect 12544 7154 12572 8486
rect 12728 8129 12756 9454
rect 12820 9450 12848 9862
rect 12900 9580 12952 9586
rect 12900 9522 12952 9528
rect 12808 9444 12860 9450
rect 12808 9386 12860 9392
rect 12806 9208 12862 9217
rect 12806 9143 12862 9152
rect 12820 8430 12848 9143
rect 12912 8838 12940 9522
rect 12900 8832 12952 8838
rect 12900 8774 12952 8780
rect 13004 8514 13032 10016
rect 13084 9648 13136 9654
rect 13084 9590 13136 9596
rect 12912 8486 13032 8514
rect 12808 8424 12860 8430
rect 12808 8366 12860 8372
rect 12714 8120 12770 8129
rect 12820 8090 12848 8366
rect 12714 8055 12770 8064
rect 12808 8084 12860 8090
rect 12452 7126 12572 7154
rect 12452 6458 12480 7126
rect 12532 6996 12584 7002
rect 12532 6938 12584 6944
rect 12440 6452 12492 6458
rect 12440 6394 12492 6400
rect 12440 6316 12492 6322
rect 12440 6258 12492 6264
rect 11888 5772 11940 5778
rect 11888 5714 11940 5720
rect 12072 5772 12124 5778
rect 12072 5714 12124 5720
rect 11900 5370 11928 5714
rect 11888 5364 11940 5370
rect 11888 5306 11940 5312
rect 11796 5160 11848 5166
rect 12164 5160 12216 5166
rect 11848 5108 11928 5114
rect 11796 5102 11928 5108
rect 12164 5102 12216 5108
rect 12346 5128 12402 5137
rect 11808 5086 11928 5102
rect 11900 4690 11928 5086
rect 11888 4684 11940 4690
rect 11888 4626 11940 4632
rect 11796 4208 11848 4214
rect 11796 4150 11848 4156
rect 11808 4078 11836 4150
rect 11796 4072 11848 4078
rect 11796 4014 11848 4020
rect 11796 3936 11848 3942
rect 11796 3878 11848 3884
rect 11808 3058 11836 3878
rect 11900 3602 11928 4626
rect 12176 4622 12204 5102
rect 12346 5063 12402 5072
rect 12256 5024 12308 5030
rect 12254 4992 12256 5001
rect 12308 4992 12310 5001
rect 12254 4927 12310 4936
rect 12254 4856 12310 4865
rect 12254 4791 12256 4800
rect 12308 4791 12310 4800
rect 12256 4762 12308 4768
rect 12164 4616 12216 4622
rect 12360 4570 12388 5063
rect 12164 4558 12216 4564
rect 12268 4542 12388 4570
rect 12268 3992 12296 4542
rect 12348 4480 12400 4486
rect 12348 4422 12400 4428
rect 12084 3964 12296 3992
rect 11980 3936 12032 3942
rect 11980 3878 12032 3884
rect 11888 3596 11940 3602
rect 11888 3538 11940 3544
rect 11992 3482 12020 3878
rect 12084 3602 12112 3964
rect 12360 3602 12388 4422
rect 12452 4078 12480 6258
rect 12544 4282 12572 6938
rect 12728 6780 12756 8055
rect 12808 8026 12860 8032
rect 12808 6792 12860 6798
rect 12728 6752 12808 6780
rect 12808 6734 12860 6740
rect 12808 6656 12860 6662
rect 12808 6598 12860 6604
rect 12716 5772 12768 5778
rect 12716 5714 12768 5720
rect 12728 5370 12756 5714
rect 12716 5364 12768 5370
rect 12716 5306 12768 5312
rect 12716 5024 12768 5030
rect 12622 4992 12678 5001
rect 12716 4966 12768 4972
rect 12622 4927 12678 4936
rect 12636 4758 12664 4927
rect 12624 4752 12676 4758
rect 12624 4694 12676 4700
rect 12728 4282 12756 4966
rect 12532 4276 12584 4282
rect 12532 4218 12584 4224
rect 12716 4276 12768 4282
rect 12716 4218 12768 4224
rect 12820 4078 12848 6598
rect 12912 6066 12940 8486
rect 13096 8430 13124 9590
rect 12992 8424 13044 8430
rect 12992 8366 13044 8372
rect 13084 8424 13136 8430
rect 13084 8366 13136 8372
rect 13004 7410 13032 8366
rect 13084 8288 13136 8294
rect 13084 8230 13136 8236
rect 12992 7404 13044 7410
rect 12992 7346 13044 7352
rect 13096 7002 13124 8230
rect 13084 6996 13136 7002
rect 13084 6938 13136 6944
rect 13084 6860 13136 6866
rect 13084 6802 13136 6808
rect 13096 6186 13124 6802
rect 13084 6180 13136 6186
rect 13084 6122 13136 6128
rect 12990 6080 13046 6089
rect 12912 6038 12990 6066
rect 12990 6015 13046 6024
rect 13004 5914 13032 6015
rect 13096 5914 13124 6122
rect 12992 5908 13044 5914
rect 12992 5850 13044 5856
rect 13084 5908 13136 5914
rect 13084 5850 13136 5856
rect 12992 5364 13044 5370
rect 12992 5306 13044 5312
rect 12900 5296 12952 5302
rect 12898 5264 12900 5273
rect 12952 5264 12954 5273
rect 13004 5234 13032 5306
rect 12898 5199 12954 5208
rect 12992 5228 13044 5234
rect 12992 5170 13044 5176
rect 13004 5114 13032 5170
rect 12912 5086 13032 5114
rect 12912 4729 12940 5086
rect 12992 5024 13044 5030
rect 12992 4966 13044 4972
rect 12898 4720 12954 4729
rect 13004 4690 13032 4966
rect 13188 4690 13216 11018
rect 13280 10470 13308 11172
rect 13360 11154 13412 11160
rect 13364 10908 13740 10917
rect 13420 10906 13444 10908
rect 13500 10906 13524 10908
rect 13580 10906 13604 10908
rect 13660 10906 13684 10908
rect 13420 10854 13430 10906
rect 13674 10854 13684 10906
rect 13420 10852 13444 10854
rect 13500 10852 13524 10854
rect 13580 10852 13604 10854
rect 13660 10852 13684 10854
rect 13364 10843 13740 10852
rect 13832 10742 13860 11512
rect 13820 10736 13872 10742
rect 13820 10678 13872 10684
rect 13924 10606 13952 12815
rect 14108 12374 14136 13398
rect 14188 13184 14240 13190
rect 14188 13126 14240 13132
rect 14200 12782 14228 13126
rect 14188 12776 14240 12782
rect 14188 12718 14240 12724
rect 14096 12368 14148 12374
rect 14096 12310 14148 12316
rect 14292 12238 14320 17478
rect 14372 17128 14424 17134
rect 14372 17070 14424 17076
rect 14384 16998 14412 17070
rect 14372 16992 14424 16998
rect 14372 16934 14424 16940
rect 14556 16992 14608 16998
rect 14556 16934 14608 16940
rect 14384 16794 14412 16934
rect 14372 16788 14424 16794
rect 14372 16730 14424 16736
rect 14568 16658 14596 16934
rect 14556 16652 14608 16658
rect 14556 16594 14608 16600
rect 14660 15994 14688 21134
rect 14740 21072 14792 21078
rect 14740 21014 14792 21020
rect 14752 20398 14780 21014
rect 14832 21004 14884 21010
rect 14832 20946 14884 20952
rect 14844 20602 14872 20946
rect 14832 20596 14884 20602
rect 14832 20538 14884 20544
rect 14844 20448 14872 20538
rect 14924 20460 14976 20466
rect 14844 20420 14924 20448
rect 14924 20402 14976 20408
rect 14740 20392 14792 20398
rect 14740 20334 14792 20340
rect 14740 19984 14792 19990
rect 14740 19926 14792 19932
rect 14752 19718 14780 19926
rect 14832 19848 14884 19854
rect 14832 19790 14884 19796
rect 14740 19712 14792 19718
rect 14740 19654 14792 19660
rect 14844 19514 14872 19790
rect 14924 19780 14976 19786
rect 14924 19722 14976 19728
rect 14832 19508 14884 19514
rect 14832 19450 14884 19456
rect 14936 19242 14964 19722
rect 14924 19236 14976 19242
rect 14924 19178 14976 19184
rect 14740 18352 14792 18358
rect 14740 18294 14792 18300
rect 14752 17066 14780 18294
rect 14832 18080 14884 18086
rect 14832 18022 14884 18028
rect 14740 17060 14792 17066
rect 14740 17002 14792 17008
rect 14752 16969 14780 17002
rect 14738 16960 14794 16969
rect 14738 16895 14794 16904
rect 14844 16658 14872 18022
rect 14924 17196 14976 17202
rect 14924 17138 14976 17144
rect 14936 16726 14964 17138
rect 14924 16720 14976 16726
rect 14924 16662 14976 16668
rect 14832 16652 14884 16658
rect 14832 16594 14884 16600
rect 14568 15966 14688 15994
rect 14372 14952 14424 14958
rect 14372 14894 14424 14900
rect 14384 14414 14412 14894
rect 14568 14822 14596 15966
rect 14648 15904 14700 15910
rect 14648 15846 14700 15852
rect 14556 14816 14608 14822
rect 14556 14758 14608 14764
rect 14372 14408 14424 14414
rect 14372 14350 14424 14356
rect 14384 14074 14412 14350
rect 14556 14272 14608 14278
rect 14554 14240 14556 14249
rect 14608 14240 14610 14249
rect 14554 14175 14610 14184
rect 14372 14068 14424 14074
rect 14372 14010 14424 14016
rect 14556 13728 14608 13734
rect 14556 13670 14608 13676
rect 14464 12912 14516 12918
rect 14568 12900 14596 13670
rect 14516 12872 14596 12900
rect 14464 12854 14516 12860
rect 14372 12640 14424 12646
rect 14372 12582 14424 12588
rect 14464 12640 14516 12646
rect 14464 12582 14516 12588
rect 14096 12232 14148 12238
rect 14096 12174 14148 12180
rect 14280 12232 14332 12238
rect 14280 12174 14332 12180
rect 14108 11558 14136 12174
rect 14186 11928 14242 11937
rect 14186 11863 14242 11872
rect 14280 11892 14332 11898
rect 14200 11694 14228 11863
rect 14280 11834 14332 11840
rect 14188 11688 14240 11694
rect 14186 11656 14188 11665
rect 14240 11656 14242 11665
rect 14186 11591 14242 11600
rect 14096 11552 14148 11558
rect 14096 11494 14148 11500
rect 14188 11552 14240 11558
rect 14188 11494 14240 11500
rect 14004 11348 14056 11354
rect 14004 11290 14056 11296
rect 14016 10810 14044 11290
rect 14200 11218 14228 11494
rect 14292 11257 14320 11834
rect 14384 11762 14412 12582
rect 14476 12306 14504 12582
rect 14464 12300 14516 12306
rect 14464 12242 14516 12248
rect 14372 11756 14424 11762
rect 14372 11698 14424 11704
rect 14370 11656 14426 11665
rect 14370 11591 14426 11600
rect 14278 11248 14334 11257
rect 14188 11212 14240 11218
rect 14278 11183 14334 11192
rect 14188 11154 14240 11160
rect 14280 11144 14332 11150
rect 14186 11112 14242 11121
rect 14280 11086 14332 11092
rect 14384 11098 14412 11591
rect 14464 11552 14516 11558
rect 14464 11494 14516 11500
rect 14476 11218 14504 11494
rect 14464 11212 14516 11218
rect 14464 11154 14516 11160
rect 14186 11047 14242 11056
rect 14004 10804 14056 10810
rect 14004 10746 14056 10752
rect 13360 10600 13412 10606
rect 13912 10600 13964 10606
rect 13360 10542 13412 10548
rect 13450 10568 13506 10577
rect 13268 10464 13320 10470
rect 13268 10406 13320 10412
rect 13280 9654 13308 10406
rect 13372 10130 13400 10542
rect 13964 10560 14044 10588
rect 13912 10542 13964 10548
rect 13450 10503 13506 10512
rect 13360 10124 13412 10130
rect 13360 10066 13412 10072
rect 13464 10062 13492 10503
rect 13912 10464 13964 10470
rect 13912 10406 13964 10412
rect 13634 10296 13690 10305
rect 13634 10231 13690 10240
rect 13648 10130 13676 10231
rect 13636 10124 13688 10130
rect 13636 10066 13688 10072
rect 13452 10056 13504 10062
rect 13452 9998 13504 10004
rect 13820 10056 13872 10062
rect 13820 9998 13872 10004
rect 13364 9820 13740 9829
rect 13420 9818 13444 9820
rect 13500 9818 13524 9820
rect 13580 9818 13604 9820
rect 13660 9818 13684 9820
rect 13420 9766 13430 9818
rect 13674 9766 13684 9818
rect 13420 9764 13444 9766
rect 13500 9764 13524 9766
rect 13580 9764 13604 9766
rect 13660 9764 13684 9766
rect 13364 9755 13740 9764
rect 13268 9648 13320 9654
rect 13268 9590 13320 9596
rect 13832 9518 13860 9998
rect 13924 9738 13952 10406
rect 14016 9874 14044 10560
rect 14016 9846 14136 9874
rect 13924 9710 14044 9738
rect 14016 9636 14044 9710
rect 14108 9654 14136 9846
rect 13924 9608 14044 9636
rect 14096 9648 14148 9654
rect 13820 9512 13872 9518
rect 13820 9454 13872 9460
rect 13268 9376 13320 9382
rect 13268 9318 13320 9324
rect 13280 5710 13308 9318
rect 13818 9208 13874 9217
rect 13818 9143 13874 9152
rect 13832 9110 13860 9143
rect 13820 9104 13872 9110
rect 13820 9046 13872 9052
rect 13820 8832 13872 8838
rect 13820 8774 13872 8780
rect 13364 8732 13740 8741
rect 13420 8730 13444 8732
rect 13500 8730 13524 8732
rect 13580 8730 13604 8732
rect 13660 8730 13684 8732
rect 13420 8678 13430 8730
rect 13674 8678 13684 8730
rect 13420 8676 13444 8678
rect 13500 8676 13524 8678
rect 13580 8676 13604 8678
rect 13660 8676 13684 8678
rect 13364 8667 13740 8676
rect 13832 8498 13860 8774
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 13544 8424 13596 8430
rect 13544 8366 13596 8372
rect 13556 7954 13584 8366
rect 13544 7948 13596 7954
rect 13544 7890 13596 7896
rect 13364 7644 13740 7653
rect 13420 7642 13444 7644
rect 13500 7642 13524 7644
rect 13580 7642 13604 7644
rect 13660 7642 13684 7644
rect 13420 7590 13430 7642
rect 13674 7590 13684 7642
rect 13420 7588 13444 7590
rect 13500 7588 13524 7590
rect 13580 7588 13604 7590
rect 13660 7588 13684 7590
rect 13364 7579 13740 7588
rect 13636 7336 13688 7342
rect 13634 7304 13636 7313
rect 13924 7313 13952 9608
rect 14096 9590 14148 9596
rect 14004 9376 14056 9382
rect 14004 9318 14056 9324
rect 13688 7304 13690 7313
rect 13634 7239 13690 7248
rect 13910 7304 13966 7313
rect 13910 7239 13966 7248
rect 13912 6792 13964 6798
rect 13910 6760 13912 6769
rect 13964 6760 13966 6769
rect 13910 6695 13966 6704
rect 13364 6556 13740 6565
rect 13420 6554 13444 6556
rect 13500 6554 13524 6556
rect 13580 6554 13604 6556
rect 13660 6554 13684 6556
rect 13420 6502 13430 6554
rect 13674 6502 13684 6554
rect 13420 6500 13444 6502
rect 13500 6500 13524 6502
rect 13580 6500 13604 6502
rect 13660 6500 13684 6502
rect 13364 6491 13740 6500
rect 14016 6254 14044 9318
rect 14108 9042 14136 9590
rect 14096 9036 14148 9042
rect 14096 8978 14148 8984
rect 14096 8424 14148 8430
rect 14096 8366 14148 8372
rect 14108 7818 14136 8366
rect 14096 7812 14148 7818
rect 14096 7754 14148 7760
rect 14200 7342 14228 11047
rect 14292 10470 14320 11086
rect 14384 11070 14504 11098
rect 14372 10736 14424 10742
rect 14372 10678 14424 10684
rect 14280 10464 14332 10470
rect 14280 10406 14332 10412
rect 14278 10024 14334 10033
rect 14278 9959 14334 9968
rect 14292 9518 14320 9959
rect 14280 9512 14332 9518
rect 14280 9454 14332 9460
rect 14280 9376 14332 9382
rect 14280 9318 14332 9324
rect 14188 7336 14240 7342
rect 14188 7278 14240 7284
rect 14096 7200 14148 7206
rect 14096 7142 14148 7148
rect 14188 7200 14240 7206
rect 14188 7142 14240 7148
rect 14108 6866 14136 7142
rect 14200 6866 14228 7142
rect 14096 6860 14148 6866
rect 14096 6802 14148 6808
rect 14188 6860 14240 6866
rect 14188 6802 14240 6808
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 14004 6248 14056 6254
rect 14004 6190 14056 6196
rect 14016 5778 14044 6190
rect 14004 5772 14056 5778
rect 14004 5714 14056 5720
rect 13268 5704 13320 5710
rect 13268 5646 13320 5652
rect 13280 5166 13308 5646
rect 13912 5568 13964 5574
rect 13912 5510 13964 5516
rect 13364 5468 13740 5477
rect 13420 5466 13444 5468
rect 13500 5466 13524 5468
rect 13580 5466 13604 5468
rect 13660 5466 13684 5468
rect 13420 5414 13430 5466
rect 13674 5414 13684 5466
rect 13420 5412 13444 5414
rect 13500 5412 13524 5414
rect 13580 5412 13604 5414
rect 13660 5412 13684 5414
rect 13364 5403 13740 5412
rect 13268 5160 13320 5166
rect 13268 5102 13320 5108
rect 13820 5160 13872 5166
rect 13820 5102 13872 5108
rect 12898 4655 12954 4664
rect 12992 4684 13044 4690
rect 12992 4626 13044 4632
rect 13176 4684 13228 4690
rect 13176 4626 13228 4632
rect 12900 4616 12952 4622
rect 12898 4584 12900 4593
rect 12952 4584 12954 4593
rect 12898 4519 12954 4528
rect 13176 4548 13228 4554
rect 13176 4490 13228 4496
rect 12440 4072 12492 4078
rect 12440 4014 12492 4020
rect 12808 4072 12860 4078
rect 12808 4014 12860 4020
rect 12900 4072 12952 4078
rect 12900 4014 12952 4020
rect 12072 3596 12124 3602
rect 12072 3538 12124 3544
rect 12348 3596 12400 3602
rect 12348 3538 12400 3544
rect 12452 3534 12480 4014
rect 12624 4004 12676 4010
rect 12624 3946 12676 3952
rect 12636 3670 12664 3946
rect 12808 3936 12860 3942
rect 12808 3878 12860 3884
rect 12624 3664 12676 3670
rect 12624 3606 12676 3612
rect 11900 3454 12020 3482
rect 12440 3528 12492 3534
rect 12440 3470 12492 3476
rect 12820 3466 12848 3878
rect 12912 3738 12940 4014
rect 13188 3942 13216 4490
rect 13268 4480 13320 4486
rect 13268 4422 13320 4428
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 13176 3936 13228 3942
rect 13176 3878 13228 3884
rect 12900 3732 12952 3738
rect 12900 3674 12952 3680
rect 12808 3460 12860 3466
rect 11900 3194 11928 3454
rect 12808 3402 12860 3408
rect 11980 3392 12032 3398
rect 11980 3334 12032 3340
rect 11888 3188 11940 3194
rect 11888 3130 11940 3136
rect 11796 3052 11848 3058
rect 11796 2994 11848 3000
rect 11334 2615 11336 2624
rect 11388 2615 11390 2624
rect 11520 2644 11572 2650
rect 11336 2586 11388 2592
rect 11520 2586 11572 2592
rect 11072 2536 11284 2564
rect 10968 2508 11020 2514
rect 10968 2450 11020 2456
rect 10980 2417 11008 2450
rect 10966 2408 11022 2417
rect 10966 2343 11022 2352
rect 10876 1896 10928 1902
rect 10928 1856 11008 1884
rect 10876 1838 10928 1844
rect 10784 1760 10836 1766
rect 9784 1720 9996 1748
rect 9588 1702 9640 1708
rect 9772 1420 9824 1426
rect 9772 1362 9824 1368
rect 9496 1352 9548 1358
rect 9496 1294 9548 1300
rect 9680 1284 9732 1290
rect 9680 1226 9732 1232
rect 9588 944 9640 950
rect 9588 886 9640 892
rect 9312 876 9364 882
rect 9312 818 9364 824
rect 9324 406 9352 818
rect 9312 400 9364 406
rect 9600 400 9628 886
rect 9692 474 9720 1226
rect 9784 814 9812 1362
rect 9968 1358 9996 1720
rect 10784 1702 10836 1708
rect 10364 1660 10740 1669
rect 10420 1658 10444 1660
rect 10500 1658 10524 1660
rect 10580 1658 10604 1660
rect 10660 1658 10684 1660
rect 10420 1606 10430 1658
rect 10674 1606 10684 1658
rect 10420 1604 10444 1606
rect 10500 1604 10524 1606
rect 10580 1604 10604 1606
rect 10660 1604 10684 1606
rect 10364 1595 10740 1604
rect 10980 1465 11008 1856
rect 10966 1456 11022 1465
rect 10704 1414 10916 1442
rect 9956 1352 10008 1358
rect 9862 1320 9918 1329
rect 9956 1294 10008 1300
rect 10048 1352 10100 1358
rect 10048 1294 10100 1300
rect 9862 1255 9864 1264
rect 9916 1255 9918 1264
rect 9864 1226 9916 1232
rect 9956 1012 10008 1018
rect 9956 954 10008 960
rect 9772 808 9824 814
rect 9772 750 9824 756
rect 9864 672 9916 678
rect 9864 614 9916 620
rect 9876 474 9904 614
rect 9680 468 9732 474
rect 9680 410 9732 416
rect 9864 468 9916 474
rect 9864 410 9916 416
rect 9968 400 9996 954
rect 9128 128 9180 134
rect 9128 70 9180 76
rect 9218 0 9274 400
rect 9312 342 9364 348
rect 9586 0 9642 400
rect 9954 0 10010 400
rect 10060 338 10088 1294
rect 10140 1216 10192 1222
rect 10140 1158 10192 1164
rect 10152 814 10180 1158
rect 10704 882 10732 1414
rect 10888 1290 10916 1414
rect 10966 1391 11022 1400
rect 10784 1284 10836 1290
rect 10784 1226 10836 1232
rect 10876 1284 10928 1290
rect 10876 1226 10928 1232
rect 10692 876 10744 882
rect 10692 818 10744 824
rect 10140 808 10192 814
rect 10140 750 10192 756
rect 10232 672 10284 678
rect 10232 614 10284 620
rect 10244 406 10272 614
rect 10364 572 10740 581
rect 10420 570 10444 572
rect 10500 570 10524 572
rect 10580 570 10604 572
rect 10660 570 10684 572
rect 10420 518 10430 570
rect 10674 518 10684 570
rect 10420 516 10444 518
rect 10500 516 10524 518
rect 10580 516 10604 518
rect 10660 516 10684 518
rect 10364 507 10740 516
rect 10416 468 10468 474
rect 10336 428 10416 456
rect 10232 400 10284 406
rect 10336 400 10364 428
rect 10416 410 10468 416
rect 10600 468 10652 474
rect 10652 428 10732 456
rect 10600 410 10652 416
rect 10704 400 10732 428
rect 10796 406 10824 1226
rect 10968 944 11020 950
rect 10968 886 11020 892
rect 10980 490 11008 886
rect 11072 814 11100 2536
rect 11244 2440 11296 2446
rect 11242 2408 11244 2417
rect 11296 2408 11298 2417
rect 11242 2343 11298 2352
rect 11428 2372 11480 2378
rect 11256 1902 11284 2343
rect 11428 2314 11480 2320
rect 11440 1902 11468 2314
rect 11520 2304 11572 2310
rect 11520 2246 11572 2252
rect 11532 1902 11560 2246
rect 11624 2106 11652 2751
rect 11716 2746 11836 2774
rect 11808 2650 11836 2746
rect 11886 2680 11942 2689
rect 11704 2644 11756 2650
rect 11704 2586 11756 2592
rect 11796 2644 11848 2650
rect 11886 2615 11888 2624
rect 11796 2586 11848 2592
rect 11940 2615 11942 2624
rect 11888 2586 11940 2592
rect 11716 2514 11744 2586
rect 11704 2508 11756 2514
rect 11704 2450 11756 2456
rect 11886 2272 11942 2281
rect 11886 2207 11942 2216
rect 11900 2106 11928 2207
rect 11612 2100 11664 2106
rect 11612 2042 11664 2048
rect 11888 2100 11940 2106
rect 11888 2042 11940 2048
rect 11244 1896 11296 1902
rect 11244 1838 11296 1844
rect 11428 1896 11480 1902
rect 11428 1838 11480 1844
rect 11520 1896 11572 1902
rect 11520 1838 11572 1844
rect 11612 1896 11664 1902
rect 11612 1838 11664 1844
rect 11888 1896 11940 1902
rect 11888 1838 11940 1844
rect 11244 1760 11296 1766
rect 11244 1702 11296 1708
rect 11428 1760 11480 1766
rect 11428 1702 11480 1708
rect 11060 808 11112 814
rect 11060 750 11112 756
rect 11256 728 11284 1702
rect 11336 1420 11388 1426
rect 11336 1362 11388 1368
rect 11348 1018 11376 1362
rect 11336 1012 11388 1018
rect 11336 954 11388 960
rect 11440 950 11468 1702
rect 11520 1216 11572 1222
rect 11520 1158 11572 1164
rect 11532 1018 11560 1158
rect 11520 1012 11572 1018
rect 11520 954 11572 960
rect 11428 944 11480 950
rect 11428 886 11480 892
rect 11336 740 11388 746
rect 11256 700 11336 728
rect 11336 682 11388 688
rect 11520 740 11572 746
rect 11624 728 11652 1838
rect 11704 1420 11756 1426
rect 11704 1362 11756 1368
rect 11716 814 11744 1362
rect 11900 814 11928 1838
rect 11992 1426 12020 3334
rect 12532 3120 12584 3126
rect 12532 3062 12584 3068
rect 12256 3052 12308 3058
rect 12256 2994 12308 3000
rect 12072 2848 12124 2854
rect 12072 2790 12124 2796
rect 12084 1601 12112 2790
rect 12268 2514 12296 2994
rect 12348 2916 12400 2922
rect 12348 2858 12400 2864
rect 12360 2650 12388 2858
rect 12348 2644 12400 2650
rect 12348 2586 12400 2592
rect 12164 2508 12216 2514
rect 12164 2450 12216 2456
rect 12256 2508 12308 2514
rect 12256 2450 12308 2456
rect 12176 2145 12204 2450
rect 12162 2136 12218 2145
rect 12162 2071 12218 2080
rect 12360 1902 12388 2586
rect 12440 2576 12492 2582
rect 12438 2544 12440 2553
rect 12492 2544 12494 2553
rect 12544 2514 12572 3062
rect 12912 2990 12940 3674
rect 12900 2984 12952 2990
rect 12900 2926 12952 2932
rect 12624 2848 12676 2854
rect 12622 2816 12624 2825
rect 12676 2816 12678 2825
rect 12622 2751 12678 2760
rect 12438 2479 12494 2488
rect 12532 2508 12584 2514
rect 12452 2281 12480 2479
rect 12532 2450 12584 2456
rect 12900 2508 12952 2514
rect 12900 2450 12952 2456
rect 12438 2272 12494 2281
rect 12438 2207 12494 2216
rect 12440 1964 12492 1970
rect 12440 1906 12492 1912
rect 12348 1896 12400 1902
rect 12452 1873 12480 1906
rect 12348 1838 12400 1844
rect 12438 1864 12494 1873
rect 12438 1799 12494 1808
rect 12070 1592 12126 1601
rect 12544 1562 12572 2450
rect 12912 2378 12940 2450
rect 12900 2372 12952 2378
rect 12900 2314 12952 2320
rect 12624 2304 12676 2310
rect 12624 2246 12676 2252
rect 12636 1873 12664 2246
rect 12912 1902 12940 2314
rect 12716 1896 12768 1902
rect 12622 1864 12678 1873
rect 12900 1896 12952 1902
rect 12716 1838 12768 1844
rect 12806 1864 12862 1873
rect 12622 1799 12678 1808
rect 12624 1760 12676 1766
rect 12624 1702 12676 1708
rect 12070 1527 12126 1536
rect 12532 1556 12584 1562
rect 12084 1426 12112 1527
rect 12532 1498 12584 1504
rect 11980 1420 12032 1426
rect 11980 1362 12032 1368
rect 12072 1420 12124 1426
rect 12072 1362 12124 1368
rect 11704 808 11756 814
rect 11704 750 11756 756
rect 11888 808 11940 814
rect 11888 750 11940 756
rect 11572 700 11652 728
rect 11520 682 11572 688
rect 11152 672 11204 678
rect 11152 614 11204 620
rect 11428 672 11480 678
rect 11428 614 11480 620
rect 10980 462 11100 490
rect 11164 474 11192 614
rect 10784 400 10836 406
rect 11072 400 11100 462
rect 11152 468 11204 474
rect 11152 410 11204 416
rect 11440 400 11468 614
rect 10232 342 10284 348
rect 10048 332 10100 338
rect 10048 274 10100 280
rect 10060 241 10088 274
rect 10046 232 10102 241
rect 10046 167 10102 176
rect 10322 0 10378 400
rect 10690 0 10746 400
rect 10784 342 10836 348
rect 11058 0 11114 400
rect 11426 0 11482 400
rect 11716 270 11744 750
rect 11796 672 11848 678
rect 11796 614 11848 620
rect 11808 400 11836 614
rect 12084 474 12112 1362
rect 12348 1284 12400 1290
rect 12348 1226 12400 1232
rect 12164 672 12216 678
rect 12164 614 12216 620
rect 12072 468 12124 474
rect 12072 410 12124 416
rect 12176 400 12204 614
rect 11704 264 11756 270
rect 11704 206 11756 212
rect 11794 0 11850 400
rect 12072 128 12124 134
rect 12070 96 12072 105
rect 12124 96 12126 105
rect 12070 31 12126 40
rect 12162 0 12218 400
rect 12360 82 12388 1226
rect 12636 814 12664 1702
rect 12624 808 12676 814
rect 12624 750 12676 756
rect 12728 746 12756 1838
rect 12900 1838 12952 1844
rect 12806 1799 12862 1808
rect 12820 1426 12848 1799
rect 13004 1426 13032 3878
rect 13280 3534 13308 4422
rect 13364 4380 13740 4389
rect 13420 4378 13444 4380
rect 13500 4378 13524 4380
rect 13580 4378 13604 4380
rect 13660 4378 13684 4380
rect 13420 4326 13430 4378
rect 13674 4326 13684 4378
rect 13420 4324 13444 4326
rect 13500 4324 13524 4326
rect 13580 4324 13604 4326
rect 13660 4324 13684 4326
rect 13364 4315 13740 4324
rect 13832 4264 13860 5102
rect 13924 4690 13952 5510
rect 14108 5234 14136 6598
rect 14292 6338 14320 9318
rect 14384 6866 14412 10678
rect 14476 10470 14504 11070
rect 14464 10464 14516 10470
rect 14464 10406 14516 10412
rect 14476 9081 14504 10406
rect 14568 10130 14596 12872
rect 14660 11218 14688 15846
rect 14844 15570 14872 16594
rect 15028 15570 15056 21830
rect 15212 21418 15240 22510
rect 15384 22432 15436 22438
rect 15488 22420 15516 22646
rect 15568 22432 15620 22438
rect 15488 22392 15568 22420
rect 15384 22374 15436 22380
rect 15568 22374 15620 22380
rect 15396 22098 15424 22374
rect 15672 22234 15700 23122
rect 15856 22234 15884 23258
rect 16212 23180 16264 23186
rect 16212 23122 16264 23128
rect 15936 23112 15988 23118
rect 15936 23054 15988 23060
rect 15948 22506 15976 23054
rect 16028 23044 16080 23050
rect 16028 22986 16080 22992
rect 15936 22500 15988 22506
rect 15936 22442 15988 22448
rect 16040 22386 16068 22986
rect 16120 22568 16172 22574
rect 16120 22510 16172 22516
rect 15948 22358 16068 22386
rect 15660 22228 15712 22234
rect 15660 22170 15712 22176
rect 15844 22228 15896 22234
rect 15844 22170 15896 22176
rect 15292 22092 15344 22098
rect 15292 22034 15344 22040
rect 15384 22092 15436 22098
rect 15384 22034 15436 22040
rect 15660 22092 15712 22098
rect 15660 22034 15712 22040
rect 15304 21554 15332 22034
rect 15384 21684 15436 21690
rect 15384 21626 15436 21632
rect 15292 21548 15344 21554
rect 15292 21490 15344 21496
rect 15396 21418 15424 21626
rect 15568 21548 15620 21554
rect 15568 21490 15620 21496
rect 15200 21412 15252 21418
rect 15200 21354 15252 21360
rect 15384 21412 15436 21418
rect 15384 21354 15436 21360
rect 15212 20942 15240 21354
rect 15384 21140 15436 21146
rect 15384 21082 15436 21088
rect 15200 20936 15252 20942
rect 15106 20904 15162 20913
rect 15200 20878 15252 20884
rect 15106 20839 15162 20848
rect 15120 19922 15148 20839
rect 15108 19916 15160 19922
rect 15108 19858 15160 19864
rect 15108 19712 15160 19718
rect 15108 19654 15160 19660
rect 15120 18222 15148 19654
rect 15212 19310 15240 20878
rect 15292 20800 15344 20806
rect 15292 20742 15344 20748
rect 15304 20398 15332 20742
rect 15292 20392 15344 20398
rect 15292 20334 15344 20340
rect 15292 20256 15344 20262
rect 15292 20198 15344 20204
rect 15304 19514 15332 20198
rect 15292 19508 15344 19514
rect 15292 19450 15344 19456
rect 15200 19304 15252 19310
rect 15200 19246 15252 19252
rect 15292 18896 15344 18902
rect 15292 18838 15344 18844
rect 15304 18426 15332 18838
rect 15292 18420 15344 18426
rect 15292 18362 15344 18368
rect 15108 18216 15160 18222
rect 15108 18158 15160 18164
rect 15200 18148 15252 18154
rect 15200 18090 15252 18096
rect 15212 15706 15240 18090
rect 15396 15978 15424 21082
rect 15580 20262 15608 21490
rect 15672 20602 15700 22034
rect 15752 21684 15804 21690
rect 15752 21626 15804 21632
rect 15764 21146 15792 21626
rect 15948 21593 15976 22358
rect 16028 22228 16080 22234
rect 16028 22170 16080 22176
rect 16040 21622 16068 22170
rect 16132 22098 16160 22510
rect 16224 22234 16252 23122
rect 17132 22772 17184 22778
rect 17132 22714 17184 22720
rect 17040 22432 17092 22438
rect 17040 22374 17092 22380
rect 16364 22332 16740 22341
rect 16420 22330 16444 22332
rect 16500 22330 16524 22332
rect 16580 22330 16604 22332
rect 16660 22330 16684 22332
rect 16420 22278 16430 22330
rect 16674 22278 16684 22330
rect 16420 22276 16444 22278
rect 16500 22276 16524 22278
rect 16580 22276 16604 22278
rect 16660 22276 16684 22278
rect 16364 22267 16740 22276
rect 16212 22228 16264 22234
rect 16212 22170 16264 22176
rect 16120 22092 16172 22098
rect 16120 22034 16172 22040
rect 16856 22092 16908 22098
rect 16856 22034 16908 22040
rect 16868 21978 16896 22034
rect 16868 21950 16988 21978
rect 16396 21888 16448 21894
rect 16396 21830 16448 21836
rect 16856 21888 16908 21894
rect 16856 21830 16908 21836
rect 16118 21720 16174 21729
rect 16118 21655 16174 21664
rect 16028 21616 16080 21622
rect 15934 21584 15990 21593
rect 16028 21558 16080 21564
rect 15934 21519 15990 21528
rect 16132 21434 16160 21655
rect 15844 21412 15896 21418
rect 15844 21354 15896 21360
rect 15948 21406 16160 21434
rect 15752 21140 15804 21146
rect 15752 21082 15804 21088
rect 15660 20596 15712 20602
rect 15660 20538 15712 20544
rect 15764 20398 15792 21082
rect 15660 20392 15712 20398
rect 15660 20334 15712 20340
rect 15752 20392 15804 20398
rect 15752 20334 15804 20340
rect 15568 20256 15620 20262
rect 15568 20198 15620 20204
rect 15568 19916 15620 19922
rect 15568 19858 15620 19864
rect 15580 19718 15608 19858
rect 15568 19712 15620 19718
rect 15568 19654 15620 19660
rect 15568 19236 15620 19242
rect 15568 19178 15620 19184
rect 15580 18222 15608 19178
rect 15568 18216 15620 18222
rect 15568 18158 15620 18164
rect 15568 17740 15620 17746
rect 15568 17682 15620 17688
rect 15580 17338 15608 17682
rect 15568 17332 15620 17338
rect 15568 17274 15620 17280
rect 15672 17218 15700 20334
rect 15856 19922 15884 21354
rect 15948 20058 15976 21406
rect 16408 21350 16436 21830
rect 16672 21480 16724 21486
rect 16724 21440 16804 21468
rect 16672 21422 16724 21428
rect 16120 21344 16172 21350
rect 16120 21286 16172 21292
rect 16396 21344 16448 21350
rect 16396 21286 16448 21292
rect 15936 20052 15988 20058
rect 15936 19994 15988 20000
rect 16028 20052 16080 20058
rect 16028 19994 16080 20000
rect 15844 19916 15896 19922
rect 15844 19858 15896 19864
rect 15752 19236 15804 19242
rect 15752 19178 15804 19184
rect 15764 18970 15792 19178
rect 15752 18964 15804 18970
rect 15752 18906 15804 18912
rect 15856 18086 15884 19858
rect 16040 19258 16068 19994
rect 16132 19786 16160 21286
rect 16364 21244 16740 21253
rect 16420 21242 16444 21244
rect 16500 21242 16524 21244
rect 16580 21242 16604 21244
rect 16660 21242 16684 21244
rect 16420 21190 16430 21242
rect 16674 21190 16684 21242
rect 16420 21188 16444 21190
rect 16500 21188 16524 21190
rect 16580 21188 16604 21190
rect 16660 21188 16684 21190
rect 16364 21179 16740 21188
rect 16776 21010 16804 21440
rect 16396 21004 16448 21010
rect 16396 20946 16448 20952
rect 16764 21004 16816 21010
rect 16764 20946 16816 20952
rect 16408 20602 16436 20946
rect 16396 20596 16448 20602
rect 16396 20538 16448 20544
rect 16210 20496 16266 20505
rect 16210 20431 16212 20440
rect 16264 20431 16266 20440
rect 16212 20402 16264 20408
rect 16364 20156 16740 20165
rect 16420 20154 16444 20156
rect 16500 20154 16524 20156
rect 16580 20154 16604 20156
rect 16660 20154 16684 20156
rect 16420 20102 16430 20154
rect 16674 20102 16684 20154
rect 16420 20100 16444 20102
rect 16500 20100 16524 20102
rect 16580 20100 16604 20102
rect 16660 20100 16684 20102
rect 16364 20091 16740 20100
rect 16776 19922 16804 20946
rect 16868 20534 16896 21830
rect 16960 21350 16988 21950
rect 16948 21344 17000 21350
rect 16948 21286 17000 21292
rect 16856 20528 16908 20534
rect 16856 20470 16908 20476
rect 16948 20460 17000 20466
rect 16948 20402 17000 20408
rect 16856 20392 16908 20398
rect 16854 20360 16856 20369
rect 16908 20360 16910 20369
rect 16854 20295 16910 20304
rect 16960 20058 16988 20402
rect 17052 20330 17080 22374
rect 17144 22030 17172 22714
rect 17236 22234 17264 23598
rect 17972 23050 18000 23666
rect 18234 23600 18290 24000
rect 18786 23600 18842 24000
rect 19338 23746 19394 24000
rect 19338 23718 19840 23746
rect 19338 23600 19394 23718
rect 18248 23254 18276 23600
rect 18800 23254 18828 23600
rect 18236 23248 18288 23254
rect 18236 23190 18288 23196
rect 18788 23248 18840 23254
rect 18788 23190 18840 23196
rect 18696 23112 18748 23118
rect 18696 23054 18748 23060
rect 17960 23044 18012 23050
rect 17960 22986 18012 22992
rect 17972 22642 18000 22986
rect 17316 22636 17368 22642
rect 17316 22578 17368 22584
rect 17960 22636 18012 22642
rect 17960 22578 18012 22584
rect 17224 22228 17276 22234
rect 17224 22170 17276 22176
rect 17328 22030 17356 22578
rect 17960 22160 18012 22166
rect 17960 22102 18012 22108
rect 17868 22092 17920 22098
rect 17868 22034 17920 22040
rect 17132 22024 17184 22030
rect 17132 21966 17184 21972
rect 17316 22024 17368 22030
rect 17316 21966 17368 21972
rect 17222 20632 17278 20641
rect 17328 20602 17356 21966
rect 17776 21412 17828 21418
rect 17776 21354 17828 21360
rect 17500 21344 17552 21350
rect 17500 21286 17552 21292
rect 17512 20874 17540 21286
rect 17592 21072 17644 21078
rect 17592 21014 17644 21020
rect 17604 20942 17632 21014
rect 17592 20936 17644 20942
rect 17592 20878 17644 20884
rect 17500 20868 17552 20874
rect 17500 20810 17552 20816
rect 17222 20567 17278 20576
rect 17316 20596 17368 20602
rect 17236 20534 17264 20567
rect 17316 20538 17368 20544
rect 17224 20528 17276 20534
rect 17224 20470 17276 20476
rect 17040 20324 17092 20330
rect 17040 20266 17092 20272
rect 17604 20058 17632 20878
rect 16948 20052 17000 20058
rect 16948 19994 17000 20000
rect 17592 20052 17644 20058
rect 17592 19994 17644 20000
rect 16764 19916 16816 19922
rect 16764 19858 16816 19864
rect 16120 19780 16172 19786
rect 16120 19722 16172 19728
rect 16212 19712 16264 19718
rect 16212 19654 16264 19660
rect 16304 19712 16356 19718
rect 16304 19654 16356 19660
rect 16580 19712 16632 19718
rect 16580 19654 16632 19660
rect 15948 19230 16068 19258
rect 16120 19304 16172 19310
rect 16120 19246 16172 19252
rect 15948 18766 15976 19230
rect 15936 18760 15988 18766
rect 15936 18702 15988 18708
rect 16132 18290 16160 19246
rect 16224 19224 16252 19654
rect 16316 19417 16344 19654
rect 16302 19408 16358 19417
rect 16302 19343 16358 19352
rect 16488 19236 16540 19242
rect 16224 19196 16488 19224
rect 16488 19178 16540 19184
rect 16592 19174 16620 19654
rect 16580 19168 16632 19174
rect 16580 19110 16632 19116
rect 16364 19068 16740 19077
rect 16420 19066 16444 19068
rect 16500 19066 16524 19068
rect 16580 19066 16604 19068
rect 16660 19066 16684 19068
rect 16420 19014 16430 19066
rect 16674 19014 16684 19066
rect 16420 19012 16444 19014
rect 16500 19012 16524 19014
rect 16580 19012 16604 19014
rect 16660 19012 16684 19014
rect 16364 19003 16740 19012
rect 16120 18284 16172 18290
rect 16120 18226 16172 18232
rect 15752 18080 15804 18086
rect 15752 18022 15804 18028
rect 15844 18080 15896 18086
rect 15844 18022 15896 18028
rect 15764 17746 15792 18022
rect 16364 17980 16740 17989
rect 16420 17978 16444 17980
rect 16500 17978 16524 17980
rect 16580 17978 16604 17980
rect 16660 17978 16684 17980
rect 16420 17926 16430 17978
rect 16674 17926 16684 17978
rect 16420 17924 16444 17926
rect 16500 17924 16524 17926
rect 16580 17924 16604 17926
rect 16660 17924 16684 17926
rect 16364 17915 16740 17924
rect 15842 17776 15898 17785
rect 15752 17740 15804 17746
rect 15898 17720 15976 17728
rect 15842 17711 15844 17720
rect 15752 17682 15804 17688
rect 15896 17700 15976 17720
rect 15844 17682 15896 17688
rect 15672 17190 15884 17218
rect 15476 17128 15528 17134
rect 15476 17070 15528 17076
rect 15752 17128 15804 17134
rect 15752 17070 15804 17076
rect 15488 16794 15516 17070
rect 15568 16992 15620 16998
rect 15764 16969 15792 17070
rect 15568 16934 15620 16940
rect 15750 16960 15806 16969
rect 15476 16788 15528 16794
rect 15476 16730 15528 16736
rect 15580 16658 15608 16934
rect 15750 16895 15806 16904
rect 15568 16652 15620 16658
rect 15568 16594 15620 16600
rect 15660 16244 15712 16250
rect 15660 16186 15712 16192
rect 15384 15972 15436 15978
rect 15384 15914 15436 15920
rect 15672 15881 15700 16186
rect 15658 15872 15714 15881
rect 15658 15807 15714 15816
rect 15200 15700 15252 15706
rect 15200 15642 15252 15648
rect 15672 15570 15700 15807
rect 15764 15570 15792 16895
rect 14832 15564 14884 15570
rect 14832 15506 14884 15512
rect 15016 15564 15068 15570
rect 15016 15506 15068 15512
rect 15660 15564 15712 15570
rect 15660 15506 15712 15512
rect 15752 15564 15804 15570
rect 15752 15506 15804 15512
rect 14844 14958 14872 15506
rect 14924 15428 14976 15434
rect 14924 15370 14976 15376
rect 15108 15428 15160 15434
rect 15108 15370 15160 15376
rect 15476 15428 15528 15434
rect 15476 15370 15528 15376
rect 14832 14952 14884 14958
rect 14832 14894 14884 14900
rect 14740 14544 14792 14550
rect 14740 14486 14792 14492
rect 14752 13870 14780 14486
rect 14936 14414 14964 15370
rect 15016 15360 15068 15366
rect 15016 15302 15068 15308
rect 15028 15026 15056 15302
rect 15016 15020 15068 15026
rect 15016 14962 15068 14968
rect 15028 14482 15056 14962
rect 15120 14958 15148 15370
rect 15292 15156 15344 15162
rect 15292 15098 15344 15104
rect 15108 14952 15160 14958
rect 15108 14894 15160 14900
rect 15108 14816 15160 14822
rect 15108 14758 15160 14764
rect 15016 14476 15068 14482
rect 15016 14418 15068 14424
rect 14924 14408 14976 14414
rect 15120 14362 15148 14758
rect 14924 14350 14976 14356
rect 15028 14334 15148 14362
rect 15198 14376 15254 14385
rect 14832 14272 14884 14278
rect 14832 14214 14884 14220
rect 14740 13864 14792 13870
rect 14740 13806 14792 13812
rect 14752 13326 14780 13806
rect 14740 13320 14792 13326
rect 14740 13262 14792 13268
rect 14844 12374 14872 14214
rect 15028 13274 15056 14334
rect 15198 14311 15254 14320
rect 15108 14272 15160 14278
rect 15108 14214 15160 14220
rect 15120 13870 15148 14214
rect 15108 13864 15160 13870
rect 15108 13806 15160 13812
rect 15108 13728 15160 13734
rect 15108 13670 15160 13676
rect 15120 13394 15148 13670
rect 15108 13388 15160 13394
rect 15108 13330 15160 13336
rect 15212 13326 15240 14311
rect 15304 13870 15332 15098
rect 15488 14074 15516 15370
rect 15856 14278 15884 17190
rect 15948 16998 15976 17700
rect 16028 17536 16080 17542
rect 16028 17478 16080 17484
rect 15936 16992 15988 16998
rect 15936 16934 15988 16940
rect 15948 16658 15976 16934
rect 15936 16652 15988 16658
rect 15936 16594 15988 16600
rect 15936 16448 15988 16454
rect 15936 16390 15988 16396
rect 15844 14272 15896 14278
rect 15844 14214 15896 14220
rect 15476 14068 15528 14074
rect 15476 14010 15528 14016
rect 15488 13870 15516 14010
rect 15842 13968 15898 13977
rect 15842 13903 15898 13912
rect 15292 13864 15344 13870
rect 15292 13806 15344 13812
rect 15476 13864 15528 13870
rect 15476 13806 15528 13812
rect 15304 13462 15332 13806
rect 15750 13696 15806 13705
rect 15750 13631 15806 13640
rect 15292 13456 15344 13462
rect 15292 13398 15344 13404
rect 15200 13320 15252 13326
rect 15028 13258 15148 13274
rect 15200 13262 15252 13268
rect 15028 13252 15160 13258
rect 15028 13246 15108 13252
rect 15108 13194 15160 13200
rect 14924 13184 14976 13190
rect 14924 13126 14976 13132
rect 15200 13184 15252 13190
rect 15200 13126 15252 13132
rect 14832 12368 14884 12374
rect 14832 12310 14884 12316
rect 14740 12096 14792 12102
rect 14740 12038 14792 12044
rect 14648 11212 14700 11218
rect 14648 11154 14700 11160
rect 14752 10674 14780 12038
rect 14844 11694 14872 12310
rect 14832 11688 14884 11694
rect 14832 11630 14884 11636
rect 14832 11552 14884 11558
rect 14832 11494 14884 11500
rect 14740 10668 14792 10674
rect 14740 10610 14792 10616
rect 14844 10577 14872 11494
rect 14936 11218 14964 13126
rect 15108 12912 15160 12918
rect 15108 12854 15160 12860
rect 15016 12844 15068 12850
rect 15016 12786 15068 12792
rect 15028 12306 15056 12786
rect 15016 12300 15068 12306
rect 15016 12242 15068 12248
rect 15016 12096 15068 12102
rect 15016 12038 15068 12044
rect 15028 11762 15056 12038
rect 15016 11756 15068 11762
rect 15016 11698 15068 11704
rect 14924 11212 14976 11218
rect 14924 11154 14976 11160
rect 15120 10674 15148 12854
rect 15212 12714 15240 13126
rect 15384 12776 15436 12782
rect 15384 12718 15436 12724
rect 15476 12776 15528 12782
rect 15476 12718 15528 12724
rect 15200 12708 15252 12714
rect 15200 12650 15252 12656
rect 15292 12708 15344 12714
rect 15292 12650 15344 12656
rect 15200 12436 15252 12442
rect 15200 12378 15252 12384
rect 15212 11762 15240 12378
rect 15304 12306 15332 12650
rect 15396 12442 15424 12718
rect 15488 12481 15516 12718
rect 15474 12472 15530 12481
rect 15384 12436 15436 12442
rect 15764 12442 15792 13631
rect 15474 12407 15530 12416
rect 15752 12436 15804 12442
rect 15384 12378 15436 12384
rect 15752 12378 15804 12384
rect 15292 12300 15344 12306
rect 15292 12242 15344 12248
rect 15660 12164 15712 12170
rect 15660 12106 15712 12112
rect 15476 12096 15528 12102
rect 15382 12064 15438 12073
rect 15476 12038 15528 12044
rect 15382 11999 15438 12008
rect 15200 11756 15252 11762
rect 15200 11698 15252 11704
rect 15212 11150 15240 11698
rect 15396 11336 15424 11999
rect 15488 11762 15516 12038
rect 15476 11756 15528 11762
rect 15476 11698 15528 11704
rect 15568 11756 15620 11762
rect 15568 11698 15620 11704
rect 15580 11642 15608 11698
rect 15488 11626 15608 11642
rect 15476 11620 15608 11626
rect 15528 11614 15608 11620
rect 15476 11562 15528 11568
rect 15568 11552 15620 11558
rect 15568 11494 15620 11500
rect 15396 11308 15516 11336
rect 15382 11248 15438 11257
rect 15382 11183 15384 11192
rect 15436 11183 15438 11192
rect 15384 11154 15436 11160
rect 15200 11144 15252 11150
rect 15200 11086 15252 11092
rect 15292 11008 15344 11014
rect 15292 10950 15344 10956
rect 15200 10804 15252 10810
rect 15200 10746 15252 10752
rect 15108 10668 15160 10674
rect 15108 10610 15160 10616
rect 14830 10568 14886 10577
rect 14830 10503 14886 10512
rect 15108 10532 15160 10538
rect 14646 10432 14702 10441
rect 14646 10367 14702 10376
rect 14556 10124 14608 10130
rect 14556 10066 14608 10072
rect 14660 9722 14688 10367
rect 14844 10062 14872 10503
rect 15108 10474 15160 10480
rect 14832 10056 14884 10062
rect 14832 9998 14884 10004
rect 14924 10056 14976 10062
rect 14924 9998 14976 10004
rect 14830 9888 14886 9897
rect 14830 9823 14886 9832
rect 14648 9716 14700 9722
rect 14648 9658 14700 9664
rect 14740 9648 14792 9654
rect 14740 9590 14792 9596
rect 14752 9518 14780 9590
rect 14740 9512 14792 9518
rect 14740 9454 14792 9460
rect 14648 9444 14700 9450
rect 14648 9386 14700 9392
rect 14462 9072 14518 9081
rect 14462 9007 14518 9016
rect 14660 8838 14688 9386
rect 14752 9042 14780 9454
rect 14740 9036 14792 9042
rect 14740 8978 14792 8984
rect 14556 8832 14608 8838
rect 14556 8774 14608 8780
rect 14648 8832 14700 8838
rect 14648 8774 14700 8780
rect 14568 8294 14596 8774
rect 14844 8650 14872 9823
rect 14660 8622 14872 8650
rect 14464 8288 14516 8294
rect 14464 8230 14516 8236
rect 14556 8288 14608 8294
rect 14556 8230 14608 8236
rect 14476 7410 14504 8230
rect 14556 7744 14608 7750
rect 14554 7712 14556 7721
rect 14608 7712 14610 7721
rect 14554 7647 14610 7656
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 14476 6866 14504 7346
rect 14660 7206 14688 8622
rect 14936 8537 14964 9998
rect 15016 9988 15068 9994
rect 15016 9930 15068 9936
rect 15028 9654 15056 9930
rect 15016 9648 15068 9654
rect 15016 9590 15068 9596
rect 15120 9353 15148 10474
rect 15106 9344 15162 9353
rect 15106 9279 15162 9288
rect 15106 9072 15162 9081
rect 15016 9036 15068 9042
rect 15106 9007 15108 9016
rect 15016 8978 15068 8984
rect 15160 9007 15162 9016
rect 15108 8978 15160 8984
rect 14922 8528 14978 8537
rect 14922 8463 14978 8472
rect 15028 8362 15056 8978
rect 15108 8832 15160 8838
rect 15106 8800 15108 8809
rect 15160 8800 15162 8809
rect 15106 8735 15162 8744
rect 15106 8528 15162 8537
rect 15106 8463 15162 8472
rect 15120 8430 15148 8463
rect 15108 8424 15160 8430
rect 15108 8366 15160 8372
rect 15016 8356 15068 8362
rect 15016 8298 15068 8304
rect 14832 8288 14884 8294
rect 14832 8230 14884 8236
rect 14844 7886 14872 8230
rect 14832 7880 14884 7886
rect 14832 7822 14884 7828
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect 14832 7744 14884 7750
rect 14832 7686 14884 7692
rect 14752 7478 14780 7686
rect 14740 7472 14792 7478
rect 14740 7414 14792 7420
rect 14648 7200 14700 7206
rect 14648 7142 14700 7148
rect 14740 6996 14792 7002
rect 14740 6938 14792 6944
rect 14372 6860 14424 6866
rect 14372 6802 14424 6808
rect 14464 6860 14516 6866
rect 14464 6802 14516 6808
rect 14648 6860 14700 6866
rect 14648 6802 14700 6808
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14200 6310 14320 6338
rect 14200 6254 14228 6310
rect 14188 6248 14240 6254
rect 14188 6190 14240 6196
rect 14372 6248 14424 6254
rect 14372 6190 14424 6196
rect 14096 5228 14148 5234
rect 14096 5170 14148 5176
rect 14004 5160 14056 5166
rect 14004 5102 14056 5108
rect 14016 4826 14044 5102
rect 14004 4820 14056 4826
rect 14004 4762 14056 4768
rect 13912 4684 13964 4690
rect 13912 4626 13964 4632
rect 13740 4236 13860 4264
rect 13740 4078 13768 4236
rect 13728 4072 13780 4078
rect 13728 4014 13780 4020
rect 13820 4072 13872 4078
rect 13924 4060 13952 4626
rect 14004 4480 14056 4486
rect 14004 4422 14056 4428
rect 14016 4146 14044 4422
rect 14108 4214 14136 5170
rect 14200 5166 14228 6190
rect 14384 5778 14412 6190
rect 14372 5772 14424 5778
rect 14372 5714 14424 5720
rect 14372 5636 14424 5642
rect 14372 5578 14424 5584
rect 14188 5160 14240 5166
rect 14188 5102 14240 5108
rect 14384 5030 14412 5578
rect 14464 5568 14516 5574
rect 14464 5510 14516 5516
rect 14476 5234 14504 5510
rect 14464 5228 14516 5234
rect 14464 5170 14516 5176
rect 14372 5024 14424 5030
rect 14372 4966 14424 4972
rect 14476 4826 14504 5170
rect 14464 4820 14516 4826
rect 14464 4762 14516 4768
rect 14186 4312 14242 4321
rect 14186 4247 14188 4256
rect 14240 4247 14242 4256
rect 14188 4218 14240 4224
rect 14096 4208 14148 4214
rect 14096 4150 14148 4156
rect 14004 4140 14056 4146
rect 14004 4082 14056 4088
rect 14200 4078 14228 4218
rect 14464 4208 14516 4214
rect 14464 4150 14516 4156
rect 14476 4078 14504 4150
rect 13872 4032 13952 4060
rect 14188 4072 14240 4078
rect 13820 4014 13872 4020
rect 14188 4014 14240 4020
rect 14464 4072 14516 4078
rect 14464 4014 14516 4020
rect 13820 3936 13872 3942
rect 13820 3878 13872 3884
rect 13832 3602 13860 3878
rect 14094 3632 14150 3641
rect 13820 3596 13872 3602
rect 14094 3567 14096 3576
rect 13820 3538 13872 3544
rect 14148 3567 14150 3576
rect 14096 3538 14148 3544
rect 13268 3528 13320 3534
rect 13268 3470 13320 3476
rect 13820 3392 13872 3398
rect 13820 3334 13872 3340
rect 13364 3292 13740 3301
rect 13420 3290 13444 3292
rect 13500 3290 13524 3292
rect 13580 3290 13604 3292
rect 13660 3290 13684 3292
rect 13420 3238 13430 3290
rect 13674 3238 13684 3290
rect 13420 3236 13444 3238
rect 13500 3236 13524 3238
rect 13580 3236 13604 3238
rect 13660 3236 13684 3238
rect 13364 3227 13740 3236
rect 13452 3120 13504 3126
rect 13452 3062 13504 3068
rect 13084 2508 13136 2514
rect 13084 2450 13136 2456
rect 13464 2496 13492 3062
rect 13728 2984 13780 2990
rect 13728 2926 13780 2932
rect 13544 2916 13596 2922
rect 13544 2858 13596 2864
rect 13556 2650 13584 2858
rect 13740 2825 13768 2926
rect 13726 2816 13782 2825
rect 13726 2751 13782 2760
rect 13544 2644 13596 2650
rect 13544 2586 13596 2592
rect 13832 2514 13860 3334
rect 14108 2990 14136 3538
rect 14188 3392 14240 3398
rect 14188 3334 14240 3340
rect 14096 2984 14148 2990
rect 14094 2952 14096 2961
rect 14148 2952 14150 2961
rect 14094 2887 14150 2896
rect 13544 2508 13596 2514
rect 13464 2468 13544 2496
rect 13096 2145 13124 2450
rect 13464 2428 13492 2468
rect 13544 2450 13596 2456
rect 13728 2508 13780 2514
rect 13728 2450 13780 2456
rect 13820 2508 13872 2514
rect 13820 2450 13872 2456
rect 13280 2400 13492 2428
rect 13082 2136 13138 2145
rect 13280 2106 13308 2400
rect 13740 2394 13768 2450
rect 14200 2417 14228 3334
rect 14476 2990 14504 4014
rect 14464 2984 14516 2990
rect 14464 2926 14516 2932
rect 14568 2514 14596 6598
rect 14660 6254 14688 6802
rect 14752 6390 14780 6938
rect 14740 6384 14792 6390
rect 14740 6326 14792 6332
rect 14648 6248 14700 6254
rect 14648 6190 14700 6196
rect 14648 6112 14700 6118
rect 14648 6054 14700 6060
rect 14660 5914 14688 6054
rect 14648 5908 14700 5914
rect 14648 5850 14700 5856
rect 14740 5704 14792 5710
rect 14740 5646 14792 5652
rect 14752 5166 14780 5646
rect 14740 5160 14792 5166
rect 14740 5102 14792 5108
rect 14648 5024 14700 5030
rect 14648 4966 14700 4972
rect 14660 4826 14688 4966
rect 14648 4820 14700 4826
rect 14648 4762 14700 4768
rect 14844 4622 14872 7686
rect 14924 7336 14976 7342
rect 14924 7278 14976 7284
rect 14936 6662 14964 7278
rect 15028 7206 15056 8298
rect 15108 7812 15160 7818
rect 15108 7754 15160 7760
rect 15016 7200 15068 7206
rect 15016 7142 15068 7148
rect 15016 6792 15068 6798
rect 15016 6734 15068 6740
rect 14924 6656 14976 6662
rect 14924 6598 14976 6604
rect 14936 6322 14964 6598
rect 15028 6458 15056 6734
rect 15016 6452 15068 6458
rect 15016 6394 15068 6400
rect 15120 6322 15148 7754
rect 15212 6866 15240 10746
rect 15304 10674 15332 10950
rect 15292 10668 15344 10674
rect 15292 10610 15344 10616
rect 15292 10532 15344 10538
rect 15292 10474 15344 10480
rect 15304 10130 15332 10474
rect 15292 10124 15344 10130
rect 15292 10066 15344 10072
rect 15292 9988 15344 9994
rect 15292 9930 15344 9936
rect 15304 9761 15332 9930
rect 15290 9752 15346 9761
rect 15290 9687 15346 9696
rect 15290 9208 15346 9217
rect 15290 9143 15346 9152
rect 15304 8362 15332 9143
rect 15292 8356 15344 8362
rect 15292 8298 15344 8304
rect 15304 8090 15332 8298
rect 15292 8084 15344 8090
rect 15292 8026 15344 8032
rect 15292 7744 15344 7750
rect 15292 7686 15344 7692
rect 15304 6866 15332 7686
rect 15396 7041 15424 11154
rect 15488 10198 15516 11308
rect 15476 10192 15528 10198
rect 15476 10134 15528 10140
rect 15488 8566 15516 10134
rect 15476 8560 15528 8566
rect 15476 8502 15528 8508
rect 15474 8392 15530 8401
rect 15474 8327 15530 8336
rect 15488 7342 15516 8327
rect 15580 7585 15608 11494
rect 15672 11218 15700 12106
rect 15752 11688 15804 11694
rect 15752 11630 15804 11636
rect 15764 11286 15792 11630
rect 15856 11370 15884 13903
rect 15948 13870 15976 16390
rect 16040 15745 16068 17478
rect 16672 17332 16724 17338
rect 16672 17274 16724 17280
rect 16684 17202 16712 17274
rect 16776 17270 16804 19858
rect 16856 19168 16908 19174
rect 16856 19110 16908 19116
rect 16868 18970 16896 19110
rect 16856 18964 16908 18970
rect 16856 18906 16908 18912
rect 16960 18834 16988 19994
rect 17040 19984 17092 19990
rect 17040 19926 17092 19932
rect 17052 18970 17080 19926
rect 17314 19816 17370 19825
rect 17314 19751 17370 19760
rect 17040 18964 17092 18970
rect 17040 18906 17092 18912
rect 17328 18834 17356 19751
rect 17592 19712 17644 19718
rect 17592 19654 17644 19660
rect 17604 18834 17632 19654
rect 17684 19168 17736 19174
rect 17684 19110 17736 19116
rect 16948 18828 17000 18834
rect 16948 18770 17000 18776
rect 17316 18828 17368 18834
rect 17592 18828 17644 18834
rect 17316 18770 17368 18776
rect 17512 18788 17592 18816
rect 16948 18624 17000 18630
rect 16948 18566 17000 18572
rect 16856 18284 16908 18290
rect 16856 18226 16908 18232
rect 16764 17264 16816 17270
rect 16764 17206 16816 17212
rect 16672 17196 16724 17202
rect 16672 17138 16724 17144
rect 16684 17054 16804 17082
rect 16684 16998 16712 17054
rect 16672 16992 16724 16998
rect 16672 16934 16724 16940
rect 16364 16892 16740 16901
rect 16420 16890 16444 16892
rect 16500 16890 16524 16892
rect 16580 16890 16604 16892
rect 16660 16890 16684 16892
rect 16420 16838 16430 16890
rect 16674 16838 16684 16890
rect 16420 16836 16444 16838
rect 16500 16836 16524 16838
rect 16580 16836 16604 16838
rect 16660 16836 16684 16838
rect 16364 16827 16740 16836
rect 16776 16726 16804 17054
rect 16868 16998 16896 18226
rect 16960 17882 16988 18566
rect 17512 18222 17540 18788
rect 17592 18770 17644 18776
rect 17592 18624 17644 18630
rect 17592 18566 17644 18572
rect 17604 18426 17632 18566
rect 17592 18420 17644 18426
rect 17592 18362 17644 18368
rect 17040 18216 17092 18222
rect 17040 18158 17092 18164
rect 17500 18216 17552 18222
rect 17500 18158 17552 18164
rect 16948 17876 17000 17882
rect 16948 17818 17000 17824
rect 17052 17814 17080 18158
rect 17316 18148 17368 18154
rect 17316 18090 17368 18096
rect 17040 17808 17092 17814
rect 17040 17750 17092 17756
rect 16948 17740 17000 17746
rect 16948 17682 17000 17688
rect 16960 17338 16988 17682
rect 16948 17332 17000 17338
rect 16948 17274 17000 17280
rect 16856 16992 16908 16998
rect 16856 16934 16908 16940
rect 16764 16720 16816 16726
rect 16764 16662 16816 16668
rect 16212 16652 16264 16658
rect 16212 16594 16264 16600
rect 16224 16250 16252 16594
rect 16212 16244 16264 16250
rect 16212 16186 16264 16192
rect 16120 15972 16172 15978
rect 16120 15914 16172 15920
rect 16026 15736 16082 15745
rect 16026 15671 16082 15680
rect 16132 15502 16160 15914
rect 16212 15904 16264 15910
rect 16212 15846 16264 15852
rect 16224 15638 16252 15846
rect 16364 15804 16740 15813
rect 16420 15802 16444 15804
rect 16500 15802 16524 15804
rect 16580 15802 16604 15804
rect 16660 15802 16684 15804
rect 16420 15750 16430 15802
rect 16674 15750 16684 15802
rect 16420 15748 16444 15750
rect 16500 15748 16524 15750
rect 16580 15748 16604 15750
rect 16660 15748 16684 15750
rect 16364 15739 16740 15748
rect 16212 15632 16264 15638
rect 16212 15574 16264 15580
rect 16120 15496 16172 15502
rect 16120 15438 16172 15444
rect 16488 15360 16540 15366
rect 16488 15302 16540 15308
rect 16764 15360 16816 15366
rect 16764 15302 16816 15308
rect 16500 15094 16528 15302
rect 16488 15088 16540 15094
rect 16488 15030 16540 15036
rect 16040 14878 16344 14906
rect 15936 13864 15988 13870
rect 15936 13806 15988 13812
rect 16040 12646 16068 14878
rect 16316 14822 16344 14878
rect 16212 14816 16264 14822
rect 16212 14758 16264 14764
rect 16304 14816 16356 14822
rect 16304 14758 16356 14764
rect 16120 13932 16172 13938
rect 16120 13874 16172 13880
rect 16028 12640 16080 12646
rect 16028 12582 16080 12588
rect 15936 12368 15988 12374
rect 15936 12310 15988 12316
rect 15948 11830 15976 12310
rect 16028 12096 16080 12102
rect 16028 12038 16080 12044
rect 15936 11824 15988 11830
rect 15936 11766 15988 11772
rect 15856 11342 15976 11370
rect 15752 11280 15804 11286
rect 15804 11240 15884 11268
rect 15752 11222 15804 11228
rect 15660 11212 15712 11218
rect 15660 11154 15712 11160
rect 15752 11144 15804 11150
rect 15752 11086 15804 11092
rect 15764 10674 15792 11086
rect 15856 10810 15884 11240
rect 15844 10804 15896 10810
rect 15844 10746 15896 10752
rect 15752 10668 15804 10674
rect 15752 10610 15804 10616
rect 15660 10600 15712 10606
rect 15856 10554 15884 10746
rect 15660 10542 15712 10548
rect 15672 10418 15700 10542
rect 15764 10538 15884 10554
rect 15752 10532 15884 10538
rect 15804 10526 15884 10532
rect 15752 10474 15804 10480
rect 15672 10390 15884 10418
rect 15856 10266 15884 10390
rect 15844 10260 15896 10266
rect 15844 10202 15896 10208
rect 15752 10192 15804 10198
rect 15752 10134 15804 10140
rect 15660 9444 15712 9450
rect 15660 9386 15712 9392
rect 15672 8673 15700 9386
rect 15764 8974 15792 10134
rect 15948 10010 15976 11342
rect 15856 9982 15976 10010
rect 15856 9586 15884 9982
rect 15934 9752 15990 9761
rect 15934 9687 15990 9696
rect 15844 9580 15896 9586
rect 15844 9522 15896 9528
rect 15856 9042 15884 9522
rect 15844 9036 15896 9042
rect 15844 8978 15896 8984
rect 15752 8968 15804 8974
rect 15752 8910 15804 8916
rect 15658 8664 15714 8673
rect 15658 8599 15714 8608
rect 15752 8560 15804 8566
rect 15752 8502 15804 8508
rect 15660 7948 15712 7954
rect 15660 7890 15712 7896
rect 15672 7818 15700 7890
rect 15660 7812 15712 7818
rect 15660 7754 15712 7760
rect 15566 7576 15622 7585
rect 15566 7511 15622 7520
rect 15476 7336 15528 7342
rect 15476 7278 15528 7284
rect 15566 7168 15622 7177
rect 15566 7103 15622 7112
rect 15382 7032 15438 7041
rect 15382 6967 15438 6976
rect 15200 6860 15252 6866
rect 15200 6802 15252 6808
rect 15292 6860 15344 6866
rect 15292 6802 15344 6808
rect 15384 6860 15436 6866
rect 15384 6802 15436 6808
rect 15476 6860 15528 6866
rect 15476 6802 15528 6808
rect 15292 6724 15344 6730
rect 15292 6666 15344 6672
rect 14924 6316 14976 6322
rect 14924 6258 14976 6264
rect 15108 6316 15160 6322
rect 15108 6258 15160 6264
rect 15120 5914 15148 6258
rect 15200 6248 15252 6254
rect 15200 6190 15252 6196
rect 15212 6089 15240 6190
rect 15198 6080 15254 6089
rect 15198 6015 15254 6024
rect 15108 5908 15160 5914
rect 15108 5850 15160 5856
rect 15200 5568 15252 5574
rect 15200 5510 15252 5516
rect 14922 4856 14978 4865
rect 14922 4791 14978 4800
rect 14832 4616 14884 4622
rect 14832 4558 14884 4564
rect 14740 4140 14792 4146
rect 14740 4082 14792 4088
rect 14752 3738 14780 4082
rect 14844 3738 14872 4558
rect 14936 4486 14964 4791
rect 14924 4480 14976 4486
rect 14924 4422 14976 4428
rect 14936 4282 14964 4422
rect 14924 4276 14976 4282
rect 14924 4218 14976 4224
rect 15212 4146 15240 5510
rect 15304 4146 15332 6666
rect 15396 6089 15424 6802
rect 15488 6662 15516 6802
rect 15580 6712 15608 7103
rect 15672 6934 15700 7754
rect 15764 7750 15792 8502
rect 15844 8492 15896 8498
rect 15844 8434 15896 8440
rect 15856 7750 15884 8434
rect 15752 7744 15804 7750
rect 15752 7686 15804 7692
rect 15844 7744 15896 7750
rect 15844 7686 15896 7692
rect 15856 7546 15884 7686
rect 15844 7540 15896 7546
rect 15844 7482 15896 7488
rect 15660 6928 15712 6934
rect 15660 6870 15712 6876
rect 15580 6684 15700 6712
rect 15476 6656 15528 6662
rect 15476 6598 15528 6604
rect 15382 6080 15438 6089
rect 15382 6015 15438 6024
rect 15488 4758 15516 6598
rect 15568 6248 15620 6254
rect 15568 6190 15620 6196
rect 15580 5710 15608 6190
rect 15568 5704 15620 5710
rect 15568 5646 15620 5652
rect 15476 4752 15528 4758
rect 15476 4694 15528 4700
rect 15384 4548 15436 4554
rect 15384 4490 15436 4496
rect 15396 4146 15424 4490
rect 15672 4146 15700 6684
rect 15752 6656 15804 6662
rect 15752 6598 15804 6604
rect 15764 4185 15792 6598
rect 15948 6322 15976 9687
rect 16040 8922 16068 12038
rect 16132 10520 16160 13874
rect 16224 13870 16252 14758
rect 16364 14716 16740 14725
rect 16420 14714 16444 14716
rect 16500 14714 16524 14716
rect 16580 14714 16604 14716
rect 16660 14714 16684 14716
rect 16420 14662 16430 14714
rect 16674 14662 16684 14714
rect 16420 14660 16444 14662
rect 16500 14660 16524 14662
rect 16580 14660 16604 14662
rect 16660 14660 16684 14662
rect 16364 14651 16740 14660
rect 16776 14346 16804 15302
rect 16764 14340 16816 14346
rect 16764 14282 16816 14288
rect 16396 13932 16448 13938
rect 16396 13874 16448 13880
rect 16212 13864 16264 13870
rect 16212 13806 16264 13812
rect 16408 13734 16436 13874
rect 16868 13870 16896 16934
rect 17052 16776 17080 17750
rect 17224 16992 17276 16998
rect 17224 16934 17276 16940
rect 16960 16748 17080 16776
rect 16960 16046 16988 16748
rect 17132 16720 17184 16726
rect 17132 16662 17184 16668
rect 17040 16652 17092 16658
rect 17040 16594 17092 16600
rect 16948 16040 17000 16046
rect 16948 15982 17000 15988
rect 16948 14000 17000 14006
rect 16948 13942 17000 13948
rect 16856 13864 16908 13870
rect 16856 13806 16908 13812
rect 16212 13728 16264 13734
rect 16212 13670 16264 13676
rect 16396 13728 16448 13734
rect 16396 13670 16448 13676
rect 16764 13728 16816 13734
rect 16764 13670 16816 13676
rect 16224 10674 16252 13670
rect 16364 13628 16740 13637
rect 16420 13626 16444 13628
rect 16500 13626 16524 13628
rect 16580 13626 16604 13628
rect 16660 13626 16684 13628
rect 16420 13574 16430 13626
rect 16674 13574 16684 13626
rect 16420 13572 16444 13574
rect 16500 13572 16524 13574
rect 16580 13572 16604 13574
rect 16660 13572 16684 13574
rect 16364 13563 16740 13572
rect 16580 13524 16632 13530
rect 16580 13466 16632 13472
rect 16592 12764 16620 13466
rect 16776 13444 16804 13670
rect 16684 13416 16804 13444
rect 16684 13326 16712 13416
rect 16672 13320 16724 13326
rect 16672 13262 16724 13268
rect 16960 12782 16988 13942
rect 17052 13530 17080 16594
rect 17144 15586 17172 16662
rect 17236 16658 17264 16934
rect 17224 16652 17276 16658
rect 17224 16594 17276 16600
rect 17144 15558 17264 15586
rect 17132 15496 17184 15502
rect 17132 15438 17184 15444
rect 17144 14958 17172 15438
rect 17132 14952 17184 14958
rect 17132 14894 17184 14900
rect 17132 14340 17184 14346
rect 17132 14282 17184 14288
rect 17144 13938 17172 14282
rect 17132 13932 17184 13938
rect 17132 13874 17184 13880
rect 17040 13524 17092 13530
rect 17040 13466 17092 13472
rect 17052 13394 17080 13466
rect 17040 13388 17092 13394
rect 17040 13330 17092 13336
rect 17132 13184 17184 13190
rect 17052 13144 17132 13172
rect 16856 12776 16908 12782
rect 16592 12736 16804 12764
rect 16364 12540 16740 12549
rect 16420 12538 16444 12540
rect 16500 12538 16524 12540
rect 16580 12538 16604 12540
rect 16660 12538 16684 12540
rect 16420 12486 16430 12538
rect 16674 12486 16684 12538
rect 16420 12484 16444 12486
rect 16500 12484 16524 12486
rect 16580 12484 16604 12486
rect 16660 12484 16684 12486
rect 16364 12475 16740 12484
rect 16304 12436 16356 12442
rect 16356 12406 16528 12434
rect 16304 12378 16356 12384
rect 16500 12374 16528 12406
rect 16488 12368 16540 12374
rect 16488 12310 16540 12316
rect 16304 12300 16356 12306
rect 16304 12242 16356 12248
rect 16396 12300 16448 12306
rect 16396 12242 16448 12248
rect 16316 11898 16344 12242
rect 16408 12102 16436 12242
rect 16670 12200 16726 12209
rect 16670 12135 16726 12144
rect 16396 12096 16448 12102
rect 16396 12038 16448 12044
rect 16304 11892 16356 11898
rect 16304 11834 16356 11840
rect 16684 11694 16712 12135
rect 16580 11688 16632 11694
rect 16578 11656 16580 11665
rect 16672 11688 16724 11694
rect 16632 11656 16634 11665
rect 16672 11630 16724 11636
rect 16578 11591 16634 11600
rect 16364 11452 16740 11461
rect 16420 11450 16444 11452
rect 16500 11450 16524 11452
rect 16580 11450 16604 11452
rect 16660 11450 16684 11452
rect 16420 11398 16430 11450
rect 16674 11398 16684 11450
rect 16420 11396 16444 11398
rect 16500 11396 16524 11398
rect 16580 11396 16604 11398
rect 16660 11396 16684 11398
rect 16364 11387 16740 11396
rect 16302 11248 16358 11257
rect 16302 11183 16304 11192
rect 16356 11183 16358 11192
rect 16304 11154 16356 11160
rect 16776 10810 16804 12736
rect 16856 12718 16908 12724
rect 16948 12776 17000 12782
rect 16948 12718 17000 12724
rect 16868 12424 16896 12718
rect 16868 12396 16988 12424
rect 16856 12300 16908 12306
rect 16856 12242 16908 12248
rect 16868 11898 16896 12242
rect 16960 11898 16988 12396
rect 16856 11892 16908 11898
rect 16856 11834 16908 11840
rect 16948 11892 17000 11898
rect 16948 11834 17000 11840
rect 16948 11620 17000 11626
rect 16948 11562 17000 11568
rect 16856 11348 16908 11354
rect 16856 11290 16908 11296
rect 16764 10804 16816 10810
rect 16764 10746 16816 10752
rect 16212 10668 16264 10674
rect 16212 10610 16264 10616
rect 16672 10668 16724 10674
rect 16724 10628 16804 10656
rect 16672 10610 16724 10616
rect 16212 10532 16264 10538
rect 16132 10492 16212 10520
rect 16212 10474 16264 10480
rect 16396 10464 16448 10470
rect 16309 10424 16396 10452
rect 16309 10418 16337 10424
rect 16224 10390 16337 10418
rect 16396 10406 16448 10412
rect 16118 10160 16174 10169
rect 16118 10095 16120 10104
rect 16172 10095 16174 10104
rect 16120 10066 16172 10072
rect 16040 8894 16160 8922
rect 16028 8832 16080 8838
rect 16028 8774 16080 8780
rect 16040 8430 16068 8774
rect 16028 8424 16080 8430
rect 16028 8366 16080 8372
rect 16026 8120 16082 8129
rect 16026 8055 16082 8064
rect 16040 7954 16068 8055
rect 16028 7948 16080 7954
rect 16028 7890 16080 7896
rect 15936 6316 15988 6322
rect 15936 6258 15988 6264
rect 15844 6248 15896 6254
rect 15844 6190 15896 6196
rect 15856 5914 15884 6190
rect 15936 6112 15988 6118
rect 15936 6054 15988 6060
rect 15844 5908 15896 5914
rect 15844 5850 15896 5856
rect 15750 4176 15806 4185
rect 15200 4140 15252 4146
rect 15200 4082 15252 4088
rect 15292 4140 15344 4146
rect 15292 4082 15344 4088
rect 15384 4140 15436 4146
rect 15384 4082 15436 4088
rect 15660 4140 15712 4146
rect 15750 4111 15806 4120
rect 15660 4082 15712 4088
rect 14924 3936 14976 3942
rect 14924 3878 14976 3884
rect 15108 3936 15160 3942
rect 15108 3878 15160 3884
rect 14740 3732 14792 3738
rect 14740 3674 14792 3680
rect 14832 3732 14884 3738
rect 14832 3674 14884 3680
rect 14556 2508 14608 2514
rect 14556 2450 14608 2456
rect 14186 2408 14242 2417
rect 13740 2366 14136 2394
rect 14108 2310 14136 2366
rect 14186 2343 14242 2352
rect 14004 2304 14056 2310
rect 14004 2246 14056 2252
rect 14096 2304 14148 2310
rect 14096 2246 14148 2252
rect 14278 2272 14334 2281
rect 13364 2204 13740 2213
rect 13420 2202 13444 2204
rect 13500 2202 13524 2204
rect 13580 2202 13604 2204
rect 13660 2202 13684 2204
rect 13420 2150 13430 2202
rect 13674 2150 13684 2202
rect 13420 2148 13444 2150
rect 13500 2148 13524 2150
rect 13580 2148 13604 2150
rect 13660 2148 13684 2150
rect 13364 2139 13740 2148
rect 13818 2136 13874 2145
rect 13082 2071 13138 2080
rect 13268 2100 13320 2106
rect 13268 2042 13320 2048
rect 13648 2080 13818 2088
rect 13648 2071 13874 2080
rect 13648 2060 13860 2071
rect 13268 1828 13320 1834
rect 13268 1770 13320 1776
rect 13084 1760 13136 1766
rect 13084 1702 13136 1708
rect 13176 1760 13228 1766
rect 13176 1702 13228 1708
rect 13096 1562 13124 1702
rect 13084 1556 13136 1562
rect 13084 1498 13136 1504
rect 12808 1420 12860 1426
rect 12808 1362 12860 1368
rect 12992 1420 13044 1426
rect 12992 1362 13044 1368
rect 13084 1420 13136 1426
rect 13084 1362 13136 1368
rect 13096 1222 13124 1362
rect 13084 1216 13136 1222
rect 13084 1158 13136 1164
rect 13188 882 13216 1702
rect 13176 876 13228 882
rect 13176 818 13228 824
rect 13280 814 13308 1770
rect 13648 1766 13676 2060
rect 14016 2038 14044 2246
rect 14108 2106 14136 2246
rect 14278 2207 14334 2216
rect 14096 2100 14148 2106
rect 14096 2042 14148 2048
rect 14004 2032 14056 2038
rect 14004 1974 14056 1980
rect 14292 1970 14320 2207
rect 14280 1964 14332 1970
rect 14280 1906 14332 1912
rect 14372 1964 14424 1970
rect 14372 1906 14424 1912
rect 13728 1828 13780 1834
rect 13728 1770 13780 1776
rect 13636 1760 13688 1766
rect 13636 1702 13688 1708
rect 13358 1456 13414 1465
rect 13648 1426 13676 1702
rect 13740 1426 13768 1770
rect 14384 1494 14412 1906
rect 14464 1896 14516 1902
rect 14464 1838 14516 1844
rect 14554 1864 14610 1873
rect 14372 1488 14424 1494
rect 14372 1430 14424 1436
rect 13358 1391 13414 1400
rect 13636 1420 13688 1426
rect 13372 1358 13400 1391
rect 13636 1362 13688 1368
rect 13728 1420 13780 1426
rect 13728 1362 13780 1368
rect 13360 1352 13412 1358
rect 13360 1294 13412 1300
rect 14280 1284 14332 1290
rect 14280 1226 14332 1232
rect 13820 1216 13872 1222
rect 13820 1158 13872 1164
rect 13364 1116 13740 1125
rect 13420 1114 13444 1116
rect 13500 1114 13524 1116
rect 13580 1114 13604 1116
rect 13660 1114 13684 1116
rect 13420 1062 13430 1114
rect 13674 1062 13684 1114
rect 13420 1060 13444 1062
rect 13500 1060 13524 1062
rect 13580 1060 13604 1062
rect 13660 1060 13684 1062
rect 13364 1051 13740 1060
rect 13832 814 13860 1158
rect 14186 1048 14242 1057
rect 14186 983 14188 992
rect 14240 983 14242 992
rect 14188 954 14240 960
rect 13268 808 13320 814
rect 13268 750 13320 756
rect 13820 808 13872 814
rect 13820 750 13872 756
rect 12716 740 12768 746
rect 12716 682 12768 688
rect 12532 672 12584 678
rect 12532 614 12584 620
rect 12900 672 12952 678
rect 12900 614 12952 620
rect 13268 672 13320 678
rect 13728 672 13780 678
rect 13268 614 13320 620
rect 13648 632 13728 660
rect 12544 400 12572 614
rect 12912 400 12940 614
rect 12992 400 13044 406
rect 13280 400 13308 614
rect 13648 400 13676 632
rect 14096 672 14148 678
rect 13728 614 13780 620
rect 14016 632 14096 660
rect 14016 400 14044 632
rect 14096 614 14148 620
rect 12268 66 12388 82
rect 12256 60 12388 66
rect 12308 54 12388 60
rect 12256 2 12308 8
rect 12530 0 12586 400
rect 12898 0 12954 400
rect 12992 342 13044 348
rect 13004 202 13032 342
rect 12992 196 13044 202
rect 12992 138 13044 144
rect 13266 0 13322 400
rect 13634 0 13690 400
rect 14002 0 14058 400
rect 14292 338 14320 1226
rect 14384 882 14412 1430
rect 14476 1290 14504 1838
rect 14554 1799 14610 1808
rect 14568 1426 14596 1799
rect 14648 1760 14700 1766
rect 14648 1702 14700 1708
rect 14556 1420 14608 1426
rect 14556 1362 14608 1368
rect 14464 1284 14516 1290
rect 14464 1226 14516 1232
rect 14372 876 14424 882
rect 14372 818 14424 824
rect 14476 814 14504 1226
rect 14568 1193 14596 1362
rect 14554 1184 14610 1193
rect 14554 1119 14610 1128
rect 14660 814 14688 1702
rect 14936 1494 14964 3878
rect 15016 2848 15068 2854
rect 15016 2790 15068 2796
rect 15028 2514 15056 2790
rect 15016 2508 15068 2514
rect 15016 2450 15068 2456
rect 15014 1728 15070 1737
rect 15014 1663 15070 1672
rect 14924 1488 14976 1494
rect 14924 1430 14976 1436
rect 15028 1306 15056 1663
rect 15120 1426 15148 3878
rect 15396 3534 15424 4082
rect 15844 4072 15896 4078
rect 15844 4014 15896 4020
rect 15660 3936 15712 3942
rect 15660 3878 15712 3884
rect 15672 3670 15700 3878
rect 15660 3664 15712 3670
rect 15660 3606 15712 3612
rect 15856 3534 15884 4014
rect 15948 3602 15976 6054
rect 16028 5092 16080 5098
rect 16028 5034 16080 5040
rect 16040 4298 16068 5034
rect 16132 4690 16160 8894
rect 16224 6322 16252 10390
rect 16364 10364 16740 10373
rect 16420 10362 16444 10364
rect 16500 10362 16524 10364
rect 16580 10362 16604 10364
rect 16660 10362 16684 10364
rect 16420 10310 16430 10362
rect 16674 10310 16684 10362
rect 16420 10308 16444 10310
rect 16500 10308 16524 10310
rect 16580 10308 16604 10310
rect 16660 10308 16684 10310
rect 16364 10299 16740 10308
rect 16304 10124 16356 10130
rect 16304 10066 16356 10072
rect 16316 9586 16344 10066
rect 16394 10024 16450 10033
rect 16394 9959 16396 9968
rect 16448 9959 16450 9968
rect 16396 9930 16448 9936
rect 16776 9761 16804 10628
rect 16762 9752 16818 9761
rect 16762 9687 16818 9696
rect 16394 9616 16450 9625
rect 16304 9580 16356 9586
rect 16394 9551 16396 9560
rect 16304 9522 16356 9528
rect 16448 9551 16450 9560
rect 16762 9616 16818 9625
rect 16762 9551 16818 9560
rect 16396 9522 16448 9528
rect 16672 9512 16724 9518
rect 16670 9480 16672 9489
rect 16724 9480 16726 9489
rect 16670 9415 16726 9424
rect 16364 9276 16740 9285
rect 16420 9274 16444 9276
rect 16500 9274 16524 9276
rect 16580 9274 16604 9276
rect 16660 9274 16684 9276
rect 16420 9222 16430 9274
rect 16674 9222 16684 9274
rect 16420 9220 16444 9222
rect 16500 9220 16524 9222
rect 16580 9220 16604 9222
rect 16660 9220 16684 9222
rect 16364 9211 16740 9220
rect 16776 9024 16804 9551
rect 16684 8996 16804 9024
rect 16304 8968 16356 8974
rect 16304 8910 16356 8916
rect 16580 8968 16632 8974
rect 16580 8910 16632 8916
rect 16316 8430 16344 8910
rect 16592 8430 16620 8910
rect 16684 8906 16712 8996
rect 16868 8922 16896 11290
rect 16960 10985 16988 11562
rect 16946 10976 17002 10985
rect 16946 10911 17002 10920
rect 16948 10804 17000 10810
rect 16948 10746 17000 10752
rect 16960 10606 16988 10746
rect 16948 10600 17000 10606
rect 16948 10542 17000 10548
rect 16672 8900 16724 8906
rect 16672 8842 16724 8848
rect 16776 8894 16896 8922
rect 16776 8566 16804 8894
rect 16856 8832 16908 8838
rect 16856 8774 16908 8780
rect 16764 8560 16816 8566
rect 16764 8502 16816 8508
rect 16868 8430 16896 8774
rect 16304 8424 16356 8430
rect 16304 8366 16356 8372
rect 16580 8424 16632 8430
rect 16580 8366 16632 8372
rect 16856 8424 16908 8430
rect 16856 8366 16908 8372
rect 16764 8356 16816 8362
rect 16764 8298 16816 8304
rect 16364 8188 16740 8197
rect 16420 8186 16444 8188
rect 16500 8186 16524 8188
rect 16580 8186 16604 8188
rect 16660 8186 16684 8188
rect 16420 8134 16430 8186
rect 16674 8134 16684 8186
rect 16420 8132 16444 8134
rect 16500 8132 16524 8134
rect 16580 8132 16604 8134
rect 16660 8132 16684 8134
rect 16364 8123 16740 8132
rect 16672 7540 16724 7546
rect 16672 7482 16724 7488
rect 16684 7342 16712 7482
rect 16672 7336 16724 7342
rect 16672 7278 16724 7284
rect 16364 7100 16740 7109
rect 16420 7098 16444 7100
rect 16500 7098 16524 7100
rect 16580 7098 16604 7100
rect 16660 7098 16684 7100
rect 16420 7046 16430 7098
rect 16674 7046 16684 7098
rect 16420 7044 16444 7046
rect 16500 7044 16524 7046
rect 16580 7044 16604 7046
rect 16660 7044 16684 7046
rect 16364 7035 16740 7044
rect 16776 6798 16804 8298
rect 16856 7200 16908 7206
rect 16856 7142 16908 7148
rect 16764 6792 16816 6798
rect 16764 6734 16816 6740
rect 16488 6724 16540 6730
rect 16488 6666 16540 6672
rect 16212 6316 16264 6322
rect 16212 6258 16264 6264
rect 16500 6254 16528 6666
rect 16304 6248 16356 6254
rect 16302 6216 16304 6225
rect 16488 6248 16540 6254
rect 16356 6216 16358 6225
rect 16488 6190 16540 6196
rect 16302 6151 16358 6160
rect 16364 6012 16740 6021
rect 16420 6010 16444 6012
rect 16500 6010 16524 6012
rect 16580 6010 16604 6012
rect 16660 6010 16684 6012
rect 16420 5958 16430 6010
rect 16674 5958 16684 6010
rect 16420 5956 16444 5958
rect 16500 5956 16524 5958
rect 16580 5956 16604 5958
rect 16660 5956 16684 5958
rect 16364 5947 16740 5956
rect 16868 5846 16896 7142
rect 16580 5840 16632 5846
rect 16580 5782 16632 5788
rect 16856 5840 16908 5846
rect 16856 5782 16908 5788
rect 16592 5234 16620 5782
rect 16580 5228 16632 5234
rect 16580 5170 16632 5176
rect 16672 5228 16724 5234
rect 16960 5216 16988 10542
rect 17052 10470 17080 13144
rect 17132 13126 17184 13132
rect 17236 12918 17264 15558
rect 17328 14618 17356 18090
rect 17408 17060 17460 17066
rect 17408 17002 17460 17008
rect 17420 16658 17448 17002
rect 17408 16652 17460 16658
rect 17408 16594 17460 16600
rect 17500 16448 17552 16454
rect 17500 16390 17552 16396
rect 17408 15972 17460 15978
rect 17408 15914 17460 15920
rect 17420 15638 17448 15914
rect 17408 15632 17460 15638
rect 17408 15574 17460 15580
rect 17420 15502 17448 15574
rect 17408 15496 17460 15502
rect 17408 15438 17460 15444
rect 17408 14816 17460 14822
rect 17408 14758 17460 14764
rect 17316 14612 17368 14618
rect 17316 14554 17368 14560
rect 17224 12912 17276 12918
rect 17224 12854 17276 12860
rect 17132 12640 17184 12646
rect 17132 12582 17184 12588
rect 17144 12306 17172 12582
rect 17132 12300 17184 12306
rect 17132 12242 17184 12248
rect 17328 12186 17356 14554
rect 17236 12158 17356 12186
rect 17132 11688 17184 11694
rect 17132 11630 17184 11636
rect 17144 11286 17172 11630
rect 17132 11280 17184 11286
rect 17132 11222 17184 11228
rect 17130 10976 17186 10985
rect 17130 10911 17186 10920
rect 17040 10464 17092 10470
rect 17040 10406 17092 10412
rect 17040 9376 17092 9382
rect 17040 9318 17092 9324
rect 17052 7886 17080 9318
rect 17144 9110 17172 10911
rect 17132 9104 17184 9110
rect 17130 9072 17132 9081
rect 17184 9072 17186 9081
rect 17130 9007 17186 9016
rect 17236 8974 17264 12158
rect 17316 12096 17368 12102
rect 17316 12038 17368 12044
rect 17328 11354 17356 12038
rect 17420 11642 17448 14758
rect 17512 13394 17540 16390
rect 17604 16017 17632 18362
rect 17696 17066 17724 19110
rect 17788 18970 17816 21354
rect 17880 21026 17908 22034
rect 17972 21729 18000 22102
rect 18708 22098 18736 23054
rect 18880 22976 18932 22982
rect 18880 22918 18932 22924
rect 18604 22092 18656 22098
rect 18604 22034 18656 22040
rect 18696 22092 18748 22098
rect 18696 22034 18748 22040
rect 17958 21720 18014 21729
rect 17958 21655 18014 21664
rect 18420 21344 18472 21350
rect 18420 21286 18472 21292
rect 17880 20998 18092 21026
rect 17868 20936 17920 20942
rect 17868 20878 17920 20884
rect 17880 20602 17908 20878
rect 17868 20596 17920 20602
rect 18064 20584 18092 20998
rect 18144 20596 18196 20602
rect 18064 20556 18144 20584
rect 17868 20538 17920 20544
rect 18432 20584 18460 21286
rect 18616 21078 18644 22034
rect 18604 21072 18656 21078
rect 18604 21014 18656 21020
rect 18708 20874 18736 22034
rect 18892 21876 18920 22918
rect 19364 22876 19740 22885
rect 19420 22874 19444 22876
rect 19500 22874 19524 22876
rect 19580 22874 19604 22876
rect 19660 22874 19684 22876
rect 19420 22822 19430 22874
rect 19674 22822 19684 22874
rect 19420 22820 19444 22822
rect 19500 22820 19524 22822
rect 19580 22820 19604 22822
rect 19660 22820 19684 22822
rect 19364 22811 19740 22820
rect 19708 22772 19760 22778
rect 19708 22714 19760 22720
rect 19064 22704 19116 22710
rect 19064 22646 19116 22652
rect 18972 22024 19024 22030
rect 19076 22012 19104 22646
rect 19720 22438 19748 22714
rect 19812 22710 19840 23718
rect 19890 23600 19946 24000
rect 20442 23746 20498 24000
rect 20272 23718 20498 23746
rect 19800 22704 19852 22710
rect 19800 22646 19852 22652
rect 19340 22432 19392 22438
rect 19340 22374 19392 22380
rect 19708 22432 19760 22438
rect 19708 22374 19760 22380
rect 19246 22128 19302 22137
rect 19156 22092 19208 22098
rect 19246 22063 19302 22072
rect 19156 22034 19208 22040
rect 19024 21984 19104 22012
rect 18972 21966 19024 21972
rect 18892 21848 19012 21876
rect 18880 21344 18932 21350
rect 18880 21286 18932 21292
rect 18892 21049 18920 21286
rect 18878 21040 18934 21049
rect 18800 20998 18878 21026
rect 18696 20868 18748 20874
rect 18696 20810 18748 20816
rect 18144 20538 18196 20544
rect 18340 20556 18460 20584
rect 17960 20256 18012 20262
rect 17960 20198 18012 20204
rect 17868 19304 17920 19310
rect 17868 19246 17920 19252
rect 17776 18964 17828 18970
rect 17776 18906 17828 18912
rect 17880 18630 17908 19246
rect 17972 18970 18000 20198
rect 18144 19712 18196 19718
rect 18144 19654 18196 19660
rect 18156 19378 18184 19654
rect 18144 19372 18196 19378
rect 18144 19314 18196 19320
rect 17960 18964 18012 18970
rect 17960 18906 18012 18912
rect 18340 18902 18368 20556
rect 18512 20392 18564 20398
rect 18512 20334 18564 20340
rect 18524 19310 18552 20334
rect 18696 20324 18748 20330
rect 18696 20266 18748 20272
rect 18708 19990 18736 20266
rect 18696 19984 18748 19990
rect 18602 19952 18658 19961
rect 18696 19926 18748 19932
rect 18602 19887 18658 19896
rect 18616 19802 18644 19887
rect 18616 19786 18736 19802
rect 18616 19780 18748 19786
rect 18616 19774 18696 19780
rect 18696 19722 18748 19728
rect 18708 19689 18736 19722
rect 18694 19680 18750 19689
rect 18694 19615 18750 19624
rect 18800 19360 18828 20998
rect 18878 20975 18934 20984
rect 18880 20324 18932 20330
rect 18880 20266 18932 20272
rect 18616 19332 18828 19360
rect 18512 19304 18564 19310
rect 18512 19246 18564 19252
rect 18328 18896 18380 18902
rect 18328 18838 18380 18844
rect 17868 18624 17920 18630
rect 17868 18566 17920 18572
rect 18420 18420 18472 18426
rect 18420 18362 18472 18368
rect 18052 18284 18104 18290
rect 18052 18226 18104 18232
rect 17960 18148 18012 18154
rect 17960 18090 18012 18096
rect 17972 17882 18000 18090
rect 17960 17876 18012 17882
rect 17960 17818 18012 17824
rect 17776 17604 17828 17610
rect 17776 17546 17828 17552
rect 17684 17060 17736 17066
rect 17684 17002 17736 17008
rect 17590 16008 17646 16017
rect 17590 15943 17646 15952
rect 17592 15700 17644 15706
rect 17592 15642 17644 15648
rect 17604 14464 17632 15642
rect 17684 15020 17736 15026
rect 17684 14962 17736 14968
rect 17696 14618 17724 14962
rect 17788 14940 17816 17546
rect 17960 17536 18012 17542
rect 17960 17478 18012 17484
rect 17972 16182 18000 17478
rect 18064 17338 18092 18226
rect 18432 18086 18460 18362
rect 18512 18216 18564 18222
rect 18512 18158 18564 18164
rect 18420 18080 18472 18086
rect 18420 18022 18472 18028
rect 18144 17808 18196 17814
rect 18144 17750 18196 17756
rect 18052 17332 18104 17338
rect 18052 17274 18104 17280
rect 18064 17134 18092 17274
rect 18052 17128 18104 17134
rect 18052 17070 18104 17076
rect 17960 16176 18012 16182
rect 17960 16118 18012 16124
rect 17868 15904 17920 15910
rect 17868 15846 17920 15852
rect 17880 15570 17908 15846
rect 18052 15700 18104 15706
rect 18052 15642 18104 15648
rect 17868 15564 17920 15570
rect 17868 15506 17920 15512
rect 17788 14912 17908 14940
rect 17684 14612 17736 14618
rect 17684 14554 17736 14560
rect 17684 14476 17736 14482
rect 17604 14436 17684 14464
rect 17500 13388 17552 13394
rect 17500 13330 17552 13336
rect 17604 13190 17632 14436
rect 17684 14418 17736 14424
rect 17776 13932 17828 13938
rect 17776 13874 17828 13880
rect 17684 13728 17736 13734
rect 17684 13670 17736 13676
rect 17696 13394 17724 13670
rect 17788 13394 17816 13874
rect 17684 13388 17736 13394
rect 17684 13330 17736 13336
rect 17776 13388 17828 13394
rect 17776 13330 17828 13336
rect 17592 13184 17644 13190
rect 17592 13126 17644 13132
rect 17592 12640 17644 12646
rect 17592 12582 17644 12588
rect 17604 12442 17632 12582
rect 17592 12436 17644 12442
rect 17592 12378 17644 12384
rect 17498 12064 17554 12073
rect 17498 11999 17554 12008
rect 17512 11762 17540 11999
rect 17592 11892 17644 11898
rect 17592 11834 17644 11840
rect 17500 11756 17552 11762
rect 17500 11698 17552 11704
rect 17420 11614 17540 11642
rect 17408 11552 17460 11558
rect 17408 11494 17460 11500
rect 17316 11348 17368 11354
rect 17316 11290 17368 11296
rect 17316 11212 17368 11218
rect 17316 11154 17368 11160
rect 17328 10606 17356 11154
rect 17316 10600 17368 10606
rect 17316 10542 17368 10548
rect 17316 10464 17368 10470
rect 17316 10406 17368 10412
rect 17328 9518 17356 10406
rect 17316 9512 17368 9518
rect 17316 9454 17368 9460
rect 17314 9208 17370 9217
rect 17314 9143 17370 9152
rect 17224 8968 17276 8974
rect 17224 8910 17276 8916
rect 17132 8560 17184 8566
rect 17132 8502 17184 8508
rect 17144 8430 17172 8502
rect 17132 8424 17184 8430
rect 17132 8366 17184 8372
rect 17040 7880 17092 7886
rect 17040 7822 17092 7828
rect 17144 7546 17172 8366
rect 17224 7948 17276 7954
rect 17224 7890 17276 7896
rect 17132 7540 17184 7546
rect 17132 7482 17184 7488
rect 17236 7002 17264 7890
rect 17224 6996 17276 7002
rect 17224 6938 17276 6944
rect 17328 6866 17356 9143
rect 17420 6866 17448 11494
rect 17512 10606 17540 11614
rect 17604 10810 17632 11834
rect 17592 10804 17644 10810
rect 17592 10746 17644 10752
rect 17590 10704 17646 10713
rect 17590 10639 17646 10648
rect 17604 10606 17632 10639
rect 17696 10606 17724 13330
rect 17776 12436 17828 12442
rect 17776 12378 17828 12384
rect 17788 12102 17816 12378
rect 17776 12096 17828 12102
rect 17776 12038 17828 12044
rect 17776 11756 17828 11762
rect 17776 11698 17828 11704
rect 17788 11354 17816 11698
rect 17776 11348 17828 11354
rect 17776 11290 17828 11296
rect 17880 11218 17908 14912
rect 18064 12345 18092 15642
rect 18156 14958 18184 17750
rect 18524 17542 18552 18158
rect 18512 17536 18564 17542
rect 18512 17478 18564 17484
rect 18420 17264 18472 17270
rect 18420 17206 18472 17212
rect 18432 17134 18460 17206
rect 18328 17128 18380 17134
rect 18328 17070 18380 17076
rect 18420 17128 18472 17134
rect 18420 17070 18472 17076
rect 18340 16998 18368 17070
rect 18328 16992 18380 16998
rect 18328 16934 18380 16940
rect 18432 16794 18460 17070
rect 18420 16788 18472 16794
rect 18420 16730 18472 16736
rect 18328 16516 18380 16522
rect 18328 16458 18380 16464
rect 18512 16516 18564 16522
rect 18512 16458 18564 16464
rect 18236 16244 18288 16250
rect 18236 16186 18288 16192
rect 18248 15502 18276 16186
rect 18236 15496 18288 15502
rect 18236 15438 18288 15444
rect 18144 14952 18196 14958
rect 18144 14894 18196 14900
rect 18236 13864 18288 13870
rect 18236 13806 18288 13812
rect 18050 12336 18106 12345
rect 18050 12271 18052 12280
rect 18104 12271 18106 12280
rect 18052 12242 18104 12248
rect 18144 12096 18196 12102
rect 18144 12038 18196 12044
rect 18156 11762 18184 12038
rect 18144 11756 18196 11762
rect 18144 11698 18196 11704
rect 18142 11656 18198 11665
rect 18052 11620 18104 11626
rect 18142 11591 18198 11600
rect 18052 11562 18104 11568
rect 17868 11212 17920 11218
rect 17868 11154 17920 11160
rect 17776 11144 17828 11150
rect 17960 11144 18012 11150
rect 17776 11086 17828 11092
rect 17880 11092 17960 11098
rect 17880 11086 18012 11092
rect 17788 10849 17816 11086
rect 17880 11070 18000 11086
rect 17774 10840 17830 10849
rect 17774 10775 17830 10784
rect 17776 10668 17828 10674
rect 17880 10656 17908 11070
rect 17828 10628 17908 10656
rect 17776 10610 17828 10616
rect 17500 10600 17552 10606
rect 17500 10542 17552 10548
rect 17592 10600 17644 10606
rect 17592 10542 17644 10548
rect 17684 10600 17736 10606
rect 17684 10542 17736 10548
rect 17960 10464 18012 10470
rect 17960 10406 18012 10412
rect 17774 10296 17830 10305
rect 17972 10266 18000 10406
rect 17774 10231 17830 10240
rect 17960 10260 18012 10266
rect 17500 9988 17552 9994
rect 17500 9930 17552 9936
rect 17512 8129 17540 9930
rect 17592 9512 17644 9518
rect 17592 9454 17644 9460
rect 17604 9110 17632 9454
rect 17684 9376 17736 9382
rect 17684 9318 17736 9324
rect 17696 9217 17724 9318
rect 17682 9208 17738 9217
rect 17788 9178 17816 10231
rect 17960 10202 18012 10208
rect 17868 9512 17920 9518
rect 17866 9480 17868 9489
rect 17920 9480 17922 9489
rect 17866 9415 17922 9424
rect 17682 9143 17738 9152
rect 17776 9172 17828 9178
rect 17776 9114 17828 9120
rect 17592 9104 17644 9110
rect 17592 9046 17644 9052
rect 17880 9024 17908 9415
rect 17788 8996 17908 9024
rect 17590 8664 17646 8673
rect 17590 8599 17646 8608
rect 17604 8498 17632 8599
rect 17592 8492 17644 8498
rect 17592 8434 17644 8440
rect 17592 8356 17644 8362
rect 17592 8298 17644 8304
rect 17498 8120 17554 8129
rect 17498 8055 17554 8064
rect 17498 7304 17554 7313
rect 17498 7239 17554 7248
rect 17512 6866 17540 7239
rect 17040 6860 17092 6866
rect 17040 6802 17092 6808
rect 17316 6860 17368 6866
rect 17316 6802 17368 6808
rect 17408 6860 17460 6866
rect 17408 6802 17460 6808
rect 17500 6860 17552 6866
rect 17500 6802 17552 6808
rect 17052 5234 17080 6802
rect 17132 6112 17184 6118
rect 17132 6054 17184 6060
rect 17144 5642 17172 6054
rect 17132 5636 17184 5642
rect 17132 5578 17184 5584
rect 17224 5568 17276 5574
rect 17224 5510 17276 5516
rect 17316 5568 17368 5574
rect 17316 5510 17368 5516
rect 16724 5188 16988 5216
rect 17040 5228 17092 5234
rect 16672 5170 16724 5176
rect 17040 5170 17092 5176
rect 16212 5024 16264 5030
rect 16212 4966 16264 4972
rect 16120 4684 16172 4690
rect 16120 4626 16172 4632
rect 16224 4486 16252 4966
rect 16364 4924 16740 4933
rect 16420 4922 16444 4924
rect 16500 4922 16524 4924
rect 16580 4922 16604 4924
rect 16660 4922 16684 4924
rect 16420 4870 16430 4922
rect 16674 4870 16684 4922
rect 16420 4868 16444 4870
rect 16500 4868 16524 4870
rect 16580 4868 16604 4870
rect 16660 4868 16684 4870
rect 16364 4859 16740 4868
rect 17236 4690 17264 5510
rect 17224 4684 17276 4690
rect 17224 4626 17276 4632
rect 16212 4480 16264 4486
rect 16212 4422 16264 4428
rect 17040 4480 17092 4486
rect 17040 4422 17092 4428
rect 16040 4270 16436 4298
rect 16302 4176 16358 4185
rect 16408 4146 16436 4270
rect 16302 4111 16304 4120
rect 16356 4111 16358 4120
rect 16396 4140 16448 4146
rect 16304 4082 16356 4088
rect 16396 4082 16448 4088
rect 16856 4140 16908 4146
rect 16856 4082 16908 4088
rect 16120 4072 16172 4078
rect 16120 4014 16172 4020
rect 16132 3738 16160 4014
rect 16764 3936 16816 3942
rect 16764 3878 16816 3884
rect 16364 3836 16740 3845
rect 16420 3834 16444 3836
rect 16500 3834 16524 3836
rect 16580 3834 16604 3836
rect 16660 3834 16684 3836
rect 16420 3782 16430 3834
rect 16674 3782 16684 3834
rect 16420 3780 16444 3782
rect 16500 3780 16524 3782
rect 16580 3780 16604 3782
rect 16660 3780 16684 3782
rect 16364 3771 16740 3780
rect 16120 3732 16172 3738
rect 16120 3674 16172 3680
rect 16672 3732 16724 3738
rect 16672 3674 16724 3680
rect 16684 3602 16712 3674
rect 15936 3596 15988 3602
rect 15936 3538 15988 3544
rect 16672 3596 16724 3602
rect 16672 3538 16724 3544
rect 15384 3528 15436 3534
rect 15384 3470 15436 3476
rect 15844 3528 15896 3534
rect 15844 3470 15896 3476
rect 15200 3392 15252 3398
rect 15200 3334 15252 3340
rect 15844 3392 15896 3398
rect 15844 3334 15896 3340
rect 15212 3126 15240 3334
rect 15200 3120 15252 3126
rect 15200 3062 15252 3068
rect 15198 2544 15254 2553
rect 15198 2479 15200 2488
rect 15252 2479 15254 2488
rect 15384 2508 15436 2514
rect 15200 2450 15252 2456
rect 15384 2450 15436 2456
rect 15396 2378 15424 2450
rect 15384 2372 15436 2378
rect 15384 2314 15436 2320
rect 15198 1592 15254 1601
rect 15198 1527 15254 1536
rect 15212 1426 15240 1527
rect 15396 1494 15424 2314
rect 15568 1896 15620 1902
rect 15568 1838 15620 1844
rect 15660 1896 15712 1902
rect 15660 1838 15712 1844
rect 15384 1488 15436 1494
rect 15384 1430 15436 1436
rect 15108 1420 15160 1426
rect 15108 1362 15160 1368
rect 15200 1420 15252 1426
rect 15200 1362 15252 1368
rect 15580 1358 15608 1838
rect 15672 1562 15700 1838
rect 15752 1760 15804 1766
rect 15752 1702 15804 1708
rect 15660 1556 15712 1562
rect 15660 1498 15712 1504
rect 15764 1426 15792 1702
rect 15856 1426 15884 3334
rect 16684 2990 16712 3538
rect 16776 3466 16804 3878
rect 16764 3460 16816 3466
rect 16764 3402 16816 3408
rect 16672 2984 16724 2990
rect 16672 2926 16724 2932
rect 16212 2848 16264 2854
rect 16212 2790 16264 2796
rect 16764 2848 16816 2854
rect 16764 2790 16816 2796
rect 16224 2582 16252 2790
rect 16364 2748 16740 2757
rect 16420 2746 16444 2748
rect 16500 2746 16524 2748
rect 16580 2746 16604 2748
rect 16660 2746 16684 2748
rect 16420 2694 16430 2746
rect 16674 2694 16684 2746
rect 16420 2692 16444 2694
rect 16500 2692 16524 2694
rect 16580 2692 16604 2694
rect 16660 2692 16684 2694
rect 16364 2683 16740 2692
rect 16580 2644 16632 2650
rect 16580 2586 16632 2592
rect 16212 2576 16264 2582
rect 16212 2518 16264 2524
rect 16302 2544 16358 2553
rect 16302 2479 16304 2488
rect 16356 2479 16358 2488
rect 16304 2450 16356 2456
rect 16212 2440 16264 2446
rect 16212 2382 16264 2388
rect 16224 2310 16252 2382
rect 16212 2304 16264 2310
rect 16212 2246 16264 2252
rect 16120 1964 16172 1970
rect 16120 1906 16172 1912
rect 15936 1828 15988 1834
rect 15936 1770 15988 1776
rect 15948 1601 15976 1770
rect 15934 1592 15990 1601
rect 15934 1527 15990 1536
rect 16132 1426 16160 1906
rect 16224 1562 16252 2246
rect 16592 2106 16620 2586
rect 16580 2100 16632 2106
rect 16580 2042 16632 2048
rect 16364 1660 16740 1669
rect 16420 1658 16444 1660
rect 16500 1658 16524 1660
rect 16580 1658 16604 1660
rect 16660 1658 16684 1660
rect 16420 1606 16430 1658
rect 16674 1606 16684 1658
rect 16420 1604 16444 1606
rect 16500 1604 16524 1606
rect 16580 1604 16604 1606
rect 16660 1604 16684 1606
rect 16364 1595 16740 1604
rect 16212 1556 16264 1562
rect 16212 1498 16264 1504
rect 15752 1420 15804 1426
rect 15752 1362 15804 1368
rect 15844 1420 15896 1426
rect 15844 1362 15896 1368
rect 16120 1420 16172 1426
rect 16120 1362 16172 1368
rect 15568 1352 15620 1358
rect 15028 1278 15240 1306
rect 15568 1294 15620 1300
rect 15016 1216 15068 1222
rect 15016 1158 15068 1164
rect 15108 1216 15160 1222
rect 15108 1158 15160 1164
rect 15028 1018 15056 1158
rect 15016 1012 15068 1018
rect 15016 954 15068 960
rect 14924 944 14976 950
rect 14752 904 14924 932
rect 14464 808 14516 814
rect 14464 750 14516 756
rect 14556 808 14608 814
rect 14556 750 14608 756
rect 14648 808 14700 814
rect 14648 750 14700 756
rect 14372 740 14424 746
rect 14372 682 14424 688
rect 14384 400 14412 682
rect 14280 332 14332 338
rect 14280 274 14332 280
rect 14370 0 14426 400
rect 14568 338 14596 750
rect 14752 400 14780 904
rect 14924 886 14976 892
rect 15120 406 15148 1158
rect 15108 400 15160 406
rect 14556 332 14608 338
rect 14556 274 14608 280
rect 14738 0 14794 400
rect 15108 342 15160 348
rect 15212 134 15240 1278
rect 15580 338 15608 1294
rect 16224 814 16252 1498
rect 16580 1420 16632 1426
rect 16580 1362 16632 1368
rect 16592 1018 16620 1362
rect 16580 1012 16632 1018
rect 16580 954 16632 960
rect 16776 814 16804 2790
rect 16868 2582 16896 4082
rect 16856 2576 16908 2582
rect 16856 2518 16908 2524
rect 17052 2514 17080 4422
rect 17328 3126 17356 5510
rect 17406 5264 17462 5273
rect 17406 5199 17462 5208
rect 17420 5166 17448 5199
rect 17604 5166 17632 8298
rect 17684 8288 17736 8294
rect 17684 8230 17736 8236
rect 17696 7410 17724 8230
rect 17788 7857 17816 8996
rect 17866 8664 17922 8673
rect 17866 8599 17922 8608
rect 17880 8566 17908 8599
rect 17868 8560 17920 8566
rect 17868 8502 17920 8508
rect 17868 8288 17920 8294
rect 17972 8265 18000 10202
rect 17868 8230 17920 8236
rect 17958 8256 18014 8265
rect 17880 8022 17908 8230
rect 17958 8191 18014 8200
rect 17868 8016 17920 8022
rect 17868 7958 17920 7964
rect 17972 7954 18000 8191
rect 17960 7948 18012 7954
rect 17960 7890 18012 7896
rect 17774 7848 17830 7857
rect 17774 7783 17830 7792
rect 17960 7744 18012 7750
rect 17960 7686 18012 7692
rect 17684 7404 17736 7410
rect 17684 7346 17736 7352
rect 17972 6390 18000 7686
rect 17960 6384 18012 6390
rect 17960 6326 18012 6332
rect 17408 5160 17460 5166
rect 17408 5102 17460 5108
rect 17592 5160 17644 5166
rect 17592 5102 17644 5108
rect 17604 4758 17632 5102
rect 17868 5092 17920 5098
rect 17868 5034 17920 5040
rect 17880 4826 17908 5034
rect 17868 4820 17920 4826
rect 17868 4762 17920 4768
rect 17592 4752 17644 4758
rect 17592 4694 17644 4700
rect 17880 4690 17908 4762
rect 17868 4684 17920 4690
rect 17868 4626 17920 4632
rect 17972 3670 18000 6326
rect 18064 5778 18092 11562
rect 18156 9994 18184 11591
rect 18248 10577 18276 13806
rect 18340 12306 18368 16458
rect 18524 15065 18552 16458
rect 18510 15056 18566 15065
rect 18510 14991 18566 15000
rect 18420 14476 18472 14482
rect 18420 14418 18472 14424
rect 18432 13802 18460 14418
rect 18420 13796 18472 13802
rect 18420 13738 18472 13744
rect 18616 13462 18644 19332
rect 18788 19236 18840 19242
rect 18788 19178 18840 19184
rect 18800 18290 18828 19178
rect 18892 18748 18920 20266
rect 18984 19938 19012 21848
rect 19076 21554 19104 21984
rect 19064 21548 19116 21554
rect 19168 21536 19196 22034
rect 19260 21690 19288 22063
rect 19352 22001 19380 22374
rect 19432 22160 19484 22166
rect 19432 22102 19484 22108
rect 19338 21992 19394 22001
rect 19338 21927 19394 21936
rect 19444 21894 19472 22102
rect 19800 21956 19852 21962
rect 19800 21898 19852 21904
rect 19432 21888 19484 21894
rect 19432 21830 19484 21836
rect 19364 21788 19740 21797
rect 19420 21786 19444 21788
rect 19500 21786 19524 21788
rect 19580 21786 19604 21788
rect 19660 21786 19684 21788
rect 19420 21734 19430 21786
rect 19674 21734 19684 21786
rect 19420 21732 19444 21734
rect 19500 21732 19524 21734
rect 19580 21732 19604 21734
rect 19660 21732 19684 21734
rect 19364 21723 19740 21732
rect 19248 21684 19300 21690
rect 19248 21626 19300 21632
rect 19524 21684 19576 21690
rect 19524 21626 19576 21632
rect 19248 21548 19300 21554
rect 19168 21508 19248 21536
rect 19064 21490 19116 21496
rect 19248 21490 19300 21496
rect 19076 21146 19104 21490
rect 19260 21418 19288 21490
rect 19536 21418 19564 21626
rect 19812 21434 19840 21898
rect 19904 21486 19932 23600
rect 20076 23520 20128 23526
rect 20076 23462 20128 23468
rect 20088 23322 20116 23462
rect 20076 23316 20128 23322
rect 20076 23258 20128 23264
rect 20088 22778 20116 23258
rect 20272 23186 20300 23718
rect 20442 23600 20498 23718
rect 20994 23600 21050 24000
rect 21546 23600 21602 24000
rect 22098 23600 22154 24000
rect 22650 23610 22706 24000
rect 22756 23718 22968 23746
rect 22756 23610 22784 23718
rect 22650 23600 22784 23610
rect 20260 23180 20312 23186
rect 20260 23122 20312 23128
rect 20812 23112 20864 23118
rect 20812 23054 20864 23060
rect 20076 22772 20128 22778
rect 20076 22714 20128 22720
rect 20444 22568 20496 22574
rect 20444 22510 20496 22516
rect 20260 22500 20312 22506
rect 20260 22442 20312 22448
rect 20272 22234 20300 22442
rect 20168 22228 20220 22234
rect 20168 22170 20220 22176
rect 20260 22228 20312 22234
rect 20260 22170 20312 22176
rect 20180 22098 20208 22170
rect 19984 22092 20036 22098
rect 19984 22034 20036 22040
rect 20168 22092 20220 22098
rect 20168 22034 20220 22040
rect 20260 22092 20312 22098
rect 20260 22034 20312 22040
rect 19996 21729 20024 22034
rect 19982 21720 20038 21729
rect 19982 21655 20038 21664
rect 20180 21622 20208 22034
rect 20168 21616 20220 21622
rect 20074 21584 20130 21593
rect 20168 21558 20220 21564
rect 20074 21519 20130 21528
rect 20088 21486 20116 21519
rect 19720 21418 19840 21434
rect 19892 21480 19944 21486
rect 19892 21422 19944 21428
rect 20076 21480 20128 21486
rect 20076 21422 20128 21428
rect 20168 21480 20220 21486
rect 20168 21422 20220 21428
rect 19248 21412 19300 21418
rect 19248 21354 19300 21360
rect 19524 21412 19576 21418
rect 19524 21354 19576 21360
rect 19708 21412 19840 21418
rect 19760 21406 19840 21412
rect 19984 21412 20036 21418
rect 19708 21354 19760 21360
rect 19984 21354 20036 21360
rect 19432 21344 19484 21350
rect 19432 21286 19484 21292
rect 19064 21140 19116 21146
rect 19064 21082 19116 21088
rect 19444 20913 19472 21286
rect 19996 21146 20024 21354
rect 20074 21312 20130 21321
rect 20074 21247 20130 21256
rect 19984 21140 20036 21146
rect 19984 21082 20036 21088
rect 20088 21078 20116 21247
rect 20076 21072 20128 21078
rect 20076 21014 20128 21020
rect 19430 20904 19486 20913
rect 20180 20874 20208 21422
rect 19430 20839 19486 20848
rect 20168 20868 20220 20874
rect 20168 20810 20220 20816
rect 19364 20700 19740 20709
rect 19420 20698 19444 20700
rect 19500 20698 19524 20700
rect 19580 20698 19604 20700
rect 19660 20698 19684 20700
rect 19420 20646 19430 20698
rect 19674 20646 19684 20698
rect 19420 20644 19444 20646
rect 19500 20644 19524 20646
rect 19580 20644 19604 20646
rect 19660 20644 19684 20646
rect 19364 20635 19740 20644
rect 19890 20360 19946 20369
rect 19890 20295 19946 20304
rect 19904 20262 19932 20295
rect 19340 20256 19392 20262
rect 19340 20198 19392 20204
rect 19524 20256 19576 20262
rect 19524 20198 19576 20204
rect 19892 20256 19944 20262
rect 19892 20198 19944 20204
rect 18984 19910 19196 19938
rect 19168 19854 19196 19910
rect 18972 19848 19024 19854
rect 18972 19790 19024 19796
rect 19064 19848 19116 19854
rect 19064 19790 19116 19796
rect 19156 19848 19208 19854
rect 19352 19802 19380 20198
rect 19536 20058 19564 20198
rect 19524 20052 19576 20058
rect 19524 19994 19576 20000
rect 20168 19916 20220 19922
rect 20168 19858 20220 19864
rect 19156 19790 19208 19796
rect 18984 19417 19012 19790
rect 18970 19408 19026 19417
rect 18970 19343 19026 19352
rect 19076 19242 19104 19790
rect 19260 19774 19380 19802
rect 19800 19848 19852 19854
rect 19800 19790 19852 19796
rect 19260 19394 19288 19774
rect 19364 19612 19740 19621
rect 19420 19610 19444 19612
rect 19500 19610 19524 19612
rect 19580 19610 19604 19612
rect 19660 19610 19684 19612
rect 19420 19558 19430 19610
rect 19674 19558 19684 19610
rect 19420 19556 19444 19558
rect 19500 19556 19524 19558
rect 19580 19556 19604 19558
rect 19660 19556 19684 19558
rect 19364 19547 19740 19556
rect 19260 19366 19380 19394
rect 18972 19236 19024 19242
rect 18972 19178 19024 19184
rect 19064 19236 19116 19242
rect 19064 19178 19116 19184
rect 18984 18970 19012 19178
rect 19248 19168 19300 19174
rect 19248 19110 19300 19116
rect 18972 18964 19024 18970
rect 18972 18906 19024 18912
rect 19260 18902 19288 19110
rect 19248 18896 19300 18902
rect 19248 18838 19300 18844
rect 18972 18760 19024 18766
rect 18892 18720 18972 18748
rect 19352 18714 19380 19366
rect 19432 19168 19484 19174
rect 19432 19110 19484 19116
rect 19708 19168 19760 19174
rect 19708 19110 19760 19116
rect 19444 18834 19472 19110
rect 19432 18828 19484 18834
rect 19432 18770 19484 18776
rect 18972 18702 19024 18708
rect 18880 18352 18932 18358
rect 18880 18294 18932 18300
rect 18788 18284 18840 18290
rect 18788 18226 18840 18232
rect 18696 18148 18748 18154
rect 18696 18090 18748 18096
rect 18708 17882 18736 18090
rect 18696 17876 18748 17882
rect 18696 17818 18748 17824
rect 18800 17746 18828 18226
rect 18892 18154 18920 18294
rect 18880 18148 18932 18154
rect 18880 18090 18932 18096
rect 18788 17740 18840 17746
rect 18788 17682 18840 17688
rect 18892 17082 18920 18090
rect 18708 17054 18920 17082
rect 18708 15609 18736 17054
rect 18788 16992 18840 16998
rect 18788 16934 18840 16940
rect 18880 16992 18932 16998
rect 18880 16934 18932 16940
rect 18800 16658 18828 16934
rect 18892 16726 18920 16934
rect 18880 16720 18932 16726
rect 18880 16662 18932 16668
rect 18788 16652 18840 16658
rect 18788 16594 18840 16600
rect 18984 15994 19012 18702
rect 19260 18686 19380 18714
rect 19720 18714 19748 19110
rect 19812 18816 19840 19790
rect 20074 19680 20130 19689
rect 20074 19615 20130 19624
rect 19892 18828 19944 18834
rect 19812 18788 19892 18816
rect 19892 18770 19944 18776
rect 19720 18686 19840 18714
rect 19260 18408 19288 18686
rect 19364 18524 19740 18533
rect 19420 18522 19444 18524
rect 19500 18522 19524 18524
rect 19580 18522 19604 18524
rect 19660 18522 19684 18524
rect 19420 18470 19430 18522
rect 19674 18470 19684 18522
rect 19420 18468 19444 18470
rect 19500 18468 19524 18470
rect 19580 18468 19604 18470
rect 19660 18468 19684 18470
rect 19364 18459 19740 18468
rect 19260 18380 19380 18408
rect 19156 18080 19208 18086
rect 19156 18022 19208 18028
rect 19168 17814 19196 18022
rect 19156 17808 19208 17814
rect 19156 17750 19208 17756
rect 19248 17808 19300 17814
rect 19248 17750 19300 17756
rect 19260 17660 19288 17750
rect 19168 17632 19288 17660
rect 19168 17066 19196 17632
rect 19352 17524 19380 18380
rect 19260 17496 19380 17524
rect 19260 17218 19288 17496
rect 19364 17436 19740 17445
rect 19420 17434 19444 17436
rect 19500 17434 19524 17436
rect 19580 17434 19604 17436
rect 19660 17434 19684 17436
rect 19420 17382 19430 17434
rect 19674 17382 19684 17434
rect 19420 17380 19444 17382
rect 19500 17380 19524 17382
rect 19580 17380 19604 17382
rect 19660 17380 19684 17382
rect 19364 17371 19740 17380
rect 19260 17190 19380 17218
rect 19352 17066 19380 17190
rect 19156 17060 19208 17066
rect 19156 17002 19208 17008
rect 19340 17060 19392 17066
rect 19340 17002 19392 17008
rect 19168 16522 19196 17002
rect 19156 16516 19208 16522
rect 19352 16504 19380 17002
rect 19156 16458 19208 16464
rect 19260 16476 19380 16504
rect 19064 16448 19116 16454
rect 19064 16390 19116 16396
rect 19076 16114 19104 16390
rect 19260 16232 19288 16476
rect 19364 16348 19740 16357
rect 19420 16346 19444 16348
rect 19500 16346 19524 16348
rect 19580 16346 19604 16348
rect 19660 16346 19684 16348
rect 19420 16294 19430 16346
rect 19674 16294 19684 16346
rect 19420 16292 19444 16294
rect 19500 16292 19524 16294
rect 19580 16292 19604 16294
rect 19660 16292 19684 16294
rect 19364 16283 19740 16292
rect 19260 16204 19380 16232
rect 19064 16108 19116 16114
rect 19064 16050 19116 16056
rect 18984 15966 19104 15994
rect 18694 15600 18750 15609
rect 18694 15535 18750 15544
rect 18696 15496 18748 15502
rect 18696 15438 18748 15444
rect 18708 15026 18736 15438
rect 18696 15020 18748 15026
rect 18696 14962 18748 14968
rect 18972 15020 19024 15026
rect 18972 14962 19024 14968
rect 18708 14906 18736 14962
rect 18708 14878 18828 14906
rect 18696 14816 18748 14822
rect 18696 14758 18748 14764
rect 18708 14550 18736 14758
rect 18696 14544 18748 14550
rect 18696 14486 18748 14492
rect 18696 14408 18748 14414
rect 18696 14350 18748 14356
rect 18708 14249 18736 14350
rect 18694 14240 18750 14249
rect 18694 14175 18750 14184
rect 18800 13870 18828 14878
rect 18984 14482 19012 14962
rect 18972 14476 19024 14482
rect 18972 14418 19024 14424
rect 18788 13864 18840 13870
rect 18788 13806 18840 13812
rect 18696 13728 18748 13734
rect 18696 13670 18748 13676
rect 18604 13456 18656 13462
rect 18604 13398 18656 13404
rect 18604 13320 18656 13326
rect 18604 13262 18656 13268
rect 18420 13252 18472 13258
rect 18420 13194 18472 13200
rect 18328 12300 18380 12306
rect 18328 12242 18380 12248
rect 18326 11928 18382 11937
rect 18326 11863 18382 11872
rect 18340 11121 18368 11863
rect 18326 11112 18382 11121
rect 18326 11047 18328 11056
rect 18380 11047 18382 11056
rect 18328 11018 18380 11024
rect 18432 10606 18460 13194
rect 18512 12912 18564 12918
rect 18512 12854 18564 12860
rect 18420 10600 18472 10606
rect 18234 10568 18290 10577
rect 18420 10542 18472 10548
rect 18234 10503 18290 10512
rect 18328 10464 18380 10470
rect 18328 10406 18380 10412
rect 18340 10130 18368 10406
rect 18420 10260 18472 10266
rect 18420 10202 18472 10208
rect 18236 10124 18288 10130
rect 18236 10066 18288 10072
rect 18328 10124 18380 10130
rect 18328 10066 18380 10072
rect 18144 9988 18196 9994
rect 18144 9930 18196 9936
rect 18248 9761 18276 10066
rect 18234 9752 18290 9761
rect 18234 9687 18290 9696
rect 18248 9450 18276 9687
rect 18236 9444 18288 9450
rect 18236 9386 18288 9392
rect 18144 9376 18196 9382
rect 18196 9324 18276 9330
rect 18144 9318 18276 9324
rect 18156 9302 18276 9318
rect 18142 9208 18198 9217
rect 18142 9143 18144 9152
rect 18196 9143 18198 9152
rect 18144 9114 18196 9120
rect 18142 9072 18198 9081
rect 18248 9042 18276 9302
rect 18142 9007 18198 9016
rect 18236 9036 18288 9042
rect 18156 8566 18184 9007
rect 18236 8978 18288 8984
rect 18234 8936 18290 8945
rect 18234 8871 18290 8880
rect 18144 8560 18196 8566
rect 18144 8502 18196 8508
rect 18142 7576 18198 7585
rect 18142 7511 18198 7520
rect 18156 6746 18184 7511
rect 18248 6866 18276 8871
rect 18340 6866 18368 10066
rect 18432 9897 18460 10202
rect 18418 9888 18474 9897
rect 18418 9823 18474 9832
rect 18524 9160 18552 12854
rect 18616 11354 18644 13262
rect 18708 12442 18736 13670
rect 18880 13184 18932 13190
rect 18880 13126 18932 13132
rect 18788 12844 18840 12850
rect 18788 12786 18840 12792
rect 18800 12646 18828 12786
rect 18892 12782 18920 13126
rect 18880 12776 18932 12782
rect 18880 12718 18932 12724
rect 18788 12640 18840 12646
rect 18788 12582 18840 12588
rect 18696 12436 18748 12442
rect 18696 12378 18748 12384
rect 18696 12300 18748 12306
rect 18696 12242 18748 12248
rect 18708 11778 18736 12242
rect 18788 12096 18840 12102
rect 18788 12038 18840 12044
rect 18880 12096 18932 12102
rect 18880 12038 18932 12044
rect 18800 11898 18828 12038
rect 18788 11892 18840 11898
rect 18788 11834 18840 11840
rect 18708 11750 18828 11778
rect 18892 11762 18920 12038
rect 18696 11620 18748 11626
rect 18696 11562 18748 11568
rect 18708 11529 18736 11562
rect 18694 11520 18750 11529
rect 18694 11455 18750 11464
rect 18604 11348 18656 11354
rect 18604 11290 18656 11296
rect 18616 11200 18644 11290
rect 18696 11212 18748 11218
rect 18616 11172 18696 11200
rect 18696 11154 18748 11160
rect 18696 11076 18748 11082
rect 18696 11018 18748 11024
rect 18708 10674 18736 11018
rect 18696 10668 18748 10674
rect 18696 10610 18748 10616
rect 18604 10600 18656 10606
rect 18604 10542 18656 10548
rect 18616 10033 18644 10542
rect 18602 10024 18658 10033
rect 18602 9959 18658 9968
rect 18800 9353 18828 11750
rect 18880 11756 18932 11762
rect 18880 11698 18932 11704
rect 19076 11694 19104 15966
rect 19352 15473 19380 16204
rect 19708 16040 19760 16046
rect 19708 15982 19760 15988
rect 19432 15904 19484 15910
rect 19432 15846 19484 15852
rect 19444 15570 19472 15846
rect 19720 15570 19748 15982
rect 19432 15564 19484 15570
rect 19432 15506 19484 15512
rect 19708 15564 19760 15570
rect 19708 15506 19760 15512
rect 19338 15464 19394 15473
rect 19156 15428 19208 15434
rect 19338 15399 19394 15408
rect 19156 15370 19208 15376
rect 19168 15026 19196 15370
rect 19248 15360 19300 15366
rect 19248 15302 19300 15308
rect 19260 15042 19288 15302
rect 19364 15260 19740 15269
rect 19420 15258 19444 15260
rect 19500 15258 19524 15260
rect 19580 15258 19604 15260
rect 19660 15258 19684 15260
rect 19420 15206 19430 15258
rect 19674 15206 19684 15258
rect 19420 15204 19444 15206
rect 19500 15204 19524 15206
rect 19580 15204 19604 15206
rect 19660 15204 19684 15206
rect 19364 15195 19740 15204
rect 19812 15094 19840 18686
rect 19904 18601 19932 18770
rect 20088 18698 20116 19615
rect 20180 18766 20208 19858
rect 20272 19786 20300 22034
rect 20352 22024 20404 22030
rect 20352 21966 20404 21972
rect 20364 20806 20392 21966
rect 20456 21146 20484 22510
rect 20628 22500 20680 22506
rect 20628 22442 20680 22448
rect 20720 22500 20772 22506
rect 20720 22442 20772 22448
rect 20640 22234 20668 22442
rect 20628 22228 20680 22234
rect 20628 22170 20680 22176
rect 20536 22024 20588 22030
rect 20536 21966 20588 21972
rect 20548 21486 20576 21966
rect 20536 21480 20588 21486
rect 20536 21422 20588 21428
rect 20444 21140 20496 21146
rect 20444 21082 20496 21088
rect 20352 20800 20404 20806
rect 20352 20742 20404 20748
rect 20364 20058 20392 20742
rect 20548 20330 20576 21422
rect 20640 20788 20668 22170
rect 20732 22166 20760 22442
rect 20720 22160 20772 22166
rect 20720 22102 20772 22108
rect 20824 21978 20852 23054
rect 20904 22704 20956 22710
rect 20904 22646 20956 22652
rect 20732 21950 20852 21978
rect 20732 21010 20760 21950
rect 20812 21888 20864 21894
rect 20812 21830 20864 21836
rect 20824 21690 20852 21830
rect 20812 21684 20864 21690
rect 20812 21626 20864 21632
rect 20812 21412 20864 21418
rect 20812 21354 20864 21360
rect 20824 21078 20852 21354
rect 20916 21078 20944 22646
rect 21008 21078 21036 23600
rect 21560 23254 21588 23600
rect 21548 23248 21600 23254
rect 21548 23190 21600 23196
rect 21364 22976 21416 22982
rect 21640 22976 21692 22982
rect 21364 22918 21416 22924
rect 21638 22944 21640 22953
rect 21692 22944 21694 22953
rect 21088 22568 21140 22574
rect 21140 22528 21220 22556
rect 21088 22510 21140 22516
rect 21088 22432 21140 22438
rect 21088 22374 21140 22380
rect 21100 22273 21128 22374
rect 21086 22264 21142 22273
rect 21086 22199 21142 22208
rect 21192 22114 21220 22528
rect 21100 22086 21220 22114
rect 21100 21622 21128 22086
rect 21272 22024 21324 22030
rect 21272 21966 21324 21972
rect 21284 21894 21312 21966
rect 21180 21888 21232 21894
rect 21180 21830 21232 21836
rect 21272 21888 21324 21894
rect 21272 21830 21324 21836
rect 21088 21616 21140 21622
rect 21088 21558 21140 21564
rect 20812 21072 20864 21078
rect 20812 21014 20864 21020
rect 20904 21072 20956 21078
rect 20904 21014 20956 21020
rect 20996 21072 21048 21078
rect 20996 21014 21048 21020
rect 20720 21004 20772 21010
rect 20720 20946 20772 20952
rect 20732 20913 20760 20946
rect 20718 20904 20774 20913
rect 20718 20839 20774 20848
rect 20824 20788 20852 21014
rect 21100 21010 21128 21558
rect 21088 21004 21140 21010
rect 21088 20946 21140 20952
rect 21088 20868 21140 20874
rect 21088 20810 21140 20816
rect 20640 20760 20852 20788
rect 20720 20528 20772 20534
rect 20812 20528 20864 20534
rect 20720 20470 20772 20476
rect 20810 20496 20812 20505
rect 20864 20496 20866 20505
rect 20732 20380 20760 20470
rect 20810 20431 20866 20440
rect 20904 20392 20956 20398
rect 20626 20360 20682 20369
rect 20444 20324 20496 20330
rect 20444 20266 20496 20272
rect 20536 20324 20588 20330
rect 20732 20352 20852 20380
rect 20626 20295 20682 20304
rect 20536 20266 20588 20272
rect 20456 20058 20484 20266
rect 20352 20052 20404 20058
rect 20352 19994 20404 20000
rect 20444 20052 20496 20058
rect 20640 20040 20668 20295
rect 20720 20256 20772 20262
rect 20720 20198 20772 20204
rect 20444 19994 20496 20000
rect 20548 20012 20668 20040
rect 20260 19780 20312 19786
rect 20260 19722 20312 19728
rect 20272 19446 20300 19722
rect 20260 19440 20312 19446
rect 20260 19382 20312 19388
rect 20260 19304 20312 19310
rect 20260 19246 20312 19252
rect 20168 18760 20220 18766
rect 20168 18702 20220 18708
rect 20076 18692 20128 18698
rect 20076 18634 20128 18640
rect 19984 18624 20036 18630
rect 19890 18592 19946 18601
rect 19984 18566 20036 18572
rect 19890 18527 19946 18536
rect 19996 18222 20024 18566
rect 20088 18222 20116 18634
rect 19984 18216 20036 18222
rect 19984 18158 20036 18164
rect 20076 18216 20128 18222
rect 20076 18158 20128 18164
rect 20088 17678 20116 18158
rect 20076 17672 20128 17678
rect 20076 17614 20128 17620
rect 19984 17536 20036 17542
rect 19984 17478 20036 17484
rect 20076 17536 20128 17542
rect 20076 17478 20128 17484
rect 19892 17332 19944 17338
rect 19892 17274 19944 17280
rect 19904 16726 19932 17274
rect 19996 17066 20024 17478
rect 19984 17060 20036 17066
rect 19984 17002 20036 17008
rect 20088 16726 20116 17478
rect 19892 16720 19944 16726
rect 19892 16662 19944 16668
rect 20076 16720 20128 16726
rect 20076 16662 20128 16668
rect 19890 16552 19946 16561
rect 19890 16487 19946 16496
rect 19340 15088 19392 15094
rect 19260 15036 19340 15042
rect 19260 15030 19392 15036
rect 19800 15088 19852 15094
rect 19800 15030 19852 15036
rect 19156 15020 19208 15026
rect 19260 15014 19380 15030
rect 19156 14962 19208 14968
rect 19248 14952 19300 14958
rect 19248 14894 19300 14900
rect 19260 14618 19288 14894
rect 19352 14890 19380 15014
rect 19524 14952 19576 14958
rect 19524 14894 19576 14900
rect 19340 14884 19392 14890
rect 19340 14826 19392 14832
rect 19536 14822 19564 14894
rect 19812 14890 19840 15030
rect 19800 14884 19852 14890
rect 19800 14826 19852 14832
rect 19524 14816 19576 14822
rect 19524 14758 19576 14764
rect 19248 14612 19300 14618
rect 19248 14554 19300 14560
rect 19338 14512 19394 14521
rect 19338 14447 19394 14456
rect 19352 14414 19380 14447
rect 19340 14408 19392 14414
rect 19340 14350 19392 14356
rect 19248 14340 19300 14346
rect 19248 14282 19300 14288
rect 19260 14056 19288 14282
rect 19536 14278 19564 14758
rect 19904 14414 19932 16487
rect 20076 16448 20128 16454
rect 20076 16390 20128 16396
rect 20088 16046 20116 16390
rect 20076 16040 20128 16046
rect 20076 15982 20128 15988
rect 20180 15722 20208 18702
rect 20272 16182 20300 19246
rect 20364 19122 20392 19994
rect 20456 19514 20484 19994
rect 20548 19854 20576 20012
rect 20626 19952 20682 19961
rect 20626 19887 20628 19896
rect 20680 19887 20682 19896
rect 20628 19858 20680 19864
rect 20536 19848 20588 19854
rect 20536 19790 20588 19796
rect 20536 19712 20588 19718
rect 20640 19689 20668 19858
rect 20536 19654 20588 19660
rect 20626 19680 20682 19689
rect 20444 19508 20496 19514
rect 20444 19450 20496 19456
rect 20548 19378 20576 19654
rect 20626 19615 20682 19624
rect 20732 19514 20760 20198
rect 20824 19922 20852 20352
rect 20904 20334 20956 20340
rect 20996 20392 21048 20398
rect 20996 20334 21048 20340
rect 20812 19916 20864 19922
rect 20812 19858 20864 19864
rect 20810 19816 20866 19825
rect 20810 19751 20812 19760
rect 20864 19751 20866 19760
rect 20812 19722 20864 19728
rect 20720 19508 20772 19514
rect 20720 19450 20772 19456
rect 20536 19372 20588 19378
rect 20536 19314 20588 19320
rect 20732 19310 20760 19450
rect 20628 19304 20680 19310
rect 20626 19272 20628 19281
rect 20720 19304 20772 19310
rect 20680 19272 20682 19281
rect 20720 19246 20772 19252
rect 20626 19207 20682 19216
rect 20364 19094 20668 19122
rect 20444 18964 20496 18970
rect 20444 18906 20496 18912
rect 20456 18766 20484 18906
rect 20536 18828 20588 18834
rect 20536 18770 20588 18776
rect 20444 18760 20496 18766
rect 20444 18702 20496 18708
rect 20456 17490 20484 18702
rect 20548 18057 20576 18770
rect 20534 18048 20590 18057
rect 20534 17983 20590 17992
rect 20456 17462 20576 17490
rect 20444 16448 20496 16454
rect 20444 16390 20496 16396
rect 20260 16176 20312 16182
rect 20260 16118 20312 16124
rect 20456 16046 20484 16390
rect 20444 16040 20496 16046
rect 20444 15982 20496 15988
rect 20352 15904 20404 15910
rect 20352 15846 20404 15852
rect 20088 15694 20208 15722
rect 19984 15088 20036 15094
rect 19984 15030 20036 15036
rect 19996 14822 20024 15030
rect 19984 14816 20036 14822
rect 19984 14758 20036 14764
rect 19984 14476 20036 14482
rect 19984 14418 20036 14424
rect 19892 14408 19944 14414
rect 19892 14350 19944 14356
rect 19524 14272 19576 14278
rect 19524 14214 19576 14220
rect 19364 14172 19740 14181
rect 19420 14170 19444 14172
rect 19500 14170 19524 14172
rect 19580 14170 19604 14172
rect 19660 14170 19684 14172
rect 19420 14118 19430 14170
rect 19674 14118 19684 14170
rect 19420 14116 19444 14118
rect 19500 14116 19524 14118
rect 19580 14116 19604 14118
rect 19660 14116 19684 14118
rect 19364 14107 19740 14116
rect 19340 14068 19392 14074
rect 19260 14028 19340 14056
rect 19340 14010 19392 14016
rect 19352 13870 19380 14010
rect 19616 14000 19668 14006
rect 19616 13942 19668 13948
rect 19340 13864 19392 13870
rect 19340 13806 19392 13812
rect 19628 13394 19656 13942
rect 19996 13938 20024 14418
rect 19708 13932 19760 13938
rect 19708 13874 19760 13880
rect 19984 13932 20036 13938
rect 19984 13874 20036 13880
rect 19720 13530 19748 13874
rect 19800 13728 19852 13734
rect 19800 13670 19852 13676
rect 19984 13728 20036 13734
rect 19984 13670 20036 13676
rect 19708 13524 19760 13530
rect 19708 13466 19760 13472
rect 19616 13388 19668 13394
rect 19616 13330 19668 13336
rect 19364 13084 19740 13093
rect 19420 13082 19444 13084
rect 19500 13082 19524 13084
rect 19580 13082 19604 13084
rect 19660 13082 19684 13084
rect 19420 13030 19430 13082
rect 19674 13030 19684 13082
rect 19420 13028 19444 13030
rect 19500 13028 19524 13030
rect 19580 13028 19604 13030
rect 19660 13028 19684 13030
rect 19364 13019 19740 13028
rect 19338 12880 19394 12889
rect 19522 12880 19578 12889
rect 19338 12815 19394 12824
rect 19432 12844 19484 12850
rect 19352 12764 19380 12815
rect 19522 12815 19578 12824
rect 19432 12786 19484 12792
rect 19306 12736 19380 12764
rect 19306 12646 19334 12736
rect 19294 12640 19346 12646
rect 19294 12582 19346 12588
rect 19444 12306 19472 12786
rect 19536 12782 19564 12815
rect 19524 12776 19576 12782
rect 19524 12718 19576 12724
rect 19432 12300 19484 12306
rect 19432 12242 19484 12248
rect 19524 12300 19576 12306
rect 19524 12242 19576 12248
rect 19444 12084 19472 12242
rect 19536 12209 19564 12242
rect 19522 12200 19578 12209
rect 19522 12135 19524 12144
rect 19576 12135 19578 12144
rect 19524 12106 19576 12112
rect 19260 12056 19472 12084
rect 19260 11778 19288 12056
rect 19364 11996 19740 12005
rect 19420 11994 19444 11996
rect 19500 11994 19524 11996
rect 19580 11994 19604 11996
rect 19660 11994 19684 11996
rect 19420 11942 19430 11994
rect 19674 11942 19684 11994
rect 19420 11940 19444 11942
rect 19500 11940 19524 11942
rect 19580 11940 19604 11942
rect 19660 11940 19684 11942
rect 19364 11931 19740 11940
rect 19522 11792 19578 11801
rect 19260 11762 19380 11778
rect 19260 11756 19392 11762
rect 19260 11750 19340 11756
rect 19340 11698 19392 11704
rect 19432 11756 19484 11762
rect 19522 11727 19578 11736
rect 19432 11698 19484 11704
rect 19064 11688 19116 11694
rect 19064 11630 19116 11636
rect 19248 11688 19300 11694
rect 19248 11630 19300 11636
rect 19064 11552 19116 11558
rect 19062 11520 19064 11529
rect 19116 11520 19118 11529
rect 19062 11455 19118 11464
rect 18878 11248 18934 11257
rect 18878 11183 18934 11192
rect 19064 11212 19116 11218
rect 18786 9344 18842 9353
rect 18786 9279 18842 9288
rect 18892 9194 18920 11183
rect 19064 11154 19116 11160
rect 19076 10538 19104 11154
rect 19260 10792 19288 11630
rect 19340 11144 19392 11150
rect 19338 11112 19340 11121
rect 19392 11112 19394 11121
rect 19338 11047 19394 11056
rect 19340 11008 19392 11014
rect 19444 10996 19472 11698
rect 19536 11014 19564 11727
rect 19392 10968 19472 10996
rect 19524 11008 19576 11014
rect 19340 10950 19392 10956
rect 19524 10950 19576 10956
rect 19364 10908 19740 10917
rect 19420 10906 19444 10908
rect 19500 10906 19524 10908
rect 19580 10906 19604 10908
rect 19660 10906 19684 10908
rect 19420 10854 19430 10906
rect 19674 10854 19684 10906
rect 19420 10852 19444 10854
rect 19500 10852 19524 10854
rect 19580 10852 19604 10854
rect 19660 10852 19684 10854
rect 19364 10843 19740 10852
rect 19260 10764 19380 10792
rect 19246 10704 19302 10713
rect 19246 10639 19302 10648
rect 19064 10532 19116 10538
rect 19064 10474 19116 10480
rect 19260 10198 19288 10639
rect 19248 10192 19300 10198
rect 19248 10134 19300 10140
rect 19064 9920 19116 9926
rect 19352 9908 19380 10764
rect 19614 10568 19670 10577
rect 19614 10503 19670 10512
rect 19432 10464 19484 10470
rect 19432 10406 19484 10412
rect 19444 9926 19472 10406
rect 19628 10130 19656 10503
rect 19616 10124 19668 10130
rect 19616 10066 19668 10072
rect 19064 9862 19116 9868
rect 19260 9880 19380 9908
rect 19432 9920 19484 9926
rect 19076 9654 19104 9862
rect 19064 9648 19116 9654
rect 19260 9636 19288 9880
rect 19432 9862 19484 9868
rect 19364 9820 19740 9829
rect 19420 9818 19444 9820
rect 19500 9818 19524 9820
rect 19580 9818 19604 9820
rect 19660 9818 19684 9820
rect 19420 9766 19430 9818
rect 19674 9766 19684 9818
rect 19420 9764 19444 9766
rect 19500 9764 19524 9766
rect 19580 9764 19604 9766
rect 19660 9764 19684 9766
rect 19364 9755 19740 9764
rect 19260 9608 19380 9636
rect 19064 9590 19116 9596
rect 19248 9376 19300 9382
rect 19248 9318 19300 9324
rect 18800 9166 18920 9194
rect 19260 9178 19288 9318
rect 19352 9217 19380 9608
rect 19432 9512 19484 9518
rect 19430 9480 19432 9489
rect 19484 9480 19486 9489
rect 19430 9415 19486 9424
rect 19338 9208 19394 9217
rect 19248 9172 19300 9178
rect 18524 9132 18644 9160
rect 18512 9036 18564 9042
rect 18512 8978 18564 8984
rect 18524 8906 18552 8978
rect 18512 8900 18564 8906
rect 18512 8842 18564 8848
rect 18420 8832 18472 8838
rect 18420 8774 18472 8780
rect 18432 8673 18460 8774
rect 18418 8664 18474 8673
rect 18418 8599 18474 8608
rect 18420 8560 18472 8566
rect 18420 8502 18472 8508
rect 18432 8430 18460 8502
rect 18420 8424 18472 8430
rect 18420 8366 18472 8372
rect 18432 7993 18460 8366
rect 18418 7984 18474 7993
rect 18418 7919 18474 7928
rect 18420 7880 18472 7886
rect 18524 7868 18552 8842
rect 18472 7840 18552 7868
rect 18420 7822 18472 7828
rect 18236 6860 18288 6866
rect 18236 6802 18288 6808
rect 18328 6860 18380 6866
rect 18328 6802 18380 6808
rect 18512 6792 18564 6798
rect 18156 6718 18276 6746
rect 18512 6734 18564 6740
rect 18144 6656 18196 6662
rect 18144 6598 18196 6604
rect 18156 6390 18184 6598
rect 18144 6384 18196 6390
rect 18144 6326 18196 6332
rect 18052 5772 18104 5778
rect 18052 5714 18104 5720
rect 18248 5030 18276 6718
rect 18524 6662 18552 6734
rect 18420 6656 18472 6662
rect 18420 6598 18472 6604
rect 18512 6656 18564 6662
rect 18512 6598 18564 6604
rect 18328 6316 18380 6322
rect 18328 6258 18380 6264
rect 18236 5024 18288 5030
rect 18236 4966 18288 4972
rect 18340 4672 18368 6258
rect 18432 5778 18460 6598
rect 18512 6112 18564 6118
rect 18512 6054 18564 6060
rect 18420 5772 18472 5778
rect 18420 5714 18472 5720
rect 18524 5574 18552 6054
rect 18616 5778 18644 9132
rect 18694 8664 18750 8673
rect 18694 8599 18750 8608
rect 18708 7954 18736 8599
rect 18696 7948 18748 7954
rect 18696 7890 18748 7896
rect 18694 7848 18750 7857
rect 18800 7834 18828 9166
rect 19338 9143 19394 9152
rect 19248 9114 19300 9120
rect 19062 9072 19118 9081
rect 19062 9007 19064 9016
rect 19116 9007 19118 9016
rect 19708 9036 19760 9042
rect 19064 8978 19116 8984
rect 19812 9024 19840 13670
rect 19892 13456 19944 13462
rect 19892 13398 19944 13404
rect 19904 12986 19932 13398
rect 19892 12980 19944 12986
rect 19892 12922 19944 12928
rect 19892 12776 19944 12782
rect 19892 12718 19944 12724
rect 19904 12442 19932 12718
rect 19892 12436 19944 12442
rect 19892 12378 19944 12384
rect 19904 11898 19932 12378
rect 19996 12306 20024 13670
rect 20088 13190 20116 15694
rect 20168 15632 20220 15638
rect 20168 15574 20220 15580
rect 20076 13184 20128 13190
rect 20076 13126 20128 13132
rect 20180 12889 20208 15574
rect 20364 15366 20392 15846
rect 20456 15502 20484 15982
rect 20444 15496 20496 15502
rect 20444 15438 20496 15444
rect 20548 15434 20576 17462
rect 20536 15428 20588 15434
rect 20536 15370 20588 15376
rect 20260 15360 20312 15366
rect 20260 15302 20312 15308
rect 20352 15360 20404 15366
rect 20352 15302 20404 15308
rect 20272 13938 20300 15302
rect 20352 14816 20404 14822
rect 20352 14758 20404 14764
rect 20444 14816 20496 14822
rect 20444 14758 20496 14764
rect 20364 14482 20392 14758
rect 20456 14482 20484 14758
rect 20352 14476 20404 14482
rect 20352 14418 20404 14424
rect 20444 14476 20496 14482
rect 20496 14436 20576 14464
rect 20444 14418 20496 14424
rect 20364 14006 20392 14418
rect 20444 14272 20496 14278
rect 20444 14214 20496 14220
rect 20352 14000 20404 14006
rect 20352 13942 20404 13948
rect 20260 13932 20312 13938
rect 20260 13874 20312 13880
rect 20260 13184 20312 13190
rect 20260 13126 20312 13132
rect 20166 12880 20222 12889
rect 20166 12815 20222 12824
rect 20076 12776 20128 12782
rect 20076 12718 20128 12724
rect 19984 12300 20036 12306
rect 19984 12242 20036 12248
rect 19996 11898 20024 12242
rect 20088 11898 20116 12718
rect 20272 12322 20300 13126
rect 20456 12968 20484 14214
rect 20548 13870 20576 14436
rect 20536 13864 20588 13870
rect 20536 13806 20588 13812
rect 20536 13728 20588 13734
rect 20536 13670 20588 13676
rect 20548 13394 20576 13670
rect 20536 13388 20588 13394
rect 20536 13330 20588 13336
rect 20640 13274 20668 19094
rect 20916 18970 20944 20334
rect 21008 19310 21036 20334
rect 21100 19922 21128 20810
rect 21192 20466 21220 21830
rect 21284 20942 21312 21830
rect 21376 21486 21404 22918
rect 21638 22879 21694 22888
rect 21652 22506 21680 22879
rect 21640 22500 21692 22506
rect 21640 22442 21692 22448
rect 21548 22092 21600 22098
rect 21548 22034 21600 22040
rect 21454 21720 21510 21729
rect 21454 21655 21510 21664
rect 21468 21622 21496 21655
rect 21456 21616 21508 21622
rect 21456 21558 21508 21564
rect 21364 21480 21416 21486
rect 21560 21457 21588 22034
rect 21364 21422 21416 21428
rect 21546 21448 21602 21457
rect 21546 21383 21602 21392
rect 21822 21448 21878 21457
rect 21822 21383 21878 21392
rect 22008 21412 22060 21418
rect 21456 21344 21508 21350
rect 21454 21312 21456 21321
rect 21508 21312 21510 21321
rect 21454 21247 21510 21256
rect 21272 20936 21324 20942
rect 21272 20878 21324 20884
rect 21640 20936 21692 20942
rect 21640 20878 21692 20884
rect 21180 20460 21232 20466
rect 21180 20402 21232 20408
rect 21272 20392 21324 20398
rect 21272 20334 21324 20340
rect 21364 20392 21416 20398
rect 21364 20334 21416 20340
rect 21548 20392 21600 20398
rect 21548 20334 21600 20340
rect 21284 20058 21312 20334
rect 21376 20058 21404 20334
rect 21456 20324 21508 20330
rect 21456 20266 21508 20272
rect 21272 20052 21324 20058
rect 21272 19994 21324 20000
rect 21364 20052 21416 20058
rect 21364 19994 21416 20000
rect 21088 19916 21140 19922
rect 21088 19858 21140 19864
rect 21180 19848 21232 19854
rect 21100 19796 21180 19802
rect 21100 19790 21232 19796
rect 21100 19774 21220 19790
rect 21100 19310 21128 19774
rect 21284 19530 21312 19994
rect 21364 19916 21416 19922
rect 21364 19858 21416 19864
rect 21376 19825 21404 19858
rect 21362 19816 21418 19825
rect 21362 19751 21418 19760
rect 21284 19502 21404 19530
rect 21270 19408 21326 19417
rect 21180 19372 21232 19378
rect 21270 19343 21326 19352
rect 21180 19314 21232 19320
rect 20996 19304 21048 19310
rect 20996 19246 21048 19252
rect 21088 19304 21140 19310
rect 21088 19246 21140 19252
rect 20904 18964 20956 18970
rect 20904 18906 20956 18912
rect 21008 18766 21036 19246
rect 21088 18896 21140 18902
rect 21088 18838 21140 18844
rect 20996 18760 21048 18766
rect 20996 18702 21048 18708
rect 21100 18426 21128 18838
rect 21192 18834 21220 19314
rect 21180 18828 21232 18834
rect 21180 18770 21232 18776
rect 21088 18420 21140 18426
rect 21088 18362 21140 18368
rect 20904 18080 20956 18086
rect 20904 18022 20956 18028
rect 20720 17740 20772 17746
rect 20720 17682 20772 17688
rect 20732 17649 20760 17682
rect 20812 17672 20864 17678
rect 20718 17640 20774 17649
rect 20812 17614 20864 17620
rect 20718 17575 20774 17584
rect 20824 17202 20852 17614
rect 20812 17196 20864 17202
rect 20812 17138 20864 17144
rect 20824 17105 20852 17138
rect 20810 17096 20866 17105
rect 20810 17031 20866 17040
rect 20718 16688 20774 16697
rect 20718 16623 20720 16632
rect 20772 16623 20774 16632
rect 20720 16594 20772 16600
rect 20812 15564 20864 15570
rect 20812 15506 20864 15512
rect 20720 15360 20772 15366
rect 20720 15302 20772 15308
rect 20732 15162 20760 15302
rect 20720 15156 20772 15162
rect 20720 15098 20772 15104
rect 20824 14958 20852 15506
rect 20812 14952 20864 14958
rect 20812 14894 20864 14900
rect 20812 14000 20864 14006
rect 20812 13942 20864 13948
rect 20364 12940 20484 12968
rect 20548 13246 20668 13274
rect 20824 13258 20852 13942
rect 20812 13252 20864 13258
rect 20364 12442 20392 12940
rect 20444 12844 20496 12850
rect 20444 12786 20496 12792
rect 20352 12436 20404 12442
rect 20352 12378 20404 12384
rect 20272 12294 20392 12322
rect 20168 12232 20220 12238
rect 20168 12174 20220 12180
rect 20260 12232 20312 12238
rect 20260 12174 20312 12180
rect 19892 11892 19944 11898
rect 19892 11834 19944 11840
rect 19984 11892 20036 11898
rect 19984 11834 20036 11840
rect 20076 11892 20128 11898
rect 20076 11834 20128 11840
rect 19892 11756 19944 11762
rect 19892 11698 19944 11704
rect 19904 10266 19932 11698
rect 20180 11694 20208 12174
rect 20272 11694 20300 12174
rect 20168 11688 20220 11694
rect 20168 11630 20220 11636
rect 20260 11688 20312 11694
rect 20260 11630 20312 11636
rect 19984 11620 20036 11626
rect 19984 11562 20036 11568
rect 19892 10260 19944 10266
rect 19892 10202 19944 10208
rect 19996 10130 20024 11562
rect 20260 11552 20312 11558
rect 20260 11494 20312 11500
rect 20168 11348 20220 11354
rect 20168 11290 20220 11296
rect 20180 11218 20208 11290
rect 20272 11257 20300 11494
rect 20258 11248 20314 11257
rect 20076 11212 20128 11218
rect 20076 11154 20128 11160
rect 20168 11212 20220 11218
rect 20258 11183 20314 11192
rect 20168 11154 20220 11160
rect 20088 10606 20116 11154
rect 20180 10810 20208 11154
rect 20272 11082 20300 11183
rect 20260 11076 20312 11082
rect 20260 11018 20312 11024
rect 20168 10804 20220 10810
rect 20168 10746 20220 10752
rect 20076 10600 20128 10606
rect 20076 10542 20128 10548
rect 20180 10538 20208 10746
rect 20168 10532 20220 10538
rect 20168 10474 20220 10480
rect 20076 10464 20128 10470
rect 20076 10406 20128 10412
rect 20088 10198 20116 10406
rect 20076 10192 20128 10198
rect 20076 10134 20128 10140
rect 19984 10124 20036 10130
rect 19984 10066 20036 10072
rect 20260 10056 20312 10062
rect 20260 9998 20312 10004
rect 20168 9988 20220 9994
rect 20168 9930 20220 9936
rect 19984 9920 20036 9926
rect 19984 9862 20036 9868
rect 19996 9738 20024 9862
rect 19904 9722 20024 9738
rect 19892 9716 20024 9722
rect 19944 9710 20024 9716
rect 20076 9716 20128 9722
rect 19892 9658 19944 9664
rect 19996 9664 20076 9674
rect 19996 9658 20128 9664
rect 19996 9646 20116 9658
rect 19892 9580 19944 9586
rect 19892 9522 19944 9528
rect 19904 9489 19932 9522
rect 19890 9480 19946 9489
rect 19890 9415 19946 9424
rect 19892 9036 19944 9042
rect 19812 8996 19892 9024
rect 19708 8978 19760 8984
rect 19892 8978 19944 8984
rect 19720 8945 19748 8978
rect 19246 8936 19302 8945
rect 19246 8871 19302 8880
rect 19706 8936 19762 8945
rect 19996 8922 20024 9646
rect 20076 9512 20128 9518
rect 20074 9480 20076 9489
rect 20128 9480 20130 9489
rect 20074 9415 20130 9424
rect 20076 9376 20128 9382
rect 20076 9318 20128 9324
rect 19904 8906 20024 8922
rect 19706 8871 19762 8880
rect 19892 8900 20024 8906
rect 18880 8832 18932 8838
rect 18880 8774 18932 8780
rect 18970 8800 19026 8809
rect 18892 7954 18920 8774
rect 18970 8735 19026 8744
rect 18984 8634 19012 8735
rect 18972 8628 19024 8634
rect 18972 8570 19024 8576
rect 19154 8256 19210 8265
rect 19154 8191 19210 8200
rect 19168 8022 19196 8191
rect 19156 8016 19208 8022
rect 19156 7958 19208 7964
rect 18880 7948 18932 7954
rect 18880 7890 18932 7896
rect 18800 7806 19196 7834
rect 18694 7783 18750 7792
rect 18708 7478 18736 7783
rect 18788 7744 18840 7750
rect 18788 7686 18840 7692
rect 18880 7744 18932 7750
rect 18880 7686 18932 7692
rect 18970 7712 19026 7721
rect 18696 7472 18748 7478
rect 18696 7414 18748 7420
rect 18800 6254 18828 7686
rect 18892 6322 18920 7686
rect 18970 7647 19026 7656
rect 18984 6798 19012 7647
rect 18972 6792 19024 6798
rect 18972 6734 19024 6740
rect 18880 6316 18932 6322
rect 18880 6258 18932 6264
rect 18788 6248 18840 6254
rect 18788 6190 18840 6196
rect 18696 6112 18748 6118
rect 18696 6054 18748 6060
rect 18708 5846 18736 6054
rect 18696 5840 18748 5846
rect 18696 5782 18748 5788
rect 18604 5772 18656 5778
rect 18604 5714 18656 5720
rect 18604 5636 18656 5642
rect 18604 5578 18656 5584
rect 18512 5568 18564 5574
rect 18512 5510 18564 5516
rect 18616 4706 18644 5578
rect 18696 5160 18748 5166
rect 18696 5102 18748 5108
rect 18524 4690 18644 4706
rect 18420 4684 18472 4690
rect 18340 4644 18420 4672
rect 18420 4626 18472 4632
rect 18512 4684 18644 4690
rect 18564 4678 18644 4684
rect 18512 4626 18564 4632
rect 18052 4616 18104 4622
rect 18050 4584 18052 4593
rect 18104 4584 18106 4593
rect 18050 4519 18106 4528
rect 18064 4214 18092 4519
rect 18052 4208 18104 4214
rect 18052 4150 18104 4156
rect 17960 3664 18012 3670
rect 17960 3606 18012 3612
rect 18524 3534 18552 4626
rect 18604 4616 18656 4622
rect 18604 4558 18656 4564
rect 18512 3528 18564 3534
rect 18512 3470 18564 3476
rect 17684 3460 17736 3466
rect 17684 3402 17736 3408
rect 18052 3460 18104 3466
rect 18052 3402 18104 3408
rect 17408 3392 17460 3398
rect 17408 3334 17460 3340
rect 17420 3126 17448 3334
rect 17132 3120 17184 3126
rect 17132 3062 17184 3068
rect 17316 3120 17368 3126
rect 17316 3062 17368 3068
rect 17408 3120 17460 3126
rect 17408 3062 17460 3068
rect 17144 2854 17172 3062
rect 17408 2984 17460 2990
rect 17592 2984 17644 2990
rect 17460 2944 17592 2972
rect 17408 2926 17460 2932
rect 17592 2926 17644 2932
rect 17132 2848 17184 2854
rect 17696 2836 17724 3402
rect 17776 3120 17828 3126
rect 17776 3062 17828 3068
rect 17132 2790 17184 2796
rect 17604 2808 17724 2836
rect 17040 2508 17092 2514
rect 17040 2450 17092 2456
rect 16856 2440 16908 2446
rect 16856 2382 16908 2388
rect 16868 1766 16896 2382
rect 17040 2304 17092 2310
rect 17040 2246 17092 2252
rect 17132 2304 17184 2310
rect 17132 2246 17184 2252
rect 17408 2304 17460 2310
rect 17408 2246 17460 2252
rect 17052 2106 17080 2246
rect 17040 2100 17092 2106
rect 17040 2042 17092 2048
rect 16856 1760 16908 1766
rect 16856 1702 16908 1708
rect 17144 1426 17172 2246
rect 17420 1902 17448 2246
rect 17408 1896 17460 1902
rect 17408 1838 17460 1844
rect 17132 1420 17184 1426
rect 17132 1362 17184 1368
rect 17604 1358 17632 2808
rect 17788 2582 17816 3062
rect 17776 2576 17828 2582
rect 17776 2518 17828 2524
rect 17684 2508 17736 2514
rect 17684 2450 17736 2456
rect 17696 2417 17724 2450
rect 17682 2408 17738 2417
rect 17682 2343 17738 2352
rect 17866 2408 17922 2417
rect 17866 2343 17868 2352
rect 17920 2343 17922 2352
rect 17868 2314 17920 2320
rect 18064 2281 18092 3402
rect 18616 2990 18644 4558
rect 18708 4554 18736 5102
rect 18800 4570 18828 6190
rect 19064 6112 19116 6118
rect 19064 6054 19116 6060
rect 19076 5914 19104 6054
rect 19064 5908 19116 5914
rect 19064 5850 19116 5856
rect 19168 5778 19196 7806
rect 19260 7449 19288 8871
rect 19944 8894 20024 8900
rect 19892 8842 19944 8848
rect 19800 8832 19852 8838
rect 19800 8774 19852 8780
rect 19364 8732 19740 8741
rect 19420 8730 19444 8732
rect 19500 8730 19524 8732
rect 19580 8730 19604 8732
rect 19660 8730 19684 8732
rect 19420 8678 19430 8730
rect 19674 8678 19684 8730
rect 19420 8676 19444 8678
rect 19500 8676 19524 8678
rect 19580 8676 19604 8678
rect 19660 8676 19684 8678
rect 19364 8667 19740 8676
rect 19812 8106 19840 8774
rect 20088 8378 20116 9318
rect 19996 8350 20116 8378
rect 19892 8288 19944 8294
rect 19892 8230 19944 8236
rect 19628 8078 19840 8106
rect 19628 7954 19656 8078
rect 19616 7948 19668 7954
rect 19616 7890 19668 7896
rect 19708 7948 19760 7954
rect 19760 7908 19840 7936
rect 19708 7890 19760 7896
rect 19364 7644 19740 7653
rect 19420 7642 19444 7644
rect 19500 7642 19524 7644
rect 19580 7642 19604 7644
rect 19660 7642 19684 7644
rect 19420 7590 19430 7642
rect 19674 7590 19684 7642
rect 19420 7588 19444 7590
rect 19500 7588 19524 7590
rect 19580 7588 19604 7590
rect 19660 7588 19684 7590
rect 19364 7579 19740 7588
rect 19812 7546 19840 7908
rect 19904 7750 19932 8230
rect 19892 7744 19944 7750
rect 19892 7686 19944 7692
rect 19800 7540 19852 7546
rect 19800 7482 19852 7488
rect 19246 7440 19302 7449
rect 19246 7375 19302 7384
rect 19614 7440 19670 7449
rect 19614 7375 19670 7384
rect 19628 7342 19656 7375
rect 19616 7336 19668 7342
rect 19616 7278 19668 7284
rect 19800 7268 19852 7274
rect 19800 7210 19852 7216
rect 19812 7002 19840 7210
rect 19800 6996 19852 7002
rect 19800 6938 19852 6944
rect 19904 6934 19932 7686
rect 19892 6928 19944 6934
rect 19798 6896 19854 6905
rect 19708 6860 19760 6866
rect 19892 6870 19944 6876
rect 19798 6831 19854 6840
rect 19708 6802 19760 6808
rect 19720 6769 19748 6802
rect 19812 6798 19840 6831
rect 19800 6792 19852 6798
rect 19706 6760 19762 6769
rect 19800 6734 19852 6740
rect 19706 6695 19762 6704
rect 19892 6656 19944 6662
rect 19892 6598 19944 6604
rect 19364 6556 19740 6565
rect 19420 6554 19444 6556
rect 19500 6554 19524 6556
rect 19580 6554 19604 6556
rect 19660 6554 19684 6556
rect 19420 6502 19430 6554
rect 19674 6502 19684 6554
rect 19420 6500 19444 6502
rect 19500 6500 19524 6502
rect 19580 6500 19604 6502
rect 19660 6500 19684 6502
rect 19364 6491 19740 6500
rect 19904 6458 19932 6598
rect 19892 6452 19944 6458
rect 19892 6394 19944 6400
rect 19430 6352 19486 6361
rect 19430 6287 19486 6296
rect 19444 5778 19472 6287
rect 19800 6112 19852 6118
rect 19800 6054 19852 6060
rect 19522 5808 19578 5817
rect 19156 5772 19208 5778
rect 19156 5714 19208 5720
rect 19432 5772 19484 5778
rect 19522 5743 19524 5752
rect 19432 5714 19484 5720
rect 19576 5743 19578 5752
rect 19524 5714 19576 5720
rect 18880 5568 18932 5574
rect 18880 5510 18932 5516
rect 18892 4690 18920 5510
rect 19064 5364 19116 5370
rect 19064 5306 19116 5312
rect 19076 5234 19104 5306
rect 19064 5228 19116 5234
rect 19064 5170 19116 5176
rect 18972 5160 19024 5166
rect 19168 5137 19196 5714
rect 19364 5468 19740 5477
rect 19420 5466 19444 5468
rect 19500 5466 19524 5468
rect 19580 5466 19604 5468
rect 19660 5466 19684 5468
rect 19420 5414 19430 5466
rect 19674 5414 19684 5466
rect 19420 5412 19444 5414
rect 19500 5412 19524 5414
rect 19580 5412 19604 5414
rect 19660 5412 19684 5414
rect 19364 5403 19740 5412
rect 19812 5370 19840 6054
rect 19800 5364 19852 5370
rect 19800 5306 19852 5312
rect 19706 5264 19762 5273
rect 19706 5199 19762 5208
rect 18972 5102 19024 5108
rect 19154 5128 19210 5137
rect 18984 4826 19012 5102
rect 19064 5092 19116 5098
rect 19154 5063 19210 5072
rect 19064 5034 19116 5040
rect 18972 4820 19024 4826
rect 18972 4762 19024 4768
rect 18880 4684 18932 4690
rect 18880 4626 18932 4632
rect 18696 4548 18748 4554
rect 18800 4542 18920 4570
rect 18696 4490 18748 4496
rect 18788 4480 18840 4486
rect 18788 4422 18840 4428
rect 18604 2984 18656 2990
rect 18604 2926 18656 2932
rect 18510 2680 18566 2689
rect 18510 2615 18566 2624
rect 18050 2272 18106 2281
rect 18050 2207 18106 2216
rect 17774 2000 17830 2009
rect 18064 1970 18092 2207
rect 17774 1935 17830 1944
rect 18052 1964 18104 1970
rect 17788 1902 17816 1935
rect 18052 1906 18104 1912
rect 17776 1896 17828 1902
rect 17776 1838 17828 1844
rect 18328 1828 18380 1834
rect 18328 1770 18380 1776
rect 16856 1352 16908 1358
rect 16856 1294 16908 1300
rect 17592 1352 17644 1358
rect 17592 1294 17644 1300
rect 16868 1193 16896 1294
rect 16854 1184 16910 1193
rect 16854 1119 16910 1128
rect 16212 808 16264 814
rect 16212 750 16264 756
rect 16764 808 16816 814
rect 16764 750 16816 756
rect 16364 572 16740 581
rect 16420 570 16444 572
rect 16500 570 16524 572
rect 16580 570 16604 572
rect 16660 570 16684 572
rect 16420 518 16430 570
rect 16674 518 16684 570
rect 16420 516 16444 518
rect 16500 516 16524 518
rect 16580 516 16604 518
rect 16660 516 16684 518
rect 16364 507 16740 516
rect 15568 332 15620 338
rect 15568 274 15620 280
rect 16868 270 16896 1119
rect 16856 264 16908 270
rect 16856 206 16908 212
rect 15200 128 15252 134
rect 17604 105 17632 1294
rect 18340 1222 18368 1770
rect 18524 1562 18552 2615
rect 18800 2514 18828 4422
rect 18892 3670 18920 4542
rect 19076 4321 19104 5034
rect 19720 5030 19748 5199
rect 19156 5024 19208 5030
rect 19156 4966 19208 4972
rect 19708 5024 19760 5030
rect 19708 4966 19760 4972
rect 19062 4312 19118 4321
rect 19062 4247 19118 4256
rect 18880 3664 18932 3670
rect 18880 3606 18932 3612
rect 18880 3528 18932 3534
rect 18878 3496 18880 3505
rect 18932 3496 18934 3505
rect 18878 3431 18934 3440
rect 19168 2514 19196 4966
rect 19708 4820 19760 4826
rect 19708 4762 19760 4768
rect 19720 4570 19748 4762
rect 19812 4690 19840 5306
rect 19904 5166 19932 6394
rect 19996 5846 20024 8350
rect 20076 8288 20128 8294
rect 20076 8230 20128 8236
rect 20088 7818 20116 8230
rect 20180 8090 20208 9930
rect 20168 8084 20220 8090
rect 20168 8026 20220 8032
rect 20076 7812 20128 7818
rect 20076 7754 20128 7760
rect 20088 7410 20116 7754
rect 20168 7744 20220 7750
rect 20168 7686 20220 7692
rect 20180 7478 20208 7686
rect 20168 7472 20220 7478
rect 20168 7414 20220 7420
rect 20076 7404 20128 7410
rect 20076 7346 20128 7352
rect 20168 7200 20220 7206
rect 20168 7142 20220 7148
rect 20180 6798 20208 7142
rect 20272 7002 20300 9998
rect 20364 9926 20392 12294
rect 20456 12238 20484 12786
rect 20444 12232 20496 12238
rect 20444 12174 20496 12180
rect 20548 12084 20576 13246
rect 20812 13194 20864 13200
rect 20720 13184 20772 13190
rect 20720 13126 20772 13132
rect 20732 12434 20760 13126
rect 20810 12880 20866 12889
rect 20810 12815 20866 12824
rect 20824 12782 20852 12815
rect 20812 12776 20864 12782
rect 20812 12718 20864 12724
rect 20732 12406 20852 12434
rect 20824 12306 20852 12406
rect 20812 12300 20864 12306
rect 20812 12242 20864 12248
rect 20628 12232 20680 12238
rect 20626 12200 20628 12209
rect 20680 12200 20682 12209
rect 20626 12135 20682 12144
rect 20456 12056 20576 12084
rect 20352 9920 20404 9926
rect 20352 9862 20404 9868
rect 20364 9518 20392 9862
rect 20456 9674 20484 12056
rect 20640 11762 20668 12135
rect 20628 11756 20680 11762
rect 20628 11698 20680 11704
rect 20628 11620 20680 11626
rect 20628 11562 20680 11568
rect 20640 11218 20668 11562
rect 20720 11552 20772 11558
rect 20720 11494 20772 11500
rect 20628 11212 20680 11218
rect 20548 11172 20628 11200
rect 20548 10606 20576 11172
rect 20628 11154 20680 11160
rect 20732 10606 20760 11494
rect 20536 10600 20588 10606
rect 20536 10542 20588 10548
rect 20720 10600 20772 10606
rect 20720 10542 20772 10548
rect 20732 10130 20760 10542
rect 20536 10124 20588 10130
rect 20720 10124 20772 10130
rect 20588 10084 20668 10112
rect 20536 10066 20588 10072
rect 20640 9722 20668 10084
rect 20720 10066 20772 10072
rect 20628 9716 20680 9722
rect 20456 9646 20576 9674
rect 20628 9658 20680 9664
rect 20352 9512 20404 9518
rect 20352 9454 20404 9460
rect 20444 9376 20496 9382
rect 20350 9344 20406 9353
rect 20444 9318 20496 9324
rect 20350 9279 20406 9288
rect 20364 8906 20392 9279
rect 20352 8900 20404 8906
rect 20352 8842 20404 8848
rect 20352 8628 20404 8634
rect 20352 8570 20404 8576
rect 20364 8498 20392 8570
rect 20456 8514 20484 9318
rect 20352 8492 20404 8498
rect 20352 8434 20404 8440
rect 20455 8486 20484 8514
rect 20352 8288 20404 8294
rect 20455 8276 20483 8486
rect 20548 8294 20576 9646
rect 20720 8900 20772 8906
rect 20720 8842 20772 8848
rect 20628 8832 20680 8838
rect 20628 8774 20680 8780
rect 20536 8288 20588 8294
rect 20455 8248 20484 8276
rect 20352 8230 20404 8236
rect 20260 6996 20312 7002
rect 20260 6938 20312 6944
rect 20258 6896 20314 6905
rect 20258 6831 20260 6840
rect 20312 6831 20314 6840
rect 20260 6802 20312 6808
rect 20168 6792 20220 6798
rect 20168 6734 20220 6740
rect 20168 6180 20220 6186
rect 20168 6122 20220 6128
rect 19984 5840 20036 5846
rect 19984 5782 20036 5788
rect 19996 5234 20024 5782
rect 20180 5778 20208 6122
rect 20168 5772 20220 5778
rect 20168 5714 20220 5720
rect 20074 5672 20130 5681
rect 20074 5607 20130 5616
rect 19984 5228 20036 5234
rect 19984 5170 20036 5176
rect 19892 5160 19944 5166
rect 19892 5102 19944 5108
rect 19904 4826 19932 5102
rect 19984 5024 20036 5030
rect 19984 4966 20036 4972
rect 19892 4820 19944 4826
rect 19892 4762 19944 4768
rect 19800 4684 19852 4690
rect 19852 4644 19932 4672
rect 19800 4626 19852 4632
rect 19720 4542 19840 4570
rect 19364 4380 19740 4389
rect 19420 4378 19444 4380
rect 19500 4378 19524 4380
rect 19580 4378 19604 4380
rect 19660 4378 19684 4380
rect 19420 4326 19430 4378
rect 19674 4326 19684 4378
rect 19420 4324 19444 4326
rect 19500 4324 19524 4326
rect 19580 4324 19604 4326
rect 19660 4324 19684 4326
rect 19364 4315 19740 4324
rect 19340 4072 19392 4078
rect 19340 4014 19392 4020
rect 19352 3942 19380 4014
rect 19340 3936 19392 3942
rect 19340 3878 19392 3884
rect 19812 3738 19840 4542
rect 19904 4146 19932 4644
rect 19892 4140 19944 4146
rect 19892 4082 19944 4088
rect 19996 4049 20024 4966
rect 19982 4040 20038 4049
rect 19982 3975 20038 3984
rect 19800 3732 19852 3738
rect 19800 3674 19852 3680
rect 19522 3632 19578 3641
rect 19890 3632 19946 3641
rect 19522 3567 19524 3576
rect 19576 3567 19578 3576
rect 19800 3596 19852 3602
rect 19524 3538 19576 3544
rect 19890 3567 19892 3576
rect 19800 3538 19852 3544
rect 19944 3567 19946 3576
rect 19892 3538 19944 3544
rect 19340 3528 19392 3534
rect 19338 3496 19340 3505
rect 19392 3496 19394 3505
rect 19338 3431 19394 3440
rect 19364 3292 19740 3301
rect 19420 3290 19444 3292
rect 19500 3290 19524 3292
rect 19580 3290 19604 3292
rect 19660 3290 19684 3292
rect 19420 3238 19430 3290
rect 19674 3238 19684 3290
rect 19420 3236 19444 3238
rect 19500 3236 19524 3238
rect 19580 3236 19604 3238
rect 19660 3236 19684 3238
rect 19364 3227 19740 3236
rect 19812 3176 19840 3538
rect 19892 3188 19944 3194
rect 19812 3148 19892 3176
rect 19812 3058 19840 3148
rect 19892 3130 19944 3136
rect 19800 3052 19852 3058
rect 19800 2994 19852 3000
rect 19996 2990 20024 3975
rect 20088 3942 20116 5607
rect 20180 5370 20208 5714
rect 20260 5704 20312 5710
rect 20260 5646 20312 5652
rect 20364 5658 20392 8230
rect 20456 6304 20484 8248
rect 20536 8230 20588 8236
rect 20536 8084 20588 8090
rect 20536 8026 20588 8032
rect 20548 6866 20576 8026
rect 20536 6860 20588 6866
rect 20536 6802 20588 6808
rect 20536 6656 20588 6662
rect 20536 6598 20588 6604
rect 20548 6458 20576 6598
rect 20536 6452 20588 6458
rect 20536 6394 20588 6400
rect 20536 6316 20588 6322
rect 20456 6276 20536 6304
rect 20536 6258 20588 6264
rect 20640 6186 20668 8774
rect 20732 8430 20760 8842
rect 20720 8424 20772 8430
rect 20720 8366 20772 8372
rect 20720 8288 20772 8294
rect 20720 8230 20772 8236
rect 20732 8022 20760 8230
rect 20720 8016 20772 8022
rect 20720 7958 20772 7964
rect 20732 6934 20760 7958
rect 20720 6928 20772 6934
rect 20720 6870 20772 6876
rect 20628 6180 20680 6186
rect 20628 6122 20680 6128
rect 20168 5364 20220 5370
rect 20168 5306 20220 5312
rect 20272 5302 20300 5646
rect 20364 5630 20576 5658
rect 20352 5568 20404 5574
rect 20352 5510 20404 5516
rect 20260 5296 20312 5302
rect 20260 5238 20312 5244
rect 20364 4078 20392 5510
rect 20444 4548 20496 4554
rect 20444 4490 20496 4496
rect 20456 4078 20484 4490
rect 20260 4072 20312 4078
rect 20258 4040 20260 4049
rect 20352 4072 20404 4078
rect 20312 4040 20314 4049
rect 20352 4014 20404 4020
rect 20444 4072 20496 4078
rect 20444 4014 20496 4020
rect 20258 3975 20314 3984
rect 20076 3936 20128 3942
rect 20076 3878 20128 3884
rect 20168 3936 20220 3942
rect 20168 3878 20220 3884
rect 20352 3936 20404 3942
rect 20352 3878 20404 3884
rect 20088 3534 20116 3878
rect 20180 3670 20208 3878
rect 20168 3664 20220 3670
rect 20168 3606 20220 3612
rect 20076 3528 20128 3534
rect 20076 3470 20128 3476
rect 20260 3460 20312 3466
rect 20260 3402 20312 3408
rect 20168 3392 20220 3398
rect 20168 3334 20220 3340
rect 19984 2984 20036 2990
rect 19984 2926 20036 2932
rect 19892 2848 19944 2854
rect 19892 2790 19944 2796
rect 19984 2848 20036 2854
rect 19984 2790 20036 2796
rect 18788 2508 18840 2514
rect 18788 2450 18840 2456
rect 19156 2508 19208 2514
rect 19156 2450 19208 2456
rect 19800 2372 19852 2378
rect 19800 2314 19852 2320
rect 18604 2304 18656 2310
rect 18604 2246 18656 2252
rect 18880 2304 18932 2310
rect 18880 2246 18932 2252
rect 18972 2304 19024 2310
rect 18972 2246 19024 2252
rect 18512 1556 18564 1562
rect 18512 1498 18564 1504
rect 18616 1426 18644 2246
rect 18694 2000 18750 2009
rect 18694 1935 18750 1944
rect 18708 1902 18736 1935
rect 18696 1896 18748 1902
rect 18696 1838 18748 1844
rect 18708 1562 18736 1838
rect 18696 1556 18748 1562
rect 18696 1498 18748 1504
rect 18604 1420 18656 1426
rect 18604 1362 18656 1368
rect 18604 1284 18656 1290
rect 18604 1226 18656 1232
rect 18696 1284 18748 1290
rect 18696 1226 18748 1232
rect 17684 1216 17736 1222
rect 17684 1158 17736 1164
rect 17776 1216 17828 1222
rect 17776 1158 17828 1164
rect 18328 1216 18380 1222
rect 18328 1158 18380 1164
rect 17696 882 17724 1158
rect 17684 876 17736 882
rect 17684 818 17736 824
rect 17684 672 17736 678
rect 17684 614 17736 620
rect 17696 406 17724 614
rect 17788 474 17816 1158
rect 17866 1048 17922 1057
rect 17866 983 17922 992
rect 17880 814 17908 983
rect 17868 808 17920 814
rect 18616 785 18644 1226
rect 17868 750 17920 756
rect 18602 776 18658 785
rect 18602 711 18658 720
rect 18144 672 18196 678
rect 18064 632 18144 660
rect 17776 468 17828 474
rect 17776 410 17828 416
rect 17868 468 17920 474
rect 17868 410 17920 416
rect 17684 400 17736 406
rect 17684 342 17736 348
rect 17880 241 17908 410
rect 18064 400 18092 632
rect 18144 614 18196 620
rect 18420 672 18472 678
rect 18420 614 18472 620
rect 18432 400 18460 614
rect 18708 474 18736 1226
rect 18788 740 18840 746
rect 18788 682 18840 688
rect 18696 468 18748 474
rect 18696 410 18748 416
rect 18800 400 18828 682
rect 17866 232 17922 241
rect 17866 167 17922 176
rect 15200 70 15252 76
rect 17590 96 17646 105
rect 17590 31 17646 40
rect 18050 0 18106 400
rect 18418 0 18474 400
rect 18786 0 18842 400
rect 18892 338 18920 2246
rect 18984 1834 19012 2246
rect 19364 2204 19740 2213
rect 19420 2202 19444 2204
rect 19500 2202 19524 2204
rect 19580 2202 19604 2204
rect 19660 2202 19684 2204
rect 19420 2150 19430 2202
rect 19674 2150 19684 2202
rect 19420 2148 19444 2150
rect 19500 2148 19524 2150
rect 19580 2148 19604 2150
rect 19660 2148 19684 2150
rect 19364 2139 19740 2148
rect 18972 1828 19024 1834
rect 18972 1770 19024 1776
rect 19248 1760 19300 1766
rect 19340 1760 19392 1766
rect 19248 1702 19300 1708
rect 19338 1728 19340 1737
rect 19392 1728 19394 1737
rect 18972 1420 19024 1426
rect 18972 1362 19024 1368
rect 19064 1420 19116 1426
rect 19064 1362 19116 1368
rect 18880 332 18932 338
rect 18880 274 18932 280
rect 18984 202 19012 1362
rect 19076 1222 19104 1362
rect 19064 1216 19116 1222
rect 19064 1158 19116 1164
rect 19076 814 19104 1158
rect 19156 944 19208 950
rect 19156 886 19208 892
rect 19064 808 19116 814
rect 19064 750 19116 756
rect 19168 400 19196 886
rect 19260 814 19288 1702
rect 19338 1663 19394 1672
rect 19706 1456 19762 1465
rect 19812 1426 19840 2314
rect 19904 2281 19932 2790
rect 19890 2272 19946 2281
rect 19890 2207 19946 2216
rect 19996 2038 20024 2790
rect 20074 2408 20130 2417
rect 20074 2343 20130 2352
rect 20088 2106 20116 2343
rect 20076 2100 20128 2106
rect 20076 2042 20128 2048
rect 19984 2032 20036 2038
rect 19984 1974 20036 1980
rect 19892 1760 19944 1766
rect 19892 1702 19944 1708
rect 19984 1760 20036 1766
rect 19984 1702 20036 1708
rect 19904 1562 19932 1702
rect 19892 1556 19944 1562
rect 19892 1498 19944 1504
rect 19706 1391 19708 1400
rect 19760 1391 19762 1400
rect 19800 1420 19852 1426
rect 19708 1362 19760 1368
rect 19800 1362 19852 1368
rect 19798 1320 19854 1329
rect 19798 1255 19854 1264
rect 19892 1284 19944 1290
rect 19364 1116 19740 1125
rect 19420 1114 19444 1116
rect 19500 1114 19524 1116
rect 19580 1114 19604 1116
rect 19660 1114 19684 1116
rect 19420 1062 19430 1114
rect 19674 1062 19684 1114
rect 19420 1060 19444 1062
rect 19500 1060 19524 1062
rect 19580 1060 19604 1062
rect 19660 1060 19684 1062
rect 19364 1051 19740 1060
rect 19812 950 19840 1255
rect 19892 1226 19944 1232
rect 19904 1057 19932 1226
rect 19890 1048 19946 1057
rect 19890 983 19946 992
rect 19800 944 19852 950
rect 19800 886 19852 892
rect 19996 882 20024 1702
rect 20074 1456 20130 1465
rect 20180 1442 20208 3334
rect 20272 2378 20300 3402
rect 20364 3097 20392 3878
rect 20456 3194 20484 4014
rect 20548 3924 20576 5630
rect 20720 5636 20772 5642
rect 20720 5578 20772 5584
rect 20732 5370 20760 5578
rect 20720 5364 20772 5370
rect 20720 5306 20772 5312
rect 20628 5024 20680 5030
rect 20628 4966 20680 4972
rect 20640 4690 20668 4966
rect 20628 4684 20680 4690
rect 20628 4626 20680 4632
rect 20628 4072 20680 4078
rect 20680 4032 20760 4060
rect 20628 4014 20680 4020
rect 20732 4026 20760 4032
rect 20824 4026 20852 12242
rect 20916 11694 20944 18022
rect 21100 16794 21128 18362
rect 21284 17338 21312 19343
rect 21376 19174 21404 19502
rect 21364 19168 21416 19174
rect 21364 19110 21416 19116
rect 21364 18352 21416 18358
rect 21364 18294 21416 18300
rect 21376 17746 21404 18294
rect 21468 18290 21496 20266
rect 21560 19310 21588 20334
rect 21652 19922 21680 20878
rect 21836 20534 21864 21383
rect 22008 21354 22060 21360
rect 21824 20528 21876 20534
rect 21824 20470 21876 20476
rect 21824 20392 21876 20398
rect 21824 20334 21876 20340
rect 21640 19916 21692 19922
rect 21640 19858 21692 19864
rect 21732 19916 21784 19922
rect 21732 19858 21784 19864
rect 21744 19378 21772 19858
rect 21836 19446 21864 20334
rect 21916 20256 21968 20262
rect 21916 20198 21968 20204
rect 21824 19440 21876 19446
rect 21824 19382 21876 19388
rect 21732 19372 21784 19378
rect 21732 19314 21784 19320
rect 21548 19304 21600 19310
rect 21548 19246 21600 19252
rect 21732 19236 21784 19242
rect 21732 19178 21784 19184
rect 21744 18970 21772 19178
rect 21732 18964 21784 18970
rect 21732 18906 21784 18912
rect 21732 18624 21784 18630
rect 21836 18601 21864 19382
rect 21732 18566 21784 18572
rect 21822 18592 21878 18601
rect 21456 18284 21508 18290
rect 21456 18226 21508 18232
rect 21456 18080 21508 18086
rect 21548 18080 21600 18086
rect 21456 18022 21508 18028
rect 21546 18048 21548 18057
rect 21600 18048 21602 18057
rect 21364 17740 21416 17746
rect 21364 17682 21416 17688
rect 21272 17332 21324 17338
rect 21272 17274 21324 17280
rect 21364 17264 21416 17270
rect 21364 17206 21416 17212
rect 21088 16788 21140 16794
rect 21088 16730 21140 16736
rect 21180 16788 21232 16794
rect 21180 16730 21232 16736
rect 21088 16652 21140 16658
rect 21088 16594 21140 16600
rect 21100 16454 21128 16594
rect 21088 16448 21140 16454
rect 21088 16390 21140 16396
rect 20996 16176 21048 16182
rect 20996 16118 21048 16124
rect 21008 12850 21036 16118
rect 21100 15570 21128 16390
rect 21192 16250 21220 16730
rect 21180 16244 21232 16250
rect 21180 16186 21232 16192
rect 21088 15564 21140 15570
rect 21088 15506 21140 15512
rect 21088 15428 21140 15434
rect 21088 15370 21140 15376
rect 21100 13190 21128 15370
rect 21192 14482 21220 16186
rect 21272 16176 21324 16182
rect 21272 16118 21324 16124
rect 21284 14618 21312 16118
rect 21376 16046 21404 17206
rect 21364 16040 21416 16046
rect 21364 15982 21416 15988
rect 21468 15314 21496 18022
rect 21546 17983 21602 17992
rect 21744 17746 21772 18566
rect 21822 18527 21878 18536
rect 21732 17740 21784 17746
rect 21732 17682 21784 17688
rect 21744 17134 21772 17682
rect 21732 17128 21784 17134
rect 21732 17070 21784 17076
rect 21744 16658 21772 17070
rect 21732 16652 21784 16658
rect 21732 16594 21784 16600
rect 21468 15286 21588 15314
rect 21364 14816 21416 14822
rect 21364 14758 21416 14764
rect 21272 14612 21324 14618
rect 21272 14554 21324 14560
rect 21376 14550 21404 14758
rect 21364 14544 21416 14550
rect 21364 14486 21416 14492
rect 21180 14476 21232 14482
rect 21180 14418 21232 14424
rect 21180 13728 21232 13734
rect 21180 13670 21232 13676
rect 21088 13184 21140 13190
rect 21088 13126 21140 13132
rect 20996 12844 21048 12850
rect 20996 12786 21048 12792
rect 20904 11688 20956 11694
rect 20904 11630 20956 11636
rect 20916 11218 20944 11630
rect 20904 11212 20956 11218
rect 20904 11154 20956 11160
rect 20904 10464 20956 10470
rect 20904 10406 20956 10412
rect 20916 9994 20944 10406
rect 20904 9988 20956 9994
rect 20904 9930 20956 9936
rect 20916 6118 20944 9930
rect 21008 9654 21036 12786
rect 21192 12288 21220 13670
rect 21456 12708 21508 12714
rect 21456 12650 21508 12656
rect 21272 12640 21324 12646
rect 21272 12582 21324 12588
rect 21284 12306 21312 12582
rect 21468 12442 21496 12650
rect 21456 12436 21508 12442
rect 21456 12378 21508 12384
rect 21100 12260 21220 12288
rect 21272 12300 21324 12306
rect 21100 11830 21128 12260
rect 21272 12242 21324 12248
rect 21560 12186 21588 15286
rect 21640 14272 21692 14278
rect 21640 14214 21692 14220
rect 21652 14074 21680 14214
rect 21640 14068 21692 14074
rect 21640 14010 21692 14016
rect 21652 13870 21680 14010
rect 21640 13864 21692 13870
rect 21640 13806 21692 13812
rect 21744 12714 21772 16594
rect 21928 16046 21956 20198
rect 22020 19514 22048 21354
rect 22112 20806 22140 23600
rect 22664 23582 22784 23600
rect 22364 23420 22740 23429
rect 22420 23418 22444 23420
rect 22500 23418 22524 23420
rect 22580 23418 22604 23420
rect 22660 23418 22684 23420
rect 22420 23366 22430 23418
rect 22674 23366 22684 23418
rect 22420 23364 22444 23366
rect 22500 23364 22524 23366
rect 22580 23364 22604 23366
rect 22660 23364 22684 23366
rect 22364 23355 22740 23364
rect 22836 23112 22888 23118
rect 22836 23054 22888 23060
rect 22848 22574 22876 23054
rect 22192 22568 22244 22574
rect 22192 22510 22244 22516
rect 22836 22568 22888 22574
rect 22836 22510 22888 22516
rect 22204 21894 22232 22510
rect 22364 22332 22740 22341
rect 22420 22330 22444 22332
rect 22500 22330 22524 22332
rect 22580 22330 22604 22332
rect 22660 22330 22684 22332
rect 22420 22278 22430 22330
rect 22674 22278 22684 22330
rect 22420 22276 22444 22278
rect 22500 22276 22524 22278
rect 22580 22276 22604 22278
rect 22660 22276 22684 22278
rect 22364 22267 22740 22276
rect 22192 21888 22244 21894
rect 22192 21830 22244 21836
rect 22284 21888 22336 21894
rect 22284 21830 22336 21836
rect 22296 21536 22324 21830
rect 22848 21554 22876 22510
rect 22940 22166 22968 23718
rect 23202 23600 23258 24000
rect 23020 22500 23072 22506
rect 23020 22442 23072 22448
rect 22928 22160 22980 22166
rect 22928 22102 22980 22108
rect 22204 21508 22324 21536
rect 22836 21548 22888 21554
rect 22100 20800 22152 20806
rect 22100 20742 22152 20748
rect 22100 20528 22152 20534
rect 22100 20470 22152 20476
rect 22008 19508 22060 19514
rect 22008 19450 22060 19456
rect 22020 19417 22048 19450
rect 22006 19408 22062 19417
rect 22006 19343 22062 19352
rect 22112 19310 22140 20470
rect 22204 19961 22232 21508
rect 22888 21508 22968 21536
rect 22836 21490 22888 21496
rect 22284 21412 22336 21418
rect 22284 21354 22336 21360
rect 22296 20602 22324 21354
rect 22364 21244 22740 21253
rect 22420 21242 22444 21244
rect 22500 21242 22524 21244
rect 22580 21242 22604 21244
rect 22660 21242 22684 21244
rect 22420 21190 22430 21242
rect 22674 21190 22684 21242
rect 22420 21188 22444 21190
rect 22500 21188 22524 21190
rect 22580 21188 22604 21190
rect 22660 21188 22684 21190
rect 22364 21179 22740 21188
rect 22940 21010 22968 21508
rect 22744 21004 22796 21010
rect 22744 20946 22796 20952
rect 22928 21004 22980 21010
rect 22928 20946 22980 20952
rect 22376 20800 22428 20806
rect 22376 20742 22428 20748
rect 22284 20596 22336 20602
rect 22284 20538 22336 20544
rect 22388 20482 22416 20742
rect 22296 20454 22416 20482
rect 22560 20460 22612 20466
rect 22190 19952 22246 19961
rect 22190 19887 22246 19896
rect 22296 19334 22324 20454
rect 22560 20402 22612 20408
rect 22376 20392 22428 20398
rect 22374 20360 22376 20369
rect 22428 20360 22430 20369
rect 22572 20330 22600 20402
rect 22374 20295 22430 20304
rect 22560 20324 22612 20330
rect 22560 20266 22612 20272
rect 22756 20244 22784 20946
rect 23032 20890 23060 22442
rect 22940 20862 23060 20890
rect 22756 20216 22876 20244
rect 22364 20156 22740 20165
rect 22420 20154 22444 20156
rect 22500 20154 22524 20156
rect 22580 20154 22604 20156
rect 22660 20154 22684 20156
rect 22420 20102 22430 20154
rect 22674 20102 22684 20154
rect 22420 20100 22444 20102
rect 22500 20100 22524 20102
rect 22580 20100 22604 20102
rect 22660 20100 22684 20102
rect 22364 20091 22740 20100
rect 22296 19310 22508 19334
rect 22100 19304 22152 19310
rect 22296 19306 22520 19310
rect 22100 19246 22152 19252
rect 22468 19304 22520 19306
rect 22468 19246 22520 19252
rect 22008 19168 22060 19174
rect 22008 19110 22060 19116
rect 22020 18748 22048 19110
rect 22112 18902 22140 19246
rect 22192 19168 22244 19174
rect 22376 19168 22428 19174
rect 22244 19128 22376 19156
rect 22192 19110 22244 19116
rect 22376 19110 22428 19116
rect 22364 19068 22740 19077
rect 22420 19066 22444 19068
rect 22500 19066 22524 19068
rect 22580 19066 22604 19068
rect 22660 19066 22684 19068
rect 22420 19014 22430 19066
rect 22674 19014 22684 19066
rect 22420 19012 22444 19014
rect 22500 19012 22524 19014
rect 22580 19012 22604 19014
rect 22660 19012 22684 19014
rect 22364 19003 22740 19012
rect 22284 18964 22336 18970
rect 22284 18906 22336 18912
rect 22100 18896 22152 18902
rect 22100 18838 22152 18844
rect 22020 18720 22140 18748
rect 22006 18592 22062 18601
rect 22006 18527 22062 18536
rect 22020 17814 22048 18527
rect 22008 17808 22060 17814
rect 22008 17750 22060 17756
rect 22020 16182 22048 17750
rect 22112 16674 22140 18720
rect 22192 17876 22244 17882
rect 22192 17818 22244 17824
rect 22204 17134 22232 17818
rect 22192 17128 22244 17134
rect 22192 17070 22244 17076
rect 22204 16794 22232 17070
rect 22192 16788 22244 16794
rect 22192 16730 22244 16736
rect 22112 16646 22232 16674
rect 22008 16176 22060 16182
rect 22008 16118 22060 16124
rect 22204 16114 22232 16646
rect 22296 16250 22324 18906
rect 22364 17980 22740 17989
rect 22420 17978 22444 17980
rect 22500 17978 22524 17980
rect 22580 17978 22604 17980
rect 22660 17978 22684 17980
rect 22420 17926 22430 17978
rect 22674 17926 22684 17978
rect 22420 17924 22444 17926
rect 22500 17924 22524 17926
rect 22580 17924 22604 17926
rect 22660 17924 22684 17926
rect 22364 17915 22740 17924
rect 22364 16892 22740 16901
rect 22420 16890 22444 16892
rect 22500 16890 22524 16892
rect 22580 16890 22604 16892
rect 22660 16890 22684 16892
rect 22420 16838 22430 16890
rect 22674 16838 22684 16890
rect 22420 16836 22444 16838
rect 22500 16836 22524 16838
rect 22580 16836 22604 16838
rect 22660 16836 22684 16838
rect 22364 16827 22740 16836
rect 22744 16788 22796 16794
rect 22744 16730 22796 16736
rect 22376 16652 22428 16658
rect 22376 16594 22428 16600
rect 22284 16244 22336 16250
rect 22284 16186 22336 16192
rect 22100 16108 22152 16114
rect 22100 16050 22152 16056
rect 22192 16108 22244 16114
rect 22192 16050 22244 16056
rect 21916 16040 21968 16046
rect 21916 15982 21968 15988
rect 22008 15972 22060 15978
rect 22008 15914 22060 15920
rect 21824 15904 21876 15910
rect 21824 15846 21876 15852
rect 21836 15570 21864 15846
rect 22020 15570 22048 15914
rect 22112 15570 22140 16050
rect 22388 16046 22416 16594
rect 22756 16046 22784 16730
rect 22376 16040 22428 16046
rect 22376 15982 22428 15988
rect 22744 16040 22796 16046
rect 22744 15982 22796 15988
rect 22364 15804 22740 15813
rect 22420 15802 22444 15804
rect 22500 15802 22524 15804
rect 22580 15802 22604 15804
rect 22660 15802 22684 15804
rect 22420 15750 22430 15802
rect 22674 15750 22684 15802
rect 22420 15748 22444 15750
rect 22500 15748 22524 15750
rect 22580 15748 22604 15750
rect 22660 15748 22684 15750
rect 22364 15739 22740 15748
rect 22848 15706 22876 20216
rect 22940 18970 22968 20862
rect 23020 20256 23072 20262
rect 23020 20198 23072 20204
rect 22928 18964 22980 18970
rect 22928 18906 22980 18912
rect 22928 18828 22980 18834
rect 22928 18770 22980 18776
rect 22940 16250 22968 18770
rect 22928 16244 22980 16250
rect 22928 16186 22980 16192
rect 22468 15700 22520 15706
rect 22468 15642 22520 15648
rect 22836 15700 22888 15706
rect 22836 15642 22888 15648
rect 21824 15564 21876 15570
rect 21824 15506 21876 15512
rect 22008 15564 22060 15570
rect 22008 15506 22060 15512
rect 22100 15564 22152 15570
rect 22100 15506 22152 15512
rect 22284 15564 22336 15570
rect 22284 15506 22336 15512
rect 22112 15450 22140 15506
rect 22020 15422 22140 15450
rect 22296 15434 22324 15506
rect 22284 15428 22336 15434
rect 21824 14816 21876 14822
rect 21824 14758 21876 14764
rect 21732 12708 21784 12714
rect 21732 12650 21784 12656
rect 21744 12434 21772 12650
rect 21836 12646 21864 14758
rect 22020 14482 22048 15422
rect 22284 15370 22336 15376
rect 22480 14958 22508 15642
rect 23032 15570 23060 20198
rect 23112 19168 23164 19174
rect 23112 19110 23164 19116
rect 23124 16046 23152 19110
rect 23216 18737 23244 23600
rect 23388 23180 23440 23186
rect 23388 23122 23440 23128
rect 23296 20324 23348 20330
rect 23296 20266 23348 20272
rect 23202 18728 23258 18737
rect 23202 18663 23258 18672
rect 23308 17882 23336 20266
rect 23400 19990 23428 23122
rect 23480 20392 23532 20398
rect 23480 20334 23532 20340
rect 23388 19984 23440 19990
rect 23388 19926 23440 19932
rect 23400 18086 23428 19926
rect 23388 18080 23440 18086
rect 23388 18022 23440 18028
rect 23296 17876 23348 17882
rect 23296 17818 23348 17824
rect 23388 17332 23440 17338
rect 23388 17274 23440 17280
rect 23204 16788 23256 16794
rect 23204 16730 23256 16736
rect 23112 16040 23164 16046
rect 23112 15982 23164 15988
rect 23020 15564 23072 15570
rect 23020 15506 23072 15512
rect 22560 15360 22612 15366
rect 22560 15302 22612 15308
rect 22572 15026 22600 15302
rect 22560 15020 22612 15026
rect 22560 14962 22612 14968
rect 22284 14952 22336 14958
rect 22284 14894 22336 14900
rect 22468 14952 22520 14958
rect 22468 14894 22520 14900
rect 22296 14482 22324 14894
rect 22364 14716 22740 14725
rect 22420 14714 22444 14716
rect 22500 14714 22524 14716
rect 22580 14714 22604 14716
rect 22660 14714 22684 14716
rect 22420 14662 22430 14714
rect 22674 14662 22684 14714
rect 22420 14660 22444 14662
rect 22500 14660 22524 14662
rect 22580 14660 22604 14662
rect 22660 14660 22684 14662
rect 22364 14651 22740 14660
rect 21916 14476 21968 14482
rect 21916 14418 21968 14424
rect 22008 14476 22060 14482
rect 22008 14418 22060 14424
rect 22284 14476 22336 14482
rect 22284 14418 22336 14424
rect 21824 12640 21876 12646
rect 21824 12582 21876 12588
rect 21652 12406 21772 12434
rect 21652 12374 21680 12406
rect 21640 12368 21692 12374
rect 21640 12310 21692 12316
rect 21192 12158 21588 12186
rect 21088 11824 21140 11830
rect 21088 11766 21140 11772
rect 21088 11212 21140 11218
rect 21088 11154 21140 11160
rect 21100 10606 21128 11154
rect 21088 10600 21140 10606
rect 21088 10542 21140 10548
rect 20996 9648 21048 9654
rect 21088 9648 21140 9654
rect 20996 9590 21048 9596
rect 21086 9616 21088 9625
rect 21140 9616 21142 9625
rect 21086 9551 21142 9560
rect 21088 8832 21140 8838
rect 21088 8774 21140 8780
rect 21100 8634 21128 8774
rect 21192 8634 21220 12158
rect 21456 12096 21508 12102
rect 21456 12038 21508 12044
rect 21548 12096 21600 12102
rect 21548 12038 21600 12044
rect 21468 11694 21496 12038
rect 21560 11762 21588 12038
rect 21548 11756 21600 11762
rect 21548 11698 21600 11704
rect 21456 11688 21508 11694
rect 21456 11630 21508 11636
rect 21548 11620 21600 11626
rect 21548 11562 21600 11568
rect 21272 11280 21324 11286
rect 21272 11222 21324 11228
rect 21284 10266 21312 11222
rect 21560 11218 21588 11562
rect 21652 11218 21680 12310
rect 21732 12300 21784 12306
rect 21732 12242 21784 12248
rect 21744 11898 21772 12242
rect 21824 12164 21876 12170
rect 21824 12106 21876 12112
rect 21732 11892 21784 11898
rect 21732 11834 21784 11840
rect 21732 11552 21784 11558
rect 21732 11494 21784 11500
rect 21744 11286 21772 11494
rect 21732 11280 21784 11286
rect 21732 11222 21784 11228
rect 21548 11212 21600 11218
rect 21548 11154 21600 11160
rect 21640 11212 21692 11218
rect 21640 11154 21692 11160
rect 21272 10260 21324 10266
rect 21272 10202 21324 10208
rect 21456 10260 21508 10266
rect 21456 10202 21508 10208
rect 21284 10062 21312 10202
rect 21468 10169 21496 10202
rect 21560 10198 21588 11154
rect 21836 10674 21864 12106
rect 21824 10668 21876 10674
rect 21824 10610 21876 10616
rect 21730 10296 21786 10305
rect 21730 10231 21786 10240
rect 21548 10192 21600 10198
rect 21454 10160 21510 10169
rect 21548 10134 21600 10140
rect 21454 10095 21510 10104
rect 21272 10056 21324 10062
rect 21272 9998 21324 10004
rect 21284 9518 21312 9998
rect 21456 9988 21508 9994
rect 21456 9930 21508 9936
rect 21272 9512 21324 9518
rect 21272 9454 21324 9460
rect 21272 9376 21324 9382
rect 21272 9318 21324 9324
rect 21088 8628 21140 8634
rect 21008 8588 21088 8616
rect 21008 7750 21036 8588
rect 21088 8570 21140 8576
rect 21180 8628 21232 8634
rect 21180 8570 21232 8576
rect 21086 8528 21142 8537
rect 21086 8463 21142 8472
rect 21100 8294 21128 8463
rect 21088 8288 21140 8294
rect 21088 8230 21140 8236
rect 21192 8022 21220 8570
rect 21284 8430 21312 9318
rect 21468 9081 21496 9930
rect 21560 9926 21588 10134
rect 21548 9920 21600 9926
rect 21548 9862 21600 9868
rect 21744 9722 21772 10231
rect 21732 9716 21784 9722
rect 21732 9658 21784 9664
rect 21548 9648 21600 9654
rect 21928 9602 21956 14418
rect 22468 14272 22520 14278
rect 22468 14214 22520 14220
rect 22480 13870 22508 14214
rect 22468 13864 22520 13870
rect 22468 13806 22520 13812
rect 22364 13628 22740 13637
rect 22420 13626 22444 13628
rect 22500 13626 22524 13628
rect 22580 13626 22604 13628
rect 22660 13626 22684 13628
rect 22420 13574 22430 13626
rect 22674 13574 22684 13626
rect 22420 13572 22444 13574
rect 22500 13572 22524 13574
rect 22580 13572 22604 13574
rect 22660 13572 22684 13574
rect 22364 13563 22740 13572
rect 22100 12640 22152 12646
rect 22100 12582 22152 12588
rect 22112 11694 22140 12582
rect 22364 12540 22740 12549
rect 22420 12538 22444 12540
rect 22500 12538 22524 12540
rect 22580 12538 22604 12540
rect 22660 12538 22684 12540
rect 22420 12486 22430 12538
rect 22674 12486 22684 12538
rect 22420 12484 22444 12486
rect 22500 12484 22524 12486
rect 22580 12484 22604 12486
rect 22660 12484 22684 12486
rect 22364 12475 22740 12484
rect 22100 11688 22152 11694
rect 22100 11630 22152 11636
rect 22284 11688 22336 11694
rect 22284 11630 22336 11636
rect 22112 10810 22140 11630
rect 22192 11552 22244 11558
rect 22192 11494 22244 11500
rect 22204 11286 22232 11494
rect 22192 11280 22244 11286
rect 22192 11222 22244 11228
rect 22296 10810 22324 11630
rect 22364 11452 22740 11461
rect 22420 11450 22444 11452
rect 22500 11450 22524 11452
rect 22580 11450 22604 11452
rect 22660 11450 22684 11452
rect 22420 11398 22430 11450
rect 22674 11398 22684 11450
rect 22420 11396 22444 11398
rect 22500 11396 22524 11398
rect 22580 11396 22604 11398
rect 22660 11396 22684 11398
rect 22364 11387 22740 11396
rect 23020 11008 23072 11014
rect 23020 10950 23072 10956
rect 22100 10804 22152 10810
rect 22100 10746 22152 10752
rect 22284 10804 22336 10810
rect 22284 10746 22336 10752
rect 23032 10606 23060 10950
rect 23020 10600 23072 10606
rect 23020 10542 23072 10548
rect 22836 10464 22888 10470
rect 22836 10406 22888 10412
rect 22928 10464 22980 10470
rect 22928 10406 22980 10412
rect 22364 10364 22740 10373
rect 22420 10362 22444 10364
rect 22500 10362 22524 10364
rect 22580 10362 22604 10364
rect 22660 10362 22684 10364
rect 22420 10310 22430 10362
rect 22674 10310 22684 10362
rect 22420 10308 22444 10310
rect 22500 10308 22524 10310
rect 22580 10308 22604 10310
rect 22660 10308 22684 10310
rect 22364 10299 22740 10308
rect 22652 10192 22704 10198
rect 22652 10134 22704 10140
rect 22468 9988 22520 9994
rect 22468 9930 22520 9936
rect 21548 9590 21600 9596
rect 21454 9072 21510 9081
rect 21454 9007 21456 9016
rect 21508 9007 21510 9016
rect 21456 8978 21508 8984
rect 21272 8424 21324 8430
rect 21456 8424 21508 8430
rect 21324 8372 21456 8378
rect 21272 8366 21508 8372
rect 21284 8350 21496 8366
rect 21180 8016 21232 8022
rect 21100 7976 21180 8004
rect 20996 7744 21048 7750
rect 20996 7686 21048 7692
rect 20904 6112 20956 6118
rect 20904 6054 20956 6060
rect 20916 5778 20944 6054
rect 20904 5772 20956 5778
rect 20904 5714 20956 5720
rect 21100 5166 21128 7976
rect 21180 7958 21232 7964
rect 21560 7546 21588 9590
rect 21744 9574 21956 9602
rect 21744 9110 21772 9574
rect 22480 9518 22508 9930
rect 22664 9518 22692 10134
rect 22848 10010 22876 10406
rect 22940 10198 22968 10406
rect 22928 10192 22980 10198
rect 22928 10134 22980 10140
rect 23216 10130 23244 16730
rect 23400 10674 23428 17274
rect 23492 15978 23520 20334
rect 23480 15972 23532 15978
rect 23480 15914 23532 15920
rect 23388 10668 23440 10674
rect 23388 10610 23440 10616
rect 23204 10124 23256 10130
rect 23204 10066 23256 10072
rect 22848 9982 22968 10010
rect 22744 9920 22796 9926
rect 22796 9868 22876 9874
rect 22744 9862 22876 9868
rect 22756 9846 22876 9862
rect 22468 9512 22520 9518
rect 22468 9454 22520 9460
rect 22652 9512 22704 9518
rect 22652 9454 22704 9460
rect 21824 9376 21876 9382
rect 22480 9364 22508 9454
rect 22848 9450 22876 9846
rect 22940 9518 22968 9982
rect 22928 9512 22980 9518
rect 22928 9454 22980 9460
rect 22836 9444 22888 9450
rect 22836 9386 22888 9392
rect 21824 9318 21876 9324
rect 22296 9336 22508 9364
rect 21732 9104 21784 9110
rect 21732 9046 21784 9052
rect 21640 8288 21692 8294
rect 21640 8230 21692 8236
rect 21456 7540 21508 7546
rect 21456 7482 21508 7488
rect 21548 7540 21600 7546
rect 21548 7482 21600 7488
rect 21468 7274 21496 7482
rect 21546 7440 21602 7449
rect 21546 7375 21602 7384
rect 21456 7268 21508 7274
rect 21456 7210 21508 7216
rect 21560 7206 21588 7375
rect 21652 7274 21680 8230
rect 21732 7472 21784 7478
rect 21732 7414 21784 7420
rect 21640 7268 21692 7274
rect 21640 7210 21692 7216
rect 21548 7200 21600 7206
rect 21600 7148 21680 7154
rect 21548 7142 21680 7148
rect 21560 7126 21680 7142
rect 21548 6996 21600 7002
rect 21548 6938 21600 6944
rect 21456 6656 21508 6662
rect 21456 6598 21508 6604
rect 21180 6384 21232 6390
rect 21180 6326 21232 6332
rect 21192 5846 21220 6326
rect 21362 6216 21418 6225
rect 21362 6151 21418 6160
rect 21272 6112 21324 6118
rect 21272 6054 21324 6060
rect 21180 5840 21232 5846
rect 21180 5782 21232 5788
rect 21180 5568 21232 5574
rect 21180 5510 21232 5516
rect 21192 5166 21220 5510
rect 21088 5160 21140 5166
rect 21088 5102 21140 5108
rect 21180 5160 21232 5166
rect 21180 5102 21232 5108
rect 21100 4690 21128 5102
rect 21192 4758 21220 5102
rect 21180 4752 21232 4758
rect 21180 4694 21232 4700
rect 21088 4684 21140 4690
rect 21088 4626 21140 4632
rect 21088 4480 21140 4486
rect 21088 4422 21140 4428
rect 21100 4185 21128 4422
rect 21086 4176 21142 4185
rect 21086 4111 21088 4120
rect 21140 4111 21142 4120
rect 21088 4082 21140 4088
rect 21180 4072 21232 4078
rect 20732 3998 21036 4026
rect 21180 4014 21232 4020
rect 20904 3936 20956 3942
rect 20548 3896 20668 3924
rect 20536 3392 20588 3398
rect 20536 3334 20588 3340
rect 20548 3194 20576 3334
rect 20444 3188 20496 3194
rect 20444 3130 20496 3136
rect 20536 3188 20588 3194
rect 20536 3130 20588 3136
rect 20350 3088 20406 3097
rect 20640 3058 20668 3896
rect 20904 3878 20956 3884
rect 20916 3602 20944 3878
rect 20904 3596 20956 3602
rect 20904 3538 20956 3544
rect 20350 3023 20406 3032
rect 20628 3052 20680 3058
rect 20628 2994 20680 3000
rect 20916 2990 20944 3538
rect 21008 3058 21036 3998
rect 21192 3942 21220 4014
rect 21180 3936 21232 3942
rect 21180 3878 21232 3884
rect 21086 3632 21142 3641
rect 21086 3567 21142 3576
rect 21100 3534 21128 3567
rect 21088 3528 21140 3534
rect 21192 3505 21220 3878
rect 21088 3470 21140 3476
rect 21178 3496 21234 3505
rect 21178 3431 21234 3440
rect 21192 3398 21220 3431
rect 21180 3392 21232 3398
rect 21180 3334 21232 3340
rect 20996 3052 21048 3058
rect 20996 2994 21048 3000
rect 21284 2990 21312 6054
rect 21376 5098 21404 6151
rect 21468 5778 21496 6598
rect 21456 5772 21508 5778
rect 21456 5714 21508 5720
rect 21456 5364 21508 5370
rect 21456 5306 21508 5312
rect 21364 5092 21416 5098
rect 21364 5034 21416 5040
rect 21468 4078 21496 5306
rect 21560 5166 21588 6938
rect 21652 6866 21680 7126
rect 21744 6882 21772 7414
rect 21836 7342 21864 9318
rect 21916 9172 21968 9178
rect 21916 9114 21968 9120
rect 21928 8430 21956 9114
rect 22296 9110 22324 9336
rect 22364 9276 22740 9285
rect 22420 9274 22444 9276
rect 22500 9274 22524 9276
rect 22580 9274 22604 9276
rect 22660 9274 22684 9276
rect 22420 9222 22430 9274
rect 22674 9222 22684 9274
rect 22420 9220 22444 9222
rect 22500 9220 22524 9222
rect 22580 9220 22604 9222
rect 22660 9220 22684 9222
rect 22364 9211 22740 9220
rect 22652 9172 22704 9178
rect 22652 9114 22704 9120
rect 22284 9104 22336 9110
rect 22284 9046 22336 9052
rect 22664 9042 22692 9114
rect 22100 9036 22152 9042
rect 22100 8978 22152 8984
rect 22652 9036 22704 9042
rect 22652 8978 22704 8984
rect 22008 8560 22060 8566
rect 22008 8502 22060 8508
rect 21916 8424 21968 8430
rect 21916 8366 21968 8372
rect 21916 8288 21968 8294
rect 21916 8230 21968 8236
rect 21928 7954 21956 8230
rect 21916 7948 21968 7954
rect 21916 7890 21968 7896
rect 21928 7342 21956 7890
rect 21824 7336 21876 7342
rect 21824 7278 21876 7284
rect 21916 7336 21968 7342
rect 21916 7278 21968 7284
rect 21914 6896 21970 6905
rect 21640 6860 21692 6866
rect 21744 6854 21864 6882
rect 21640 6802 21692 6808
rect 21836 6662 21864 6854
rect 22020 6866 22048 8502
rect 22112 8412 22140 8978
rect 22192 8424 22244 8430
rect 22112 8384 22192 8412
rect 22848 8401 22876 9386
rect 22940 9178 22968 9454
rect 22928 9172 22980 9178
rect 22928 9114 22980 9120
rect 22192 8366 22244 8372
rect 22834 8392 22890 8401
rect 22834 8327 22890 8336
rect 22364 8188 22740 8197
rect 22420 8186 22444 8188
rect 22500 8186 22524 8188
rect 22580 8186 22604 8188
rect 22660 8186 22684 8188
rect 22420 8134 22430 8186
rect 22674 8134 22684 8186
rect 22420 8132 22444 8134
rect 22500 8132 22524 8134
rect 22580 8132 22604 8134
rect 22660 8132 22684 8134
rect 22364 8123 22740 8132
rect 22284 7744 22336 7750
rect 22284 7686 22336 7692
rect 22296 7410 22324 7686
rect 22284 7404 22336 7410
rect 22284 7346 22336 7352
rect 22100 7268 22152 7274
rect 22100 7210 22152 7216
rect 22112 6905 22140 7210
rect 22364 7100 22740 7109
rect 22420 7098 22444 7100
rect 22500 7098 22524 7100
rect 22580 7098 22604 7100
rect 22660 7098 22684 7100
rect 22420 7046 22430 7098
rect 22674 7046 22684 7098
rect 22420 7044 22444 7046
rect 22500 7044 22524 7046
rect 22580 7044 22604 7046
rect 22660 7044 22684 7046
rect 22364 7035 22740 7044
rect 22098 6896 22154 6905
rect 21914 6831 21970 6840
rect 22008 6860 22060 6866
rect 21928 6730 21956 6831
rect 22098 6831 22154 6840
rect 22008 6802 22060 6808
rect 21916 6724 21968 6730
rect 21916 6666 21968 6672
rect 21824 6656 21876 6662
rect 21824 6598 21876 6604
rect 21914 6624 21970 6633
rect 21914 6559 21970 6568
rect 21640 5772 21692 5778
rect 21640 5714 21692 5720
rect 21548 5160 21600 5166
rect 21548 5102 21600 5108
rect 21652 4690 21680 5714
rect 21732 5092 21784 5098
rect 21732 5034 21784 5040
rect 21744 4758 21772 5034
rect 21928 4826 21956 6559
rect 22112 5658 22140 6831
rect 22192 6112 22244 6118
rect 22192 6054 22244 6060
rect 22284 6112 22336 6118
rect 22284 6054 22336 6060
rect 22204 5846 22232 6054
rect 22296 5914 22324 6054
rect 22364 6012 22740 6021
rect 22420 6010 22444 6012
rect 22500 6010 22524 6012
rect 22580 6010 22604 6012
rect 22660 6010 22684 6012
rect 22420 5958 22430 6010
rect 22674 5958 22684 6010
rect 22420 5956 22444 5958
rect 22500 5956 22524 5958
rect 22580 5956 22604 5958
rect 22660 5956 22684 5958
rect 22364 5947 22740 5956
rect 22284 5908 22336 5914
rect 22284 5850 22336 5856
rect 22192 5840 22244 5846
rect 22192 5782 22244 5788
rect 22112 5630 22232 5658
rect 22008 5568 22060 5574
rect 22008 5510 22060 5516
rect 22020 5370 22048 5510
rect 22008 5364 22060 5370
rect 22008 5306 22060 5312
rect 21824 4820 21876 4826
rect 21824 4762 21876 4768
rect 21916 4820 21968 4826
rect 21916 4762 21968 4768
rect 21732 4752 21784 4758
rect 21732 4694 21784 4700
rect 21548 4684 21600 4690
rect 21548 4626 21600 4632
rect 21640 4684 21692 4690
rect 21640 4626 21692 4632
rect 21560 4282 21588 4626
rect 21640 4480 21692 4486
rect 21640 4422 21692 4428
rect 21548 4276 21600 4282
rect 21548 4218 21600 4224
rect 21364 4072 21416 4078
rect 21364 4014 21416 4020
rect 21456 4072 21508 4078
rect 21456 4014 21508 4020
rect 21376 3738 21404 4014
rect 21364 3732 21416 3738
rect 21364 3674 21416 3680
rect 20904 2984 20956 2990
rect 20904 2926 20956 2932
rect 21272 2984 21324 2990
rect 21272 2926 21324 2932
rect 20812 2916 20864 2922
rect 20812 2858 20864 2864
rect 20824 2774 20852 2858
rect 20904 2848 20956 2854
rect 20904 2790 20956 2796
rect 21456 2848 21508 2854
rect 21456 2790 21508 2796
rect 20732 2746 20852 2774
rect 20732 2514 20760 2746
rect 20720 2508 20772 2514
rect 20720 2450 20772 2456
rect 20260 2372 20312 2378
rect 20260 2314 20312 2320
rect 20272 1970 20300 2314
rect 20444 2304 20496 2310
rect 20444 2246 20496 2252
rect 20260 1964 20312 1970
rect 20260 1906 20312 1912
rect 20456 1873 20484 2246
rect 20442 1864 20498 1873
rect 20442 1799 20498 1808
rect 20350 1728 20406 1737
rect 20350 1663 20406 1672
rect 20130 1414 20208 1442
rect 20364 1426 20392 1663
rect 20732 1494 20760 2450
rect 20812 2440 20864 2446
rect 20812 2382 20864 2388
rect 20824 2310 20852 2382
rect 20812 2304 20864 2310
rect 20812 2246 20864 2252
rect 20824 1902 20852 2246
rect 20812 1896 20864 1902
rect 20812 1838 20864 1844
rect 20720 1488 20772 1494
rect 20720 1430 20772 1436
rect 20824 1426 20852 1838
rect 20352 1420 20404 1426
rect 20074 1391 20130 1400
rect 20088 1358 20116 1391
rect 20352 1362 20404 1368
rect 20812 1420 20864 1426
rect 20812 1362 20864 1368
rect 20076 1352 20128 1358
rect 20444 1352 20496 1358
rect 20076 1294 20128 1300
rect 20166 1320 20222 1329
rect 20166 1255 20222 1264
rect 20272 1300 20444 1306
rect 20628 1352 20680 1358
rect 20272 1294 20496 1300
rect 20626 1320 20628 1329
rect 20680 1320 20682 1329
rect 20916 1306 20944 2790
rect 21468 2582 21496 2790
rect 21456 2576 21508 2582
rect 21456 2518 21508 2524
rect 21652 2514 21680 4422
rect 21732 3392 21784 3398
rect 21732 3334 21784 3340
rect 21640 2508 21692 2514
rect 21640 2450 21692 2456
rect 21364 2304 21416 2310
rect 21364 2246 21416 2252
rect 21376 1902 21404 2246
rect 21744 1902 21772 3334
rect 21836 2990 21864 4762
rect 22008 4616 22060 4622
rect 22008 4558 22060 4564
rect 22020 4078 22048 4558
rect 22100 4480 22152 4486
rect 22100 4422 22152 4428
rect 22112 4078 22140 4422
rect 21916 4072 21968 4078
rect 21916 4014 21968 4020
rect 22008 4072 22060 4078
rect 22008 4014 22060 4020
rect 22100 4072 22152 4078
rect 22100 4014 22152 4020
rect 21928 3602 21956 4014
rect 21916 3596 21968 3602
rect 21916 3538 21968 3544
rect 21916 3120 21968 3126
rect 21916 3062 21968 3068
rect 21824 2984 21876 2990
rect 21824 2926 21876 2932
rect 21824 2848 21876 2854
rect 21824 2790 21876 2796
rect 21836 2689 21864 2790
rect 21822 2680 21878 2689
rect 21822 2615 21878 2624
rect 21928 2446 21956 3062
rect 22020 3058 22048 4014
rect 22204 4010 22232 5630
rect 22284 5228 22336 5234
rect 22284 5170 22336 5176
rect 22296 4690 22324 5170
rect 22364 4924 22740 4933
rect 22420 4922 22444 4924
rect 22500 4922 22524 4924
rect 22580 4922 22604 4924
rect 22660 4922 22684 4924
rect 22420 4870 22430 4922
rect 22674 4870 22684 4922
rect 22420 4868 22444 4870
rect 22500 4868 22524 4870
rect 22580 4868 22604 4870
rect 22660 4868 22684 4870
rect 22364 4859 22740 4868
rect 22284 4684 22336 4690
rect 22284 4626 22336 4632
rect 23400 4622 23428 10610
rect 23388 4616 23440 4622
rect 23388 4558 23440 4564
rect 22284 4548 22336 4554
rect 22284 4490 22336 4496
rect 22192 4004 22244 4010
rect 22192 3946 22244 3952
rect 22296 3670 22324 4490
rect 22928 4208 22980 4214
rect 22928 4150 22980 4156
rect 22836 3936 22888 3942
rect 22836 3878 22888 3884
rect 22364 3836 22740 3845
rect 22420 3834 22444 3836
rect 22500 3834 22524 3836
rect 22580 3834 22604 3836
rect 22660 3834 22684 3836
rect 22420 3782 22430 3834
rect 22674 3782 22684 3834
rect 22420 3780 22444 3782
rect 22500 3780 22524 3782
rect 22580 3780 22604 3782
rect 22660 3780 22684 3782
rect 22364 3771 22740 3780
rect 22284 3664 22336 3670
rect 22284 3606 22336 3612
rect 22284 3392 22336 3398
rect 22284 3334 22336 3340
rect 22744 3392 22796 3398
rect 22744 3334 22796 3340
rect 22008 3052 22060 3058
rect 22008 2994 22060 3000
rect 22192 2508 22244 2514
rect 22192 2450 22244 2456
rect 21916 2440 21968 2446
rect 22204 2417 22232 2450
rect 21916 2382 21968 2388
rect 22190 2408 22246 2417
rect 22190 2343 22246 2352
rect 21916 2304 21968 2310
rect 21916 2246 21968 2252
rect 22100 2304 22152 2310
rect 22100 2246 22152 2252
rect 21364 1896 21416 1902
rect 21364 1838 21416 1844
rect 21548 1896 21600 1902
rect 21548 1838 21600 1844
rect 21732 1896 21784 1902
rect 21732 1838 21784 1844
rect 21560 1426 21588 1838
rect 21640 1828 21692 1834
rect 21640 1770 21692 1776
rect 21548 1420 21600 1426
rect 21548 1362 21600 1368
rect 20272 1278 20484 1294
rect 20076 1216 20128 1222
rect 20076 1158 20128 1164
rect 19984 876 20036 882
rect 19984 818 20036 824
rect 19248 808 19300 814
rect 19248 750 19300 756
rect 19800 808 19852 814
rect 19800 750 19852 756
rect 19524 740 19576 746
rect 19524 682 19576 688
rect 19536 400 19564 682
rect 19812 474 19840 750
rect 19800 468 19852 474
rect 19984 468 20036 474
rect 19800 410 19852 416
rect 19904 428 19984 456
rect 19904 400 19932 428
rect 19984 410 20036 416
rect 18972 196 19024 202
rect 18972 138 19024 144
rect 19154 0 19210 400
rect 19522 0 19578 400
rect 19890 0 19946 400
rect 20088 134 20116 1158
rect 20180 814 20208 1255
rect 20272 1018 20300 1278
rect 20682 1278 20944 1306
rect 20626 1255 20682 1264
rect 20352 1216 20404 1222
rect 20444 1216 20496 1222
rect 20352 1158 20404 1164
rect 20442 1184 20444 1193
rect 20536 1216 20588 1222
rect 20496 1184 20498 1193
rect 20260 1012 20312 1018
rect 20260 954 20312 960
rect 20364 814 20392 1158
rect 20536 1158 20588 1164
rect 20812 1216 20864 1222
rect 20812 1158 20864 1164
rect 20904 1216 20956 1222
rect 20904 1158 20956 1164
rect 20442 1119 20498 1128
rect 20444 944 20496 950
rect 20444 886 20496 892
rect 20168 808 20220 814
rect 20168 750 20220 756
rect 20352 808 20404 814
rect 20352 750 20404 756
rect 20076 128 20128 134
rect 20076 70 20128 76
rect 20180 66 20208 750
rect 20456 474 20484 886
rect 20548 882 20576 1158
rect 20718 1048 20774 1057
rect 20718 983 20774 992
rect 20536 876 20588 882
rect 20536 818 20588 824
rect 20732 814 20760 983
rect 20720 808 20772 814
rect 20720 750 20772 756
rect 20628 672 20680 678
rect 20548 632 20628 660
rect 20444 468 20496 474
rect 20272 428 20392 456
rect 20272 400 20300 428
rect 20168 60 20220 66
rect 20168 2 20220 8
rect 20258 0 20314 400
rect 20364 354 20392 428
rect 20444 410 20496 416
rect 20548 354 20576 632
rect 20628 614 20680 620
rect 20626 504 20682 513
rect 20626 439 20682 448
rect 20640 400 20668 439
rect 20364 326 20576 354
rect 20626 0 20682 400
rect 20824 270 20852 1158
rect 20916 338 20944 1158
rect 20996 944 21048 950
rect 21652 921 21680 1770
rect 21744 1494 21772 1838
rect 21824 1760 21876 1766
rect 21824 1702 21876 1708
rect 21732 1488 21784 1494
rect 21732 1430 21784 1436
rect 21836 1204 21864 1702
rect 21928 1358 21956 2246
rect 22112 2122 22140 2246
rect 22020 2094 22140 2122
rect 22192 2100 22244 2106
rect 22020 2038 22048 2094
rect 22192 2042 22244 2048
rect 22008 2032 22060 2038
rect 22008 1974 22060 1980
rect 22100 2032 22152 2038
rect 22100 1974 22152 1980
rect 21916 1352 21968 1358
rect 21916 1294 21968 1300
rect 21836 1176 21956 1204
rect 21824 1012 21876 1018
rect 21824 954 21876 960
rect 21732 944 21784 950
rect 20996 886 21048 892
rect 21638 912 21694 921
rect 21008 400 21036 886
rect 21732 886 21784 892
rect 21638 847 21694 856
rect 21548 672 21600 678
rect 21376 632 21548 660
rect 21376 400 21404 632
rect 21548 614 21600 620
rect 21744 400 21772 886
rect 21836 513 21864 954
rect 21928 814 21956 1176
rect 21916 808 21968 814
rect 21916 750 21968 756
rect 21822 504 21878 513
rect 21822 439 21878 448
rect 22112 400 22140 1974
rect 22204 1850 22232 2042
rect 22296 1952 22324 3334
rect 22756 2990 22784 3334
rect 22848 3058 22876 3878
rect 22836 3052 22888 3058
rect 22836 2994 22888 3000
rect 22744 2984 22796 2990
rect 22744 2926 22796 2932
rect 22836 2848 22888 2854
rect 22836 2790 22888 2796
rect 22364 2748 22740 2757
rect 22420 2746 22444 2748
rect 22500 2746 22524 2748
rect 22580 2746 22604 2748
rect 22660 2746 22684 2748
rect 22420 2694 22430 2746
rect 22674 2694 22684 2746
rect 22420 2692 22444 2694
rect 22500 2692 22524 2694
rect 22580 2692 22604 2694
rect 22660 2692 22684 2694
rect 22364 2683 22740 2692
rect 22376 2644 22428 2650
rect 22376 2586 22428 2592
rect 22388 2310 22416 2586
rect 22468 2508 22520 2514
rect 22468 2450 22520 2456
rect 22376 2304 22428 2310
rect 22480 2281 22508 2450
rect 22560 2304 22612 2310
rect 22376 2246 22428 2252
rect 22466 2272 22522 2281
rect 22388 2106 22416 2246
rect 22560 2246 22612 2252
rect 22466 2207 22522 2216
rect 22572 2106 22600 2246
rect 22376 2100 22428 2106
rect 22376 2042 22428 2048
rect 22560 2100 22612 2106
rect 22560 2042 22612 2048
rect 22376 1964 22428 1970
rect 22296 1924 22376 1952
rect 22376 1906 22428 1912
rect 22480 1958 22784 1986
rect 22480 1850 22508 1958
rect 22756 1902 22784 1958
rect 22560 1896 22612 1902
rect 22204 1822 22508 1850
rect 22558 1864 22560 1873
rect 22744 1896 22796 1902
rect 22612 1864 22614 1873
rect 22744 1838 22796 1844
rect 22558 1799 22614 1808
rect 22192 1760 22244 1766
rect 22192 1702 22244 1708
rect 22204 932 22232 1702
rect 22364 1660 22740 1669
rect 22420 1658 22444 1660
rect 22500 1658 22524 1660
rect 22580 1658 22604 1660
rect 22660 1658 22684 1660
rect 22420 1606 22430 1658
rect 22674 1606 22684 1658
rect 22420 1604 22444 1606
rect 22500 1604 22524 1606
rect 22580 1604 22604 1606
rect 22660 1604 22684 1606
rect 22364 1595 22740 1604
rect 22284 1556 22336 1562
rect 22284 1498 22336 1504
rect 22376 1556 22428 1562
rect 22376 1498 22428 1504
rect 22296 1306 22324 1498
rect 22388 1426 22416 1498
rect 22376 1420 22428 1426
rect 22376 1362 22428 1368
rect 22296 1278 22416 1306
rect 22204 904 22324 932
rect 22192 808 22244 814
rect 22192 750 22244 756
rect 22204 406 22232 750
rect 22296 456 22324 904
rect 22388 796 22416 1278
rect 22468 808 22520 814
rect 22388 768 22468 796
rect 22468 750 22520 756
rect 22364 572 22740 581
rect 22420 570 22444 572
rect 22500 570 22524 572
rect 22580 570 22604 572
rect 22660 570 22684 572
rect 22420 518 22430 570
rect 22674 518 22684 570
rect 22420 516 22444 518
rect 22500 516 22524 518
rect 22580 516 22604 518
rect 22660 516 22684 518
rect 22364 507 22740 516
rect 22296 428 22508 456
rect 22192 400 22244 406
rect 22480 400 22508 428
rect 22848 400 22876 2790
rect 22940 2514 22968 4150
rect 23112 4072 23164 4078
rect 23112 4014 23164 4020
rect 23020 3596 23072 3602
rect 23020 3538 23072 3544
rect 22928 2508 22980 2514
rect 22928 2450 22980 2456
rect 22928 1828 22980 1834
rect 22928 1770 22980 1776
rect 22940 1426 22968 1770
rect 23032 1766 23060 3538
rect 23124 2650 23152 4014
rect 23388 4004 23440 4010
rect 23388 3946 23440 3952
rect 23204 3528 23256 3534
rect 23204 3470 23256 3476
rect 23112 2644 23164 2650
rect 23112 2586 23164 2592
rect 23216 1986 23244 3470
rect 23296 2916 23348 2922
rect 23296 2858 23348 2864
rect 23124 1958 23244 1986
rect 23020 1760 23072 1766
rect 23020 1702 23072 1708
rect 23032 1494 23060 1702
rect 23020 1488 23072 1494
rect 23020 1430 23072 1436
rect 22928 1420 22980 1426
rect 22928 1362 22980 1368
rect 23124 814 23152 1958
rect 23204 1896 23256 1902
rect 23204 1838 23256 1844
rect 23112 808 23164 814
rect 23112 750 23164 756
rect 23216 400 23244 1838
rect 23308 1562 23336 2858
rect 23296 1556 23348 1562
rect 23296 1498 23348 1504
rect 23400 1358 23428 3946
rect 23572 3120 23624 3126
rect 23572 3062 23624 3068
rect 23388 1352 23440 1358
rect 23388 1294 23440 1300
rect 20904 332 20956 338
rect 20904 274 20956 280
rect 20812 264 20864 270
rect 20812 206 20864 212
rect 20994 0 21050 400
rect 21362 0 21418 400
rect 21730 0 21786 400
rect 22098 0 22154 400
rect 22192 342 22244 348
rect 22466 0 22522 400
rect 22834 0 22890 400
rect 23202 0 23258 400
rect 23400 202 23428 1294
rect 23584 400 23612 3062
rect 23388 196 23440 202
rect 23388 138 23440 144
rect 23570 0 23626 400
<< via2 >>
rect 1364 22874 1420 22876
rect 1444 22874 1500 22876
rect 1524 22874 1580 22876
rect 1604 22874 1660 22876
rect 1684 22874 1740 22876
rect 1364 22822 1366 22874
rect 1366 22822 1418 22874
rect 1418 22822 1420 22874
rect 1444 22822 1482 22874
rect 1482 22822 1494 22874
rect 1494 22822 1500 22874
rect 1524 22822 1546 22874
rect 1546 22822 1558 22874
rect 1558 22822 1580 22874
rect 1604 22822 1610 22874
rect 1610 22822 1622 22874
rect 1622 22822 1660 22874
rect 1684 22822 1686 22874
rect 1686 22822 1738 22874
rect 1738 22822 1740 22874
rect 1364 22820 1420 22822
rect 1444 22820 1500 22822
rect 1524 22820 1580 22822
rect 1604 22820 1660 22822
rect 1684 22820 1740 22822
rect 1364 21786 1420 21788
rect 1444 21786 1500 21788
rect 1524 21786 1580 21788
rect 1604 21786 1660 21788
rect 1684 21786 1740 21788
rect 1364 21734 1366 21786
rect 1366 21734 1418 21786
rect 1418 21734 1420 21786
rect 1444 21734 1482 21786
rect 1482 21734 1494 21786
rect 1494 21734 1500 21786
rect 1524 21734 1546 21786
rect 1546 21734 1558 21786
rect 1558 21734 1580 21786
rect 1604 21734 1610 21786
rect 1610 21734 1622 21786
rect 1622 21734 1660 21786
rect 1684 21734 1686 21786
rect 1686 21734 1738 21786
rect 1738 21734 1740 21786
rect 1364 21732 1420 21734
rect 1444 21732 1500 21734
rect 1524 21732 1580 21734
rect 1604 21732 1660 21734
rect 1684 21732 1740 21734
rect 1364 20698 1420 20700
rect 1444 20698 1500 20700
rect 1524 20698 1580 20700
rect 1604 20698 1660 20700
rect 1684 20698 1740 20700
rect 1364 20646 1366 20698
rect 1366 20646 1418 20698
rect 1418 20646 1420 20698
rect 1444 20646 1482 20698
rect 1482 20646 1494 20698
rect 1494 20646 1500 20698
rect 1524 20646 1546 20698
rect 1546 20646 1558 20698
rect 1558 20646 1580 20698
rect 1604 20646 1610 20698
rect 1610 20646 1622 20698
rect 1622 20646 1660 20698
rect 1684 20646 1686 20698
rect 1686 20646 1738 20698
rect 1738 20646 1740 20698
rect 1364 20644 1420 20646
rect 1444 20644 1500 20646
rect 1524 20644 1580 20646
rect 1604 20644 1660 20646
rect 1684 20644 1740 20646
rect 2962 22344 3018 22400
rect 2778 21392 2834 21448
rect 4364 23418 4420 23420
rect 4444 23418 4500 23420
rect 4524 23418 4580 23420
rect 4604 23418 4660 23420
rect 4684 23418 4740 23420
rect 4364 23366 4366 23418
rect 4366 23366 4418 23418
rect 4418 23366 4420 23418
rect 4444 23366 4482 23418
rect 4482 23366 4494 23418
rect 4494 23366 4500 23418
rect 4524 23366 4546 23418
rect 4546 23366 4558 23418
rect 4558 23366 4580 23418
rect 4604 23366 4610 23418
rect 4610 23366 4622 23418
rect 4622 23366 4660 23418
rect 4684 23366 4686 23418
rect 4686 23366 4738 23418
rect 4738 23366 4740 23418
rect 4364 23364 4420 23366
rect 4444 23364 4500 23366
rect 4524 23364 4580 23366
rect 4604 23364 4660 23366
rect 4684 23364 4740 23366
rect 2134 20440 2190 20496
rect 2042 20340 2044 20360
rect 2044 20340 2096 20360
rect 2096 20340 2098 20360
rect 2042 20304 2098 20340
rect 1364 19610 1420 19612
rect 1444 19610 1500 19612
rect 1524 19610 1580 19612
rect 1604 19610 1660 19612
rect 1684 19610 1740 19612
rect 1364 19558 1366 19610
rect 1366 19558 1418 19610
rect 1418 19558 1420 19610
rect 1444 19558 1482 19610
rect 1482 19558 1494 19610
rect 1494 19558 1500 19610
rect 1524 19558 1546 19610
rect 1546 19558 1558 19610
rect 1558 19558 1580 19610
rect 1604 19558 1610 19610
rect 1610 19558 1622 19610
rect 1622 19558 1660 19610
rect 1684 19558 1686 19610
rect 1686 19558 1738 19610
rect 1738 19558 1740 19610
rect 1364 19556 1420 19558
rect 1444 19556 1500 19558
rect 1524 19556 1580 19558
rect 1604 19556 1660 19558
rect 1684 19556 1740 19558
rect 1950 19216 2006 19272
rect 1364 18522 1420 18524
rect 1444 18522 1500 18524
rect 1524 18522 1580 18524
rect 1604 18522 1660 18524
rect 1684 18522 1740 18524
rect 1364 18470 1366 18522
rect 1366 18470 1418 18522
rect 1418 18470 1420 18522
rect 1444 18470 1482 18522
rect 1482 18470 1494 18522
rect 1494 18470 1500 18522
rect 1524 18470 1546 18522
rect 1546 18470 1558 18522
rect 1558 18470 1580 18522
rect 1604 18470 1610 18522
rect 1610 18470 1622 18522
rect 1622 18470 1660 18522
rect 1684 18470 1686 18522
rect 1686 18470 1738 18522
rect 1738 18470 1740 18522
rect 1364 18468 1420 18470
rect 1444 18468 1500 18470
rect 1524 18468 1580 18470
rect 1604 18468 1660 18470
rect 1684 18468 1740 18470
rect 4364 22330 4420 22332
rect 4444 22330 4500 22332
rect 4524 22330 4580 22332
rect 4604 22330 4660 22332
rect 4684 22330 4740 22332
rect 4364 22278 4366 22330
rect 4366 22278 4418 22330
rect 4418 22278 4420 22330
rect 4444 22278 4482 22330
rect 4482 22278 4494 22330
rect 4494 22278 4500 22330
rect 4524 22278 4546 22330
rect 4546 22278 4558 22330
rect 4558 22278 4580 22330
rect 4604 22278 4610 22330
rect 4610 22278 4622 22330
rect 4622 22278 4660 22330
rect 4684 22278 4686 22330
rect 4686 22278 4738 22330
rect 4738 22278 4740 22330
rect 4364 22276 4420 22278
rect 4444 22276 4500 22278
rect 4524 22276 4580 22278
rect 4604 22276 4660 22278
rect 4684 22276 4740 22278
rect 5354 22072 5410 22128
rect 3882 21528 3938 21584
rect 3514 21004 3570 21040
rect 3514 20984 3516 21004
rect 3516 20984 3568 21004
rect 3568 20984 3570 21004
rect 4066 20848 4122 20904
rect 4364 21242 4420 21244
rect 4444 21242 4500 21244
rect 4524 21242 4580 21244
rect 4604 21242 4660 21244
rect 4684 21242 4740 21244
rect 4364 21190 4366 21242
rect 4366 21190 4418 21242
rect 4418 21190 4420 21242
rect 4444 21190 4482 21242
rect 4482 21190 4494 21242
rect 4494 21190 4500 21242
rect 4524 21190 4546 21242
rect 4546 21190 4558 21242
rect 4558 21190 4580 21242
rect 4604 21190 4610 21242
rect 4610 21190 4622 21242
rect 4622 21190 4660 21242
rect 4684 21190 4686 21242
rect 4686 21190 4738 21242
rect 4738 21190 4740 21242
rect 4364 21188 4420 21190
rect 4444 21188 4500 21190
rect 4524 21188 4580 21190
rect 4604 21188 4660 21190
rect 4684 21188 4740 21190
rect 4986 21120 5042 21176
rect 2226 19080 2282 19136
rect 4710 20848 4766 20904
rect 4364 20154 4420 20156
rect 4444 20154 4500 20156
rect 4524 20154 4580 20156
rect 4604 20154 4660 20156
rect 4684 20154 4740 20156
rect 4364 20102 4366 20154
rect 4366 20102 4418 20154
rect 4418 20102 4420 20154
rect 4444 20102 4482 20154
rect 4482 20102 4494 20154
rect 4494 20102 4500 20154
rect 4524 20102 4546 20154
rect 4546 20102 4558 20154
rect 4558 20102 4580 20154
rect 4604 20102 4610 20154
rect 4610 20102 4622 20154
rect 4622 20102 4660 20154
rect 4684 20102 4686 20154
rect 4686 20102 4738 20154
rect 4738 20102 4740 20154
rect 4364 20100 4420 20102
rect 4444 20100 4500 20102
rect 4524 20100 4580 20102
rect 4604 20100 4660 20102
rect 4684 20100 4740 20102
rect 3422 19352 3478 19408
rect 4066 19252 4068 19272
rect 4068 19252 4120 19272
rect 4120 19252 4122 19272
rect 3790 19080 3846 19136
rect 4066 19216 4122 19252
rect 4364 19066 4420 19068
rect 4444 19066 4500 19068
rect 4524 19066 4580 19068
rect 4604 19066 4660 19068
rect 4684 19066 4740 19068
rect 4364 19014 4366 19066
rect 4366 19014 4418 19066
rect 4418 19014 4420 19066
rect 4444 19014 4482 19066
rect 4482 19014 4494 19066
rect 4494 19014 4500 19066
rect 4524 19014 4546 19066
rect 4546 19014 4558 19066
rect 4558 19014 4580 19066
rect 4604 19014 4610 19066
rect 4610 19014 4622 19066
rect 4622 19014 4660 19066
rect 4684 19014 4686 19066
rect 4686 19014 4738 19066
rect 4738 19014 4740 19066
rect 4364 19012 4420 19014
rect 4444 19012 4500 19014
rect 4524 19012 4580 19014
rect 4604 19012 4660 19014
rect 4684 19012 4740 19014
rect 5446 19916 5502 19952
rect 5446 19896 5448 19916
rect 5448 19896 5500 19916
rect 5500 19896 5502 19916
rect 6090 21004 6146 21040
rect 6090 20984 6092 21004
rect 6092 20984 6144 21004
rect 6144 20984 6146 21004
rect 6274 20848 6330 20904
rect 7364 22874 7420 22876
rect 7444 22874 7500 22876
rect 7524 22874 7580 22876
rect 7604 22874 7660 22876
rect 7684 22874 7740 22876
rect 7364 22822 7366 22874
rect 7366 22822 7418 22874
rect 7418 22822 7420 22874
rect 7444 22822 7482 22874
rect 7482 22822 7494 22874
rect 7494 22822 7500 22874
rect 7524 22822 7546 22874
rect 7546 22822 7558 22874
rect 7558 22822 7580 22874
rect 7604 22822 7610 22874
rect 7610 22822 7622 22874
rect 7622 22822 7660 22874
rect 7684 22822 7686 22874
rect 7686 22822 7738 22874
rect 7738 22822 7740 22874
rect 7364 22820 7420 22822
rect 7444 22820 7500 22822
rect 7524 22820 7580 22822
rect 7604 22820 7660 22822
rect 7684 22820 7740 22822
rect 1364 17434 1420 17436
rect 1444 17434 1500 17436
rect 1524 17434 1580 17436
rect 1604 17434 1660 17436
rect 1684 17434 1740 17436
rect 1364 17382 1366 17434
rect 1366 17382 1418 17434
rect 1418 17382 1420 17434
rect 1444 17382 1482 17434
rect 1482 17382 1494 17434
rect 1494 17382 1500 17434
rect 1524 17382 1546 17434
rect 1546 17382 1558 17434
rect 1558 17382 1580 17434
rect 1604 17382 1610 17434
rect 1610 17382 1622 17434
rect 1622 17382 1660 17434
rect 1684 17382 1686 17434
rect 1686 17382 1738 17434
rect 1738 17382 1740 17434
rect 1364 17380 1420 17382
rect 1444 17380 1500 17382
rect 1524 17380 1580 17382
rect 1604 17380 1660 17382
rect 1684 17380 1740 17382
rect 1364 16346 1420 16348
rect 1444 16346 1500 16348
rect 1524 16346 1580 16348
rect 1604 16346 1660 16348
rect 1684 16346 1740 16348
rect 1364 16294 1366 16346
rect 1366 16294 1418 16346
rect 1418 16294 1420 16346
rect 1444 16294 1482 16346
rect 1482 16294 1494 16346
rect 1494 16294 1500 16346
rect 1524 16294 1546 16346
rect 1546 16294 1558 16346
rect 1558 16294 1580 16346
rect 1604 16294 1610 16346
rect 1610 16294 1622 16346
rect 1622 16294 1660 16346
rect 1684 16294 1686 16346
rect 1686 16294 1738 16346
rect 1738 16294 1740 16346
rect 1364 16292 1420 16294
rect 1444 16292 1500 16294
rect 1524 16292 1580 16294
rect 1604 16292 1660 16294
rect 1684 16292 1740 16294
rect 1214 15952 1270 16008
rect 2410 16652 2466 16688
rect 2410 16632 2412 16652
rect 2412 16632 2464 16652
rect 2464 16632 2466 16652
rect 2502 16496 2558 16552
rect 1364 15258 1420 15260
rect 1444 15258 1500 15260
rect 1524 15258 1580 15260
rect 1604 15258 1660 15260
rect 1684 15258 1740 15260
rect 1364 15206 1366 15258
rect 1366 15206 1418 15258
rect 1418 15206 1420 15258
rect 1444 15206 1482 15258
rect 1482 15206 1494 15258
rect 1494 15206 1500 15258
rect 1524 15206 1546 15258
rect 1546 15206 1558 15258
rect 1558 15206 1580 15258
rect 1604 15206 1610 15258
rect 1610 15206 1622 15258
rect 1622 15206 1660 15258
rect 1684 15206 1686 15258
rect 1686 15206 1738 15258
rect 1738 15206 1740 15258
rect 1364 15204 1420 15206
rect 1444 15204 1500 15206
rect 1524 15204 1580 15206
rect 1604 15204 1660 15206
rect 1684 15204 1740 15206
rect 1364 14170 1420 14172
rect 1444 14170 1500 14172
rect 1524 14170 1580 14172
rect 1604 14170 1660 14172
rect 1684 14170 1740 14172
rect 1364 14118 1366 14170
rect 1366 14118 1418 14170
rect 1418 14118 1420 14170
rect 1444 14118 1482 14170
rect 1482 14118 1494 14170
rect 1494 14118 1500 14170
rect 1524 14118 1546 14170
rect 1546 14118 1558 14170
rect 1558 14118 1580 14170
rect 1604 14118 1610 14170
rect 1610 14118 1622 14170
rect 1622 14118 1660 14170
rect 1684 14118 1686 14170
rect 1686 14118 1738 14170
rect 1738 14118 1740 14170
rect 1364 14116 1420 14118
rect 1444 14116 1500 14118
rect 1524 14116 1580 14118
rect 1604 14116 1660 14118
rect 1684 14116 1740 14118
rect 2686 17620 2688 17640
rect 2688 17620 2740 17640
rect 2740 17620 2742 17640
rect 2686 17584 2742 17620
rect 3054 17040 3110 17096
rect 3790 17176 3846 17232
rect 5078 18264 5134 18320
rect 4066 18164 4068 18184
rect 4068 18164 4120 18184
rect 4120 18164 4122 18184
rect 4066 18128 4122 18164
rect 2594 16088 2650 16144
rect 3790 16652 3846 16688
rect 3790 16632 3792 16652
rect 3792 16632 3844 16652
rect 3844 16632 3846 16652
rect 2962 16496 3018 16552
rect 3514 16496 3570 16552
rect 2870 15408 2926 15464
rect 3330 15444 3332 15464
rect 3332 15444 3384 15464
rect 3384 15444 3386 15464
rect 3330 15408 3386 15444
rect 1364 13082 1420 13084
rect 1444 13082 1500 13084
rect 1524 13082 1580 13084
rect 1604 13082 1660 13084
rect 1684 13082 1740 13084
rect 1364 13030 1366 13082
rect 1366 13030 1418 13082
rect 1418 13030 1420 13082
rect 1444 13030 1482 13082
rect 1482 13030 1494 13082
rect 1494 13030 1500 13082
rect 1524 13030 1546 13082
rect 1546 13030 1558 13082
rect 1558 13030 1580 13082
rect 1604 13030 1610 13082
rect 1610 13030 1622 13082
rect 1622 13030 1660 13082
rect 1684 13030 1686 13082
rect 1686 13030 1738 13082
rect 1738 13030 1740 13082
rect 1364 13028 1420 13030
rect 1444 13028 1500 13030
rect 1524 13028 1580 13030
rect 1604 13028 1660 13030
rect 1684 13028 1740 13030
rect 1490 12144 1546 12200
rect 1364 11994 1420 11996
rect 1444 11994 1500 11996
rect 1524 11994 1580 11996
rect 1604 11994 1660 11996
rect 1684 11994 1740 11996
rect 1364 11942 1366 11994
rect 1366 11942 1418 11994
rect 1418 11942 1420 11994
rect 1444 11942 1482 11994
rect 1482 11942 1494 11994
rect 1494 11942 1500 11994
rect 1524 11942 1546 11994
rect 1546 11942 1558 11994
rect 1558 11942 1580 11994
rect 1604 11942 1610 11994
rect 1610 11942 1622 11994
rect 1622 11942 1660 11994
rect 1684 11942 1686 11994
rect 1686 11942 1738 11994
rect 1738 11942 1740 11994
rect 1364 11940 1420 11942
rect 1444 11940 1500 11942
rect 1524 11940 1580 11942
rect 1604 11940 1660 11942
rect 1684 11940 1740 11942
rect 1364 10906 1420 10908
rect 1444 10906 1500 10908
rect 1524 10906 1580 10908
rect 1604 10906 1660 10908
rect 1684 10906 1740 10908
rect 1364 10854 1366 10906
rect 1366 10854 1418 10906
rect 1418 10854 1420 10906
rect 1444 10854 1482 10906
rect 1482 10854 1494 10906
rect 1494 10854 1500 10906
rect 1524 10854 1546 10906
rect 1546 10854 1558 10906
rect 1558 10854 1580 10906
rect 1604 10854 1610 10906
rect 1610 10854 1622 10906
rect 1622 10854 1660 10906
rect 1684 10854 1686 10906
rect 1686 10854 1738 10906
rect 1738 10854 1740 10906
rect 1364 10852 1420 10854
rect 1444 10852 1500 10854
rect 1524 10852 1580 10854
rect 1604 10852 1660 10854
rect 1684 10852 1740 10854
rect 1364 9818 1420 9820
rect 1444 9818 1500 9820
rect 1524 9818 1580 9820
rect 1604 9818 1660 9820
rect 1684 9818 1740 9820
rect 1364 9766 1366 9818
rect 1366 9766 1418 9818
rect 1418 9766 1420 9818
rect 1444 9766 1482 9818
rect 1482 9766 1494 9818
rect 1494 9766 1500 9818
rect 1524 9766 1546 9818
rect 1546 9766 1558 9818
rect 1558 9766 1580 9818
rect 1604 9766 1610 9818
rect 1610 9766 1622 9818
rect 1622 9766 1660 9818
rect 1684 9766 1686 9818
rect 1686 9766 1738 9818
rect 1738 9766 1740 9818
rect 1364 9764 1420 9766
rect 1444 9764 1500 9766
rect 1524 9764 1580 9766
rect 1604 9764 1660 9766
rect 1684 9764 1740 9766
rect 1398 9460 1400 9480
rect 1400 9460 1452 9480
rect 1452 9460 1454 9480
rect 1398 9424 1454 9460
rect 1582 9172 1638 9208
rect 1582 9152 1584 9172
rect 1584 9152 1636 9172
rect 1636 9152 1638 9172
rect 1950 12144 2006 12200
rect 2318 12860 2320 12880
rect 2320 12860 2372 12880
rect 2372 12860 2374 12880
rect 2318 12824 2374 12860
rect 1950 9152 2006 9208
rect 1364 8730 1420 8732
rect 1444 8730 1500 8732
rect 1524 8730 1580 8732
rect 1604 8730 1660 8732
rect 1684 8730 1740 8732
rect 1364 8678 1366 8730
rect 1366 8678 1418 8730
rect 1418 8678 1420 8730
rect 1444 8678 1482 8730
rect 1482 8678 1494 8730
rect 1494 8678 1500 8730
rect 1524 8678 1546 8730
rect 1546 8678 1558 8730
rect 1558 8678 1580 8730
rect 1604 8678 1610 8730
rect 1610 8678 1622 8730
rect 1622 8678 1660 8730
rect 1684 8678 1686 8730
rect 1686 8678 1738 8730
rect 1738 8678 1740 8730
rect 1364 8676 1420 8678
rect 1444 8676 1500 8678
rect 1524 8676 1580 8678
rect 1604 8676 1660 8678
rect 1684 8676 1740 8678
rect 1364 7642 1420 7644
rect 1444 7642 1500 7644
rect 1524 7642 1580 7644
rect 1604 7642 1660 7644
rect 1684 7642 1740 7644
rect 1364 7590 1366 7642
rect 1366 7590 1418 7642
rect 1418 7590 1420 7642
rect 1444 7590 1482 7642
rect 1482 7590 1494 7642
rect 1494 7590 1500 7642
rect 1524 7590 1546 7642
rect 1546 7590 1558 7642
rect 1558 7590 1580 7642
rect 1604 7590 1610 7642
rect 1610 7590 1622 7642
rect 1622 7590 1660 7642
rect 1684 7590 1686 7642
rect 1686 7590 1738 7642
rect 1738 7590 1740 7642
rect 1364 7588 1420 7590
rect 1444 7588 1500 7590
rect 1524 7588 1580 7590
rect 1604 7588 1660 7590
rect 1684 7588 1740 7590
rect 2318 8608 2374 8664
rect 1364 6554 1420 6556
rect 1444 6554 1500 6556
rect 1524 6554 1580 6556
rect 1604 6554 1660 6556
rect 1684 6554 1740 6556
rect 1364 6502 1366 6554
rect 1366 6502 1418 6554
rect 1418 6502 1420 6554
rect 1444 6502 1482 6554
rect 1482 6502 1494 6554
rect 1494 6502 1500 6554
rect 1524 6502 1546 6554
rect 1546 6502 1558 6554
rect 1558 6502 1580 6554
rect 1604 6502 1610 6554
rect 1610 6502 1622 6554
rect 1622 6502 1660 6554
rect 1684 6502 1686 6554
rect 1686 6502 1738 6554
rect 1738 6502 1740 6554
rect 1364 6500 1420 6502
rect 1444 6500 1500 6502
rect 1524 6500 1580 6502
rect 1604 6500 1660 6502
rect 1684 6500 1740 6502
rect 1364 5466 1420 5468
rect 1444 5466 1500 5468
rect 1524 5466 1580 5468
rect 1604 5466 1660 5468
rect 1684 5466 1740 5468
rect 1364 5414 1366 5466
rect 1366 5414 1418 5466
rect 1418 5414 1420 5466
rect 1444 5414 1482 5466
rect 1482 5414 1494 5466
rect 1494 5414 1500 5466
rect 1524 5414 1546 5466
rect 1546 5414 1558 5466
rect 1558 5414 1580 5466
rect 1604 5414 1610 5466
rect 1610 5414 1622 5466
rect 1622 5414 1660 5466
rect 1684 5414 1686 5466
rect 1686 5414 1738 5466
rect 1738 5414 1740 5466
rect 1364 5412 1420 5414
rect 1444 5412 1500 5414
rect 1524 5412 1580 5414
rect 1604 5412 1660 5414
rect 1684 5412 1740 5414
rect 1364 4378 1420 4380
rect 1444 4378 1500 4380
rect 1524 4378 1580 4380
rect 1604 4378 1660 4380
rect 1684 4378 1740 4380
rect 1364 4326 1366 4378
rect 1366 4326 1418 4378
rect 1418 4326 1420 4378
rect 1444 4326 1482 4378
rect 1482 4326 1494 4378
rect 1494 4326 1500 4378
rect 1524 4326 1546 4378
rect 1546 4326 1558 4378
rect 1558 4326 1580 4378
rect 1604 4326 1610 4378
rect 1610 4326 1622 4378
rect 1622 4326 1660 4378
rect 1684 4326 1686 4378
rect 1686 4326 1738 4378
rect 1738 4326 1740 4378
rect 1364 4324 1420 4326
rect 1444 4324 1500 4326
rect 1524 4324 1580 4326
rect 1604 4324 1660 4326
rect 1684 4324 1740 4326
rect 1364 3290 1420 3292
rect 1444 3290 1500 3292
rect 1524 3290 1580 3292
rect 1604 3290 1660 3292
rect 1684 3290 1740 3292
rect 1364 3238 1366 3290
rect 1366 3238 1418 3290
rect 1418 3238 1420 3290
rect 1444 3238 1482 3290
rect 1482 3238 1494 3290
rect 1494 3238 1500 3290
rect 1524 3238 1546 3290
rect 1546 3238 1558 3290
rect 1558 3238 1580 3290
rect 1604 3238 1610 3290
rect 1610 3238 1622 3290
rect 1622 3238 1660 3290
rect 1684 3238 1686 3290
rect 1686 3238 1738 3290
rect 1738 3238 1740 3290
rect 1364 3236 1420 3238
rect 1444 3236 1500 3238
rect 1524 3236 1580 3238
rect 1604 3236 1660 3238
rect 1684 3236 1740 3238
rect 1364 2202 1420 2204
rect 1444 2202 1500 2204
rect 1524 2202 1580 2204
rect 1604 2202 1660 2204
rect 1684 2202 1740 2204
rect 1364 2150 1366 2202
rect 1366 2150 1418 2202
rect 1418 2150 1420 2202
rect 1444 2150 1482 2202
rect 1482 2150 1494 2202
rect 1494 2150 1500 2202
rect 1524 2150 1546 2202
rect 1546 2150 1558 2202
rect 1558 2150 1580 2202
rect 1604 2150 1610 2202
rect 1610 2150 1622 2202
rect 1622 2150 1660 2202
rect 1684 2150 1686 2202
rect 1686 2150 1738 2202
rect 1738 2150 1740 2202
rect 1364 2148 1420 2150
rect 1444 2148 1500 2150
rect 1524 2148 1580 2150
rect 1604 2148 1660 2150
rect 1684 2148 1740 2150
rect 3146 8372 3148 8392
rect 3148 8372 3200 8392
rect 3200 8372 3202 8392
rect 3146 8336 3202 8372
rect 3146 7948 3202 7984
rect 3146 7928 3148 7948
rect 3148 7928 3200 7948
rect 3200 7928 3202 7948
rect 3330 9424 3386 9480
rect 3882 14476 3938 14512
rect 3882 14456 3884 14476
rect 3884 14456 3936 14476
rect 3936 14456 3938 14476
rect 4364 17978 4420 17980
rect 4444 17978 4500 17980
rect 4524 17978 4580 17980
rect 4604 17978 4660 17980
rect 4684 17978 4740 17980
rect 4364 17926 4366 17978
rect 4366 17926 4418 17978
rect 4418 17926 4420 17978
rect 4444 17926 4482 17978
rect 4482 17926 4494 17978
rect 4494 17926 4500 17978
rect 4524 17926 4546 17978
rect 4546 17926 4558 17978
rect 4558 17926 4580 17978
rect 4604 17926 4610 17978
rect 4610 17926 4622 17978
rect 4622 17926 4660 17978
rect 4684 17926 4686 17978
rect 4686 17926 4738 17978
rect 4738 17926 4740 17978
rect 4364 17924 4420 17926
rect 4444 17924 4500 17926
rect 4524 17924 4580 17926
rect 4604 17924 4660 17926
rect 4684 17924 4740 17926
rect 4364 16890 4420 16892
rect 4444 16890 4500 16892
rect 4524 16890 4580 16892
rect 4604 16890 4660 16892
rect 4684 16890 4740 16892
rect 4364 16838 4366 16890
rect 4366 16838 4418 16890
rect 4418 16838 4420 16890
rect 4444 16838 4482 16890
rect 4482 16838 4494 16890
rect 4494 16838 4500 16890
rect 4524 16838 4546 16890
rect 4546 16838 4558 16890
rect 4558 16838 4580 16890
rect 4604 16838 4610 16890
rect 4610 16838 4622 16890
rect 4622 16838 4660 16890
rect 4684 16838 4686 16890
rect 4686 16838 4738 16890
rect 4738 16838 4740 16890
rect 4364 16836 4420 16838
rect 4444 16836 4500 16838
rect 4524 16836 4580 16838
rect 4604 16836 4660 16838
rect 4684 16836 4740 16838
rect 4802 16516 4858 16552
rect 4802 16496 4804 16516
rect 4804 16496 4856 16516
rect 4856 16496 4858 16516
rect 5078 17176 5134 17232
rect 5262 17040 5318 17096
rect 4364 15802 4420 15804
rect 4444 15802 4500 15804
rect 4524 15802 4580 15804
rect 4604 15802 4660 15804
rect 4684 15802 4740 15804
rect 4364 15750 4366 15802
rect 4366 15750 4418 15802
rect 4418 15750 4420 15802
rect 4444 15750 4482 15802
rect 4482 15750 4494 15802
rect 4494 15750 4500 15802
rect 4524 15750 4546 15802
rect 4546 15750 4558 15802
rect 4558 15750 4580 15802
rect 4604 15750 4610 15802
rect 4610 15750 4622 15802
rect 4622 15750 4660 15802
rect 4684 15750 4686 15802
rect 4686 15750 4738 15802
rect 4738 15750 4740 15802
rect 4364 15748 4420 15750
rect 4444 15748 4500 15750
rect 4524 15748 4580 15750
rect 4604 15748 4660 15750
rect 4684 15748 4740 15750
rect 4250 15136 4306 15192
rect 4434 15000 4490 15056
rect 4986 15408 5042 15464
rect 4710 14884 4766 14920
rect 4710 14864 4712 14884
rect 4712 14864 4764 14884
rect 4764 14864 4766 14884
rect 4364 14714 4420 14716
rect 4444 14714 4500 14716
rect 4524 14714 4580 14716
rect 4604 14714 4660 14716
rect 4684 14714 4740 14716
rect 4364 14662 4366 14714
rect 4366 14662 4418 14714
rect 4418 14662 4420 14714
rect 4444 14662 4482 14714
rect 4482 14662 4494 14714
rect 4494 14662 4500 14714
rect 4524 14662 4546 14714
rect 4546 14662 4558 14714
rect 4558 14662 4580 14714
rect 4604 14662 4610 14714
rect 4610 14662 4622 14714
rect 4622 14662 4660 14714
rect 4684 14662 4686 14714
rect 4686 14662 4738 14714
rect 4738 14662 4740 14714
rect 4364 14660 4420 14662
rect 4444 14660 4500 14662
rect 4524 14660 4580 14662
rect 4604 14660 4660 14662
rect 4684 14660 4740 14662
rect 4618 14320 4674 14376
rect 3606 9460 3608 9480
rect 3608 9460 3660 9480
rect 3660 9460 3662 9480
rect 3606 9424 3662 9460
rect 3790 8336 3846 8392
rect 4364 13626 4420 13628
rect 4444 13626 4500 13628
rect 4524 13626 4580 13628
rect 4604 13626 4660 13628
rect 4684 13626 4740 13628
rect 4364 13574 4366 13626
rect 4366 13574 4418 13626
rect 4418 13574 4420 13626
rect 4444 13574 4482 13626
rect 4482 13574 4494 13626
rect 4494 13574 4500 13626
rect 4524 13574 4546 13626
rect 4546 13574 4558 13626
rect 4558 13574 4580 13626
rect 4604 13574 4610 13626
rect 4610 13574 4622 13626
rect 4622 13574 4660 13626
rect 4684 13574 4686 13626
rect 4686 13574 4738 13626
rect 4738 13574 4740 13626
rect 4364 13572 4420 13574
rect 4444 13572 4500 13574
rect 4524 13572 4580 13574
rect 4604 13572 4660 13574
rect 4684 13572 4740 13574
rect 4250 13388 4306 13424
rect 4250 13368 4252 13388
rect 4252 13368 4304 13388
rect 4304 13368 4306 13388
rect 6550 20712 6606 20768
rect 6550 20032 6606 20088
rect 5722 18572 5724 18592
rect 5724 18572 5776 18592
rect 5776 18572 5778 18592
rect 5722 18536 5778 18572
rect 5354 15816 5410 15872
rect 5814 17584 5870 17640
rect 5814 17076 5816 17096
rect 5816 17076 5868 17096
rect 5868 17076 5870 17096
rect 5814 17040 5870 17076
rect 7102 21256 7158 21312
rect 6918 20168 6974 20224
rect 6918 19236 6974 19272
rect 6918 19216 6920 19236
rect 6920 19216 6972 19236
rect 6972 19216 6974 19236
rect 6826 19080 6882 19136
rect 7364 21786 7420 21788
rect 7444 21786 7500 21788
rect 7524 21786 7580 21788
rect 7604 21786 7660 21788
rect 7684 21786 7740 21788
rect 7364 21734 7366 21786
rect 7366 21734 7418 21786
rect 7418 21734 7420 21786
rect 7444 21734 7482 21786
rect 7482 21734 7494 21786
rect 7494 21734 7500 21786
rect 7524 21734 7546 21786
rect 7546 21734 7558 21786
rect 7558 21734 7580 21786
rect 7604 21734 7610 21786
rect 7610 21734 7622 21786
rect 7622 21734 7660 21786
rect 7684 21734 7686 21786
rect 7686 21734 7738 21786
rect 7738 21734 7740 21786
rect 7364 21732 7420 21734
rect 7444 21732 7500 21734
rect 7524 21732 7580 21734
rect 7604 21732 7660 21734
rect 7684 21732 7740 21734
rect 7378 20984 7434 21040
rect 8022 21956 8078 21992
rect 8022 21936 8024 21956
rect 8024 21936 8076 21956
rect 8076 21936 8078 21956
rect 8574 21528 8630 21584
rect 7364 20698 7420 20700
rect 7444 20698 7500 20700
rect 7524 20698 7580 20700
rect 7604 20698 7660 20700
rect 7684 20698 7740 20700
rect 7364 20646 7366 20698
rect 7366 20646 7418 20698
rect 7418 20646 7420 20698
rect 7444 20646 7482 20698
rect 7482 20646 7494 20698
rect 7494 20646 7500 20698
rect 7524 20646 7546 20698
rect 7546 20646 7558 20698
rect 7558 20646 7580 20698
rect 7604 20646 7610 20698
rect 7610 20646 7622 20698
rect 7622 20646 7660 20698
rect 7684 20646 7686 20698
rect 7686 20646 7738 20698
rect 7738 20646 7740 20698
rect 7364 20644 7420 20646
rect 7444 20644 7500 20646
rect 7524 20644 7580 20646
rect 7604 20644 7660 20646
rect 7684 20644 7740 20646
rect 7378 19760 7434 19816
rect 8022 19896 8078 19952
rect 7930 19760 7986 19816
rect 8206 20032 8262 20088
rect 7364 19610 7420 19612
rect 7444 19610 7500 19612
rect 7524 19610 7580 19612
rect 7604 19610 7660 19612
rect 7684 19610 7740 19612
rect 7364 19558 7366 19610
rect 7366 19558 7418 19610
rect 7418 19558 7420 19610
rect 7444 19558 7482 19610
rect 7482 19558 7494 19610
rect 7494 19558 7500 19610
rect 7524 19558 7546 19610
rect 7546 19558 7558 19610
rect 7558 19558 7580 19610
rect 7604 19558 7610 19610
rect 7610 19558 7622 19610
rect 7622 19558 7660 19610
rect 7684 19558 7686 19610
rect 7686 19558 7738 19610
rect 7738 19558 7740 19610
rect 7364 19556 7420 19558
rect 7444 19556 7500 19558
rect 7524 19556 7580 19558
rect 7604 19556 7660 19558
rect 7684 19556 7740 19558
rect 7010 18536 7066 18592
rect 7364 18522 7420 18524
rect 7444 18522 7500 18524
rect 7524 18522 7580 18524
rect 7604 18522 7660 18524
rect 7684 18522 7740 18524
rect 7364 18470 7366 18522
rect 7366 18470 7418 18522
rect 7418 18470 7420 18522
rect 7444 18470 7482 18522
rect 7482 18470 7494 18522
rect 7494 18470 7500 18522
rect 7524 18470 7546 18522
rect 7546 18470 7558 18522
rect 7558 18470 7580 18522
rect 7604 18470 7610 18522
rect 7610 18470 7622 18522
rect 7622 18470 7660 18522
rect 7684 18470 7686 18522
rect 7686 18470 7738 18522
rect 7738 18470 7740 18522
rect 7364 18468 7420 18470
rect 7444 18468 7500 18470
rect 7524 18468 7580 18470
rect 7604 18468 7660 18470
rect 7684 18468 7740 18470
rect 8758 21256 8814 21312
rect 8942 21120 8998 21176
rect 10364 23418 10420 23420
rect 10444 23418 10500 23420
rect 10524 23418 10580 23420
rect 10604 23418 10660 23420
rect 10684 23418 10740 23420
rect 10364 23366 10366 23418
rect 10366 23366 10418 23418
rect 10418 23366 10420 23418
rect 10444 23366 10482 23418
rect 10482 23366 10494 23418
rect 10494 23366 10500 23418
rect 10524 23366 10546 23418
rect 10546 23366 10558 23418
rect 10558 23366 10580 23418
rect 10604 23366 10610 23418
rect 10610 23366 10622 23418
rect 10622 23366 10660 23418
rect 10684 23366 10686 23418
rect 10686 23366 10738 23418
rect 10738 23366 10740 23418
rect 10364 23364 10420 23366
rect 10444 23364 10500 23366
rect 10524 23364 10580 23366
rect 10604 23364 10660 23366
rect 10684 23364 10740 23366
rect 10782 22616 10838 22672
rect 10046 22480 10102 22536
rect 9678 22344 9734 22400
rect 9402 21936 9458 21992
rect 9034 20984 9090 21040
rect 8758 20712 8814 20768
rect 8574 20168 8630 20224
rect 8666 19236 8722 19272
rect 8666 19216 8668 19236
rect 8668 19216 8720 19236
rect 8720 19216 8722 19236
rect 6642 17856 6698 17912
rect 6366 17620 6368 17640
rect 6368 17620 6420 17640
rect 6420 17620 6422 17640
rect 6366 17584 6422 17620
rect 6274 16904 6330 16960
rect 5998 15680 6054 15736
rect 5446 15544 5502 15600
rect 5262 14864 5318 14920
rect 6366 16632 6422 16688
rect 7378 17856 7434 17912
rect 6918 17584 6974 17640
rect 7654 17992 7710 18048
rect 7010 17060 7066 17096
rect 7010 17040 7012 17060
rect 7012 17040 7064 17060
rect 7064 17040 7066 17060
rect 6734 16108 6790 16144
rect 6734 16088 6736 16108
rect 6736 16088 6788 16108
rect 6788 16088 6790 16108
rect 5262 14456 5318 14512
rect 4364 12538 4420 12540
rect 4444 12538 4500 12540
rect 4524 12538 4580 12540
rect 4604 12538 4660 12540
rect 4684 12538 4740 12540
rect 4364 12486 4366 12538
rect 4366 12486 4418 12538
rect 4418 12486 4420 12538
rect 4444 12486 4482 12538
rect 4482 12486 4494 12538
rect 4494 12486 4500 12538
rect 4524 12486 4546 12538
rect 4546 12486 4558 12538
rect 4558 12486 4580 12538
rect 4604 12486 4610 12538
rect 4610 12486 4622 12538
rect 4622 12486 4660 12538
rect 4684 12486 4686 12538
rect 4686 12486 4738 12538
rect 4738 12486 4740 12538
rect 4364 12484 4420 12486
rect 4444 12484 4500 12486
rect 4524 12484 4580 12486
rect 4604 12484 4660 12486
rect 4684 12484 4740 12486
rect 4250 11756 4306 11792
rect 4250 11736 4252 11756
rect 4252 11736 4304 11756
rect 4304 11736 4306 11756
rect 4364 11450 4420 11452
rect 4444 11450 4500 11452
rect 4524 11450 4580 11452
rect 4604 11450 4660 11452
rect 4684 11450 4740 11452
rect 4364 11398 4366 11450
rect 4366 11398 4418 11450
rect 4418 11398 4420 11450
rect 4444 11398 4482 11450
rect 4482 11398 4494 11450
rect 4494 11398 4500 11450
rect 4524 11398 4546 11450
rect 4546 11398 4558 11450
rect 4558 11398 4580 11450
rect 4604 11398 4610 11450
rect 4610 11398 4622 11450
rect 4622 11398 4660 11450
rect 4684 11398 4686 11450
rect 4686 11398 4738 11450
rect 4738 11398 4740 11450
rect 4364 11396 4420 11398
rect 4444 11396 4500 11398
rect 4524 11396 4580 11398
rect 4604 11396 4660 11398
rect 4684 11396 4740 11398
rect 4364 10362 4420 10364
rect 4444 10362 4500 10364
rect 4524 10362 4580 10364
rect 4604 10362 4660 10364
rect 4684 10362 4740 10364
rect 4364 10310 4366 10362
rect 4366 10310 4418 10362
rect 4418 10310 4420 10362
rect 4444 10310 4482 10362
rect 4482 10310 4494 10362
rect 4494 10310 4500 10362
rect 4524 10310 4546 10362
rect 4546 10310 4558 10362
rect 4558 10310 4580 10362
rect 4604 10310 4610 10362
rect 4610 10310 4622 10362
rect 4622 10310 4660 10362
rect 4684 10310 4686 10362
rect 4686 10310 4738 10362
rect 4738 10310 4740 10362
rect 4364 10308 4420 10310
rect 4444 10308 4500 10310
rect 4524 10308 4580 10310
rect 4604 10308 4660 10310
rect 4684 10308 4740 10310
rect 4342 10104 4398 10160
rect 4066 9596 4068 9616
rect 4068 9596 4120 9616
rect 4120 9596 4122 9616
rect 4066 9560 4122 9596
rect 3974 9152 4030 9208
rect 5538 14320 5594 14376
rect 5538 13776 5594 13832
rect 4364 9274 4420 9276
rect 4444 9274 4500 9276
rect 4524 9274 4580 9276
rect 4604 9274 4660 9276
rect 4684 9274 4740 9276
rect 4364 9222 4366 9274
rect 4366 9222 4418 9274
rect 4418 9222 4420 9274
rect 4444 9222 4482 9274
rect 4482 9222 4494 9274
rect 4494 9222 4500 9274
rect 4524 9222 4546 9274
rect 4546 9222 4558 9274
rect 4558 9222 4580 9274
rect 4604 9222 4610 9274
rect 4610 9222 4622 9274
rect 4622 9222 4660 9274
rect 4684 9222 4686 9274
rect 4686 9222 4738 9274
rect 4738 9222 4740 9274
rect 4364 9220 4420 9222
rect 4444 9220 4500 9222
rect 4524 9220 4580 9222
rect 4604 9220 4660 9222
rect 4684 9220 4740 9222
rect 3606 5616 3662 5672
rect 1364 1114 1420 1116
rect 1444 1114 1500 1116
rect 1524 1114 1580 1116
rect 1604 1114 1660 1116
rect 1684 1114 1740 1116
rect 1364 1062 1366 1114
rect 1366 1062 1418 1114
rect 1418 1062 1420 1114
rect 1444 1062 1482 1114
rect 1482 1062 1494 1114
rect 1494 1062 1500 1114
rect 1524 1062 1546 1114
rect 1546 1062 1558 1114
rect 1558 1062 1580 1114
rect 1604 1062 1610 1114
rect 1610 1062 1622 1114
rect 1622 1062 1660 1114
rect 1684 1062 1686 1114
rect 1686 1062 1738 1114
rect 1738 1062 1740 1114
rect 1364 1060 1420 1062
rect 1444 1060 1500 1062
rect 1524 1060 1580 1062
rect 1604 1060 1660 1062
rect 1684 1060 1740 1062
rect 3698 4684 3754 4720
rect 3698 4664 3700 4684
rect 3700 4664 3752 4684
rect 3752 4664 3754 4684
rect 4802 8628 4858 8664
rect 4802 8608 4804 8628
rect 4804 8608 4856 8628
rect 4856 8608 4858 8628
rect 4364 8186 4420 8188
rect 4444 8186 4500 8188
rect 4524 8186 4580 8188
rect 4604 8186 4660 8188
rect 4684 8186 4740 8188
rect 4364 8134 4366 8186
rect 4366 8134 4418 8186
rect 4418 8134 4420 8186
rect 4444 8134 4482 8186
rect 4482 8134 4494 8186
rect 4494 8134 4500 8186
rect 4524 8134 4546 8186
rect 4546 8134 4558 8186
rect 4558 8134 4580 8186
rect 4604 8134 4610 8186
rect 4610 8134 4622 8186
rect 4622 8134 4660 8186
rect 4684 8134 4686 8186
rect 4686 8134 4738 8186
rect 4738 8134 4740 8186
rect 4364 8132 4420 8134
rect 4444 8132 4500 8134
rect 4524 8132 4580 8134
rect 4604 8132 4660 8134
rect 4684 8132 4740 8134
rect 4894 8372 4896 8392
rect 4896 8372 4948 8392
rect 4948 8372 4950 8392
rect 4894 8336 4950 8372
rect 4364 7098 4420 7100
rect 4444 7098 4500 7100
rect 4524 7098 4580 7100
rect 4604 7098 4660 7100
rect 4684 7098 4740 7100
rect 4364 7046 4366 7098
rect 4366 7046 4418 7098
rect 4418 7046 4420 7098
rect 4444 7046 4482 7098
rect 4482 7046 4494 7098
rect 4494 7046 4500 7098
rect 4524 7046 4546 7098
rect 4546 7046 4558 7098
rect 4558 7046 4580 7098
rect 4604 7046 4610 7098
rect 4610 7046 4622 7098
rect 4622 7046 4660 7098
rect 4684 7046 4686 7098
rect 4686 7046 4738 7098
rect 4738 7046 4740 7098
rect 4364 7044 4420 7046
rect 4444 7044 4500 7046
rect 4524 7044 4580 7046
rect 4604 7044 4660 7046
rect 4684 7044 4740 7046
rect 4364 6010 4420 6012
rect 4444 6010 4500 6012
rect 4524 6010 4580 6012
rect 4604 6010 4660 6012
rect 4684 6010 4740 6012
rect 4364 5958 4366 6010
rect 4366 5958 4418 6010
rect 4418 5958 4420 6010
rect 4444 5958 4482 6010
rect 4482 5958 4494 6010
rect 4494 5958 4500 6010
rect 4524 5958 4546 6010
rect 4546 5958 4558 6010
rect 4558 5958 4580 6010
rect 4604 5958 4610 6010
rect 4610 5958 4622 6010
rect 4622 5958 4660 6010
rect 4684 5958 4686 6010
rect 4686 5958 4738 6010
rect 4738 5958 4740 6010
rect 4364 5956 4420 5958
rect 4444 5956 4500 5958
rect 4524 5956 4580 5958
rect 4604 5956 4660 5958
rect 4684 5956 4740 5958
rect 4342 5072 4398 5128
rect 4364 4922 4420 4924
rect 4444 4922 4500 4924
rect 4524 4922 4580 4924
rect 4604 4922 4660 4924
rect 4684 4922 4740 4924
rect 4364 4870 4366 4922
rect 4366 4870 4418 4922
rect 4418 4870 4420 4922
rect 4444 4870 4482 4922
rect 4482 4870 4494 4922
rect 4494 4870 4500 4922
rect 4524 4870 4546 4922
rect 4546 4870 4558 4922
rect 4558 4870 4580 4922
rect 4604 4870 4610 4922
rect 4610 4870 4622 4922
rect 4622 4870 4660 4922
rect 4684 4870 4686 4922
rect 4686 4870 4738 4922
rect 4738 4870 4740 4922
rect 4364 4868 4420 4870
rect 4444 4868 4500 4870
rect 4524 4868 4580 4870
rect 4604 4868 4660 4870
rect 4684 4868 4740 4870
rect 5446 12144 5502 12200
rect 5262 11056 5318 11112
rect 4342 4664 4398 4720
rect 4986 4020 4988 4040
rect 4988 4020 5040 4040
rect 5040 4020 5042 4040
rect 4986 3984 5042 4020
rect 4364 3834 4420 3836
rect 4444 3834 4500 3836
rect 4524 3834 4580 3836
rect 4604 3834 4660 3836
rect 4684 3834 4740 3836
rect 4364 3782 4366 3834
rect 4366 3782 4418 3834
rect 4418 3782 4420 3834
rect 4444 3782 4482 3834
rect 4482 3782 4494 3834
rect 4494 3782 4500 3834
rect 4524 3782 4546 3834
rect 4546 3782 4558 3834
rect 4558 3782 4580 3834
rect 4604 3782 4610 3834
rect 4610 3782 4622 3834
rect 4622 3782 4660 3834
rect 4684 3782 4686 3834
rect 4686 3782 4738 3834
rect 4738 3782 4740 3834
rect 4364 3780 4420 3782
rect 4444 3780 4500 3782
rect 4524 3780 4580 3782
rect 4604 3780 4660 3782
rect 4684 3780 4740 3782
rect 4986 3052 5042 3088
rect 4986 3032 4988 3052
rect 4988 3032 5040 3052
rect 5040 3032 5042 3052
rect 4364 2746 4420 2748
rect 4444 2746 4500 2748
rect 4524 2746 4580 2748
rect 4604 2746 4660 2748
rect 4684 2746 4740 2748
rect 4364 2694 4366 2746
rect 4366 2694 4418 2746
rect 4418 2694 4420 2746
rect 4444 2694 4482 2746
rect 4482 2694 4494 2746
rect 4494 2694 4500 2746
rect 4524 2694 4546 2746
rect 4546 2694 4558 2746
rect 4558 2694 4580 2746
rect 4604 2694 4610 2746
rect 4610 2694 4622 2746
rect 4622 2694 4660 2746
rect 4684 2694 4686 2746
rect 4686 2694 4738 2746
rect 4738 2694 4740 2746
rect 4364 2692 4420 2694
rect 4444 2692 4500 2694
rect 4524 2692 4580 2694
rect 4604 2692 4660 2694
rect 4684 2692 4740 2694
rect 5998 14592 6054 14648
rect 6642 15544 6698 15600
rect 5354 9016 5410 9072
rect 6090 13912 6146 13968
rect 6458 15036 6460 15056
rect 6460 15036 6512 15056
rect 6512 15036 6514 15056
rect 6458 15000 6514 15036
rect 7364 17434 7420 17436
rect 7444 17434 7500 17436
rect 7524 17434 7580 17436
rect 7604 17434 7660 17436
rect 7684 17434 7740 17436
rect 7364 17382 7366 17434
rect 7366 17382 7418 17434
rect 7418 17382 7420 17434
rect 7444 17382 7482 17434
rect 7482 17382 7494 17434
rect 7494 17382 7500 17434
rect 7524 17382 7546 17434
rect 7546 17382 7558 17434
rect 7558 17382 7580 17434
rect 7604 17382 7610 17434
rect 7610 17382 7622 17434
rect 7622 17382 7660 17434
rect 7684 17382 7686 17434
rect 7686 17382 7738 17434
rect 7738 17382 7740 17434
rect 7364 17380 7420 17382
rect 7444 17380 7500 17382
rect 7524 17380 7580 17382
rect 7604 17380 7660 17382
rect 7684 17380 7740 17382
rect 7286 16496 7342 16552
rect 7470 16496 7526 16552
rect 7364 16346 7420 16348
rect 7444 16346 7500 16348
rect 7524 16346 7580 16348
rect 7604 16346 7660 16348
rect 7684 16346 7740 16348
rect 7364 16294 7366 16346
rect 7366 16294 7418 16346
rect 7418 16294 7420 16346
rect 7444 16294 7482 16346
rect 7482 16294 7494 16346
rect 7494 16294 7500 16346
rect 7524 16294 7546 16346
rect 7546 16294 7558 16346
rect 7558 16294 7580 16346
rect 7604 16294 7610 16346
rect 7610 16294 7622 16346
rect 7622 16294 7660 16346
rect 7684 16294 7686 16346
rect 7686 16294 7738 16346
rect 7738 16294 7740 16346
rect 7364 16292 7420 16294
rect 7444 16292 7500 16294
rect 7524 16292 7580 16294
rect 7604 16292 7660 16294
rect 7684 16292 7740 16294
rect 6826 13232 6882 13288
rect 5630 8880 5686 8936
rect 5538 6976 5594 7032
rect 5722 8628 5778 8664
rect 5722 8608 5724 8628
rect 5724 8608 5776 8628
rect 5776 8608 5778 8628
rect 6550 10648 6606 10704
rect 6274 9016 6330 9072
rect 6274 7948 6330 7984
rect 6274 7928 6276 7948
rect 6276 7928 6328 7948
rect 6328 7928 6330 7948
rect 6366 7384 6422 7440
rect 6550 9016 6606 9072
rect 6550 7248 6606 7304
rect 6458 6976 6514 7032
rect 6458 6724 6514 6760
rect 6458 6704 6460 6724
rect 6460 6704 6512 6724
rect 6512 6704 6514 6724
rect 4364 1658 4420 1660
rect 4444 1658 4500 1660
rect 4524 1658 4580 1660
rect 4604 1658 4660 1660
rect 4684 1658 4740 1660
rect 4364 1606 4366 1658
rect 4366 1606 4418 1658
rect 4418 1606 4420 1658
rect 4444 1606 4482 1658
rect 4482 1606 4494 1658
rect 4494 1606 4500 1658
rect 4524 1606 4546 1658
rect 4546 1606 4558 1658
rect 4558 1606 4580 1658
rect 4604 1606 4610 1658
rect 4610 1606 4622 1658
rect 4622 1606 4660 1658
rect 4684 1606 4686 1658
rect 4686 1606 4738 1658
rect 4738 1606 4740 1658
rect 4364 1604 4420 1606
rect 4444 1604 4500 1606
rect 4524 1604 4580 1606
rect 4604 1604 4660 1606
rect 4684 1604 4740 1606
rect 4526 756 4528 776
rect 4528 756 4580 776
rect 4580 756 4582 776
rect 4526 720 4582 756
rect 4364 570 4420 572
rect 4444 570 4500 572
rect 4524 570 4580 572
rect 4604 570 4660 572
rect 4684 570 4740 572
rect 4364 518 4366 570
rect 4366 518 4418 570
rect 4418 518 4420 570
rect 4444 518 4482 570
rect 4482 518 4494 570
rect 4494 518 4500 570
rect 4524 518 4546 570
rect 4546 518 4558 570
rect 4558 518 4580 570
rect 4604 518 4610 570
rect 4610 518 4622 570
rect 4622 518 4660 570
rect 4684 518 4686 570
rect 4686 518 4738 570
rect 4738 518 4740 570
rect 4364 516 4420 518
rect 4444 516 4500 518
rect 4524 516 4580 518
rect 4604 516 4660 518
rect 4684 516 4740 518
rect 5446 1536 5502 1592
rect 7378 15564 7434 15600
rect 7378 15544 7380 15564
rect 7380 15544 7432 15564
rect 7432 15544 7434 15564
rect 7364 15258 7420 15260
rect 7444 15258 7500 15260
rect 7524 15258 7580 15260
rect 7604 15258 7660 15260
rect 7684 15258 7740 15260
rect 7364 15206 7366 15258
rect 7366 15206 7418 15258
rect 7418 15206 7420 15258
rect 7444 15206 7482 15258
rect 7482 15206 7494 15258
rect 7494 15206 7500 15258
rect 7524 15206 7546 15258
rect 7546 15206 7558 15258
rect 7558 15206 7580 15258
rect 7604 15206 7610 15258
rect 7610 15206 7622 15258
rect 7622 15206 7660 15258
rect 7684 15206 7686 15258
rect 7686 15206 7738 15258
rect 7738 15206 7740 15258
rect 7364 15204 7420 15206
rect 7444 15204 7500 15206
rect 7524 15204 7580 15206
rect 7604 15204 7660 15206
rect 7684 15204 7740 15206
rect 7364 14170 7420 14172
rect 7444 14170 7500 14172
rect 7524 14170 7580 14172
rect 7604 14170 7660 14172
rect 7684 14170 7740 14172
rect 7364 14118 7366 14170
rect 7366 14118 7418 14170
rect 7418 14118 7420 14170
rect 7444 14118 7482 14170
rect 7482 14118 7494 14170
rect 7494 14118 7500 14170
rect 7524 14118 7546 14170
rect 7546 14118 7558 14170
rect 7558 14118 7580 14170
rect 7604 14118 7610 14170
rect 7610 14118 7622 14170
rect 7622 14118 7660 14170
rect 7684 14118 7686 14170
rect 7686 14118 7738 14170
rect 7738 14118 7740 14170
rect 7364 14116 7420 14118
rect 7444 14116 7500 14118
rect 7524 14116 7580 14118
rect 7604 14116 7660 14118
rect 7684 14116 7740 14118
rect 7378 13912 7434 13968
rect 7654 13268 7656 13288
rect 7656 13268 7708 13288
rect 7708 13268 7710 13288
rect 7654 13232 7710 13268
rect 7364 13082 7420 13084
rect 7444 13082 7500 13084
rect 7524 13082 7580 13084
rect 7604 13082 7660 13084
rect 7684 13082 7740 13084
rect 7364 13030 7366 13082
rect 7366 13030 7418 13082
rect 7418 13030 7420 13082
rect 7444 13030 7482 13082
rect 7482 13030 7494 13082
rect 7494 13030 7500 13082
rect 7524 13030 7546 13082
rect 7546 13030 7558 13082
rect 7558 13030 7580 13082
rect 7604 13030 7610 13082
rect 7610 13030 7622 13082
rect 7622 13030 7660 13082
rect 7684 13030 7686 13082
rect 7686 13030 7738 13082
rect 7738 13030 7740 13082
rect 7364 13028 7420 13030
rect 7444 13028 7500 13030
rect 7524 13028 7580 13030
rect 7604 13028 7660 13030
rect 7684 13028 7740 13030
rect 7364 11994 7420 11996
rect 7444 11994 7500 11996
rect 7524 11994 7580 11996
rect 7604 11994 7660 11996
rect 7684 11994 7740 11996
rect 7364 11942 7366 11994
rect 7366 11942 7418 11994
rect 7418 11942 7420 11994
rect 7444 11942 7482 11994
rect 7482 11942 7494 11994
rect 7494 11942 7500 11994
rect 7524 11942 7546 11994
rect 7546 11942 7558 11994
rect 7558 11942 7580 11994
rect 7604 11942 7610 11994
rect 7610 11942 7622 11994
rect 7622 11942 7660 11994
rect 7684 11942 7686 11994
rect 7686 11942 7738 11994
rect 7738 11942 7740 11994
rect 7364 11940 7420 11942
rect 7444 11940 7500 11942
rect 7524 11940 7580 11942
rect 7604 11940 7660 11942
rect 7684 11940 7740 11942
rect 7838 11056 7894 11112
rect 7364 10906 7420 10908
rect 7444 10906 7500 10908
rect 7524 10906 7580 10908
rect 7604 10906 7660 10908
rect 7684 10906 7740 10908
rect 7364 10854 7366 10906
rect 7366 10854 7418 10906
rect 7418 10854 7420 10906
rect 7444 10854 7482 10906
rect 7482 10854 7494 10906
rect 7494 10854 7500 10906
rect 7524 10854 7546 10906
rect 7546 10854 7558 10906
rect 7558 10854 7580 10906
rect 7604 10854 7610 10906
rect 7610 10854 7622 10906
rect 7622 10854 7660 10906
rect 7684 10854 7686 10906
rect 7686 10854 7738 10906
rect 7738 10854 7740 10906
rect 7364 10852 7420 10854
rect 7444 10852 7500 10854
rect 7524 10852 7580 10854
rect 7604 10852 7660 10854
rect 7684 10852 7740 10854
rect 6734 10104 6790 10160
rect 6918 9968 6974 10024
rect 6734 7384 6790 7440
rect 6826 7112 6882 7168
rect 7364 9818 7420 9820
rect 7444 9818 7500 9820
rect 7524 9818 7580 9820
rect 7604 9818 7660 9820
rect 7684 9818 7740 9820
rect 7364 9766 7366 9818
rect 7366 9766 7418 9818
rect 7418 9766 7420 9818
rect 7444 9766 7482 9818
rect 7482 9766 7494 9818
rect 7494 9766 7500 9818
rect 7524 9766 7546 9818
rect 7546 9766 7558 9818
rect 7558 9766 7580 9818
rect 7604 9766 7610 9818
rect 7610 9766 7622 9818
rect 7622 9766 7660 9818
rect 7684 9766 7686 9818
rect 7686 9766 7738 9818
rect 7738 9766 7740 9818
rect 7364 9764 7420 9766
rect 7444 9764 7500 9766
rect 7524 9764 7580 9766
rect 7604 9764 7660 9766
rect 7684 9764 7740 9766
rect 7654 9152 7710 9208
rect 7102 8880 7158 8936
rect 7838 8744 7894 8800
rect 7364 8730 7420 8732
rect 7444 8730 7500 8732
rect 7524 8730 7580 8732
rect 7604 8730 7660 8732
rect 7684 8730 7740 8732
rect 7364 8678 7366 8730
rect 7366 8678 7418 8730
rect 7418 8678 7420 8730
rect 7444 8678 7482 8730
rect 7482 8678 7494 8730
rect 7494 8678 7500 8730
rect 7524 8678 7546 8730
rect 7546 8678 7558 8730
rect 7558 8678 7580 8730
rect 7604 8678 7610 8730
rect 7610 8678 7622 8730
rect 7622 8678 7660 8730
rect 7684 8678 7686 8730
rect 7686 8678 7738 8730
rect 7738 8678 7740 8730
rect 7364 8676 7420 8678
rect 7444 8676 7500 8678
rect 7524 8676 7580 8678
rect 7604 8676 7660 8678
rect 7684 8676 7740 8678
rect 7470 7792 7526 7848
rect 8298 15816 8354 15872
rect 8298 15408 8354 15464
rect 8206 14728 8262 14784
rect 8666 16632 8722 16688
rect 8482 14728 8538 14784
rect 8298 14456 8354 14512
rect 8114 13948 8116 13968
rect 8116 13948 8168 13968
rect 8168 13948 8170 13968
rect 8114 13912 8170 13948
rect 8022 13640 8078 13696
rect 8298 12688 8354 12744
rect 8758 15680 8814 15736
rect 9126 19216 9182 19272
rect 9218 19080 9274 19136
rect 10046 21392 10102 21448
rect 9586 20712 9642 20768
rect 9862 20848 9918 20904
rect 9954 20576 10010 20632
rect 10364 22330 10420 22332
rect 10444 22330 10500 22332
rect 10524 22330 10580 22332
rect 10604 22330 10660 22332
rect 10684 22330 10740 22332
rect 10364 22278 10366 22330
rect 10366 22278 10418 22330
rect 10418 22278 10420 22330
rect 10444 22278 10482 22330
rect 10482 22278 10494 22330
rect 10494 22278 10500 22330
rect 10524 22278 10546 22330
rect 10546 22278 10558 22330
rect 10558 22278 10580 22330
rect 10604 22278 10610 22330
rect 10610 22278 10622 22330
rect 10622 22278 10660 22330
rect 10684 22278 10686 22330
rect 10686 22278 10738 22330
rect 10738 22278 10740 22330
rect 10364 22276 10420 22278
rect 10444 22276 10500 22278
rect 10524 22276 10580 22278
rect 10604 22276 10660 22278
rect 10684 22276 10740 22278
rect 11150 21528 11206 21584
rect 10364 21242 10420 21244
rect 10444 21242 10500 21244
rect 10524 21242 10580 21244
rect 10604 21242 10660 21244
rect 10684 21242 10740 21244
rect 10364 21190 10366 21242
rect 10366 21190 10418 21242
rect 10418 21190 10420 21242
rect 10444 21190 10482 21242
rect 10482 21190 10494 21242
rect 10494 21190 10500 21242
rect 10524 21190 10546 21242
rect 10546 21190 10558 21242
rect 10558 21190 10580 21242
rect 10604 21190 10610 21242
rect 10610 21190 10622 21242
rect 10622 21190 10660 21242
rect 10684 21190 10686 21242
rect 10686 21190 10738 21242
rect 10738 21190 10740 21242
rect 10364 21188 10420 21190
rect 10444 21188 10500 21190
rect 10524 21188 10580 21190
rect 10604 21188 10660 21190
rect 10684 21188 10740 21190
rect 9678 19488 9734 19544
rect 9862 19116 9864 19136
rect 9864 19116 9916 19136
rect 9916 19116 9918 19136
rect 9862 19080 9918 19116
rect 9310 18264 9366 18320
rect 9310 18128 9366 18184
rect 9218 17992 9274 18048
rect 9310 17720 9366 17776
rect 8942 16668 8944 16688
rect 8944 16668 8996 16688
rect 8996 16668 8998 16688
rect 8942 16632 8998 16668
rect 8942 15272 8998 15328
rect 8850 14864 8906 14920
rect 10364 20154 10420 20156
rect 10444 20154 10500 20156
rect 10524 20154 10580 20156
rect 10604 20154 10660 20156
rect 10684 20154 10740 20156
rect 10364 20102 10366 20154
rect 10366 20102 10418 20154
rect 10418 20102 10420 20154
rect 10444 20102 10482 20154
rect 10482 20102 10494 20154
rect 10494 20102 10500 20154
rect 10524 20102 10546 20154
rect 10546 20102 10558 20154
rect 10558 20102 10580 20154
rect 10604 20102 10610 20154
rect 10610 20102 10622 20154
rect 10622 20102 10660 20154
rect 10684 20102 10686 20154
rect 10686 20102 10738 20154
rect 10738 20102 10740 20154
rect 10364 20100 10420 20102
rect 10444 20100 10500 20102
rect 10524 20100 10580 20102
rect 10604 20100 10660 20102
rect 10684 20100 10740 20102
rect 10506 19624 10562 19680
rect 10966 20168 11022 20224
rect 10364 19066 10420 19068
rect 10444 19066 10500 19068
rect 10524 19066 10580 19068
rect 10604 19066 10660 19068
rect 10684 19066 10740 19068
rect 10364 19014 10366 19066
rect 10366 19014 10418 19066
rect 10418 19014 10420 19066
rect 10444 19014 10482 19066
rect 10482 19014 10494 19066
rect 10494 19014 10500 19066
rect 10524 19014 10546 19066
rect 10546 19014 10558 19066
rect 10558 19014 10580 19066
rect 10604 19014 10610 19066
rect 10610 19014 10622 19066
rect 10622 19014 10660 19066
rect 10684 19014 10686 19066
rect 10686 19014 10738 19066
rect 10738 19014 10740 19066
rect 10364 19012 10420 19014
rect 10444 19012 10500 19014
rect 10524 19012 10580 19014
rect 10604 19012 10660 19014
rect 10684 19012 10740 19014
rect 10230 18264 10286 18320
rect 9494 15816 9550 15872
rect 10364 17978 10420 17980
rect 10444 17978 10500 17980
rect 10524 17978 10580 17980
rect 10604 17978 10660 17980
rect 10684 17978 10740 17980
rect 10364 17926 10366 17978
rect 10366 17926 10418 17978
rect 10418 17926 10420 17978
rect 10444 17926 10482 17978
rect 10482 17926 10494 17978
rect 10494 17926 10500 17978
rect 10524 17926 10546 17978
rect 10546 17926 10558 17978
rect 10558 17926 10580 17978
rect 10604 17926 10610 17978
rect 10610 17926 10622 17978
rect 10622 17926 10660 17978
rect 10684 17926 10686 17978
rect 10686 17926 10738 17978
rect 10738 17926 10740 17978
rect 10364 17924 10420 17926
rect 10444 17924 10500 17926
rect 10524 17924 10580 17926
rect 10604 17924 10660 17926
rect 10684 17924 10740 17926
rect 13174 21936 13230 21992
rect 16364 23418 16420 23420
rect 16444 23418 16500 23420
rect 16524 23418 16580 23420
rect 16604 23418 16660 23420
rect 16684 23418 16740 23420
rect 16364 23366 16366 23418
rect 16366 23366 16418 23418
rect 16418 23366 16420 23418
rect 16444 23366 16482 23418
rect 16482 23366 16494 23418
rect 16494 23366 16500 23418
rect 16524 23366 16546 23418
rect 16546 23366 16558 23418
rect 16558 23366 16580 23418
rect 16604 23366 16610 23418
rect 16610 23366 16622 23418
rect 16622 23366 16660 23418
rect 16684 23366 16686 23418
rect 16686 23366 16738 23418
rect 16738 23366 16740 23418
rect 16364 23364 16420 23366
rect 16444 23364 16500 23366
rect 16524 23364 16580 23366
rect 16604 23364 16660 23366
rect 16684 23364 16740 23366
rect 13364 22874 13420 22876
rect 13444 22874 13500 22876
rect 13524 22874 13580 22876
rect 13604 22874 13660 22876
rect 13684 22874 13740 22876
rect 13364 22822 13366 22874
rect 13366 22822 13418 22874
rect 13418 22822 13420 22874
rect 13444 22822 13482 22874
rect 13482 22822 13494 22874
rect 13494 22822 13500 22874
rect 13524 22822 13546 22874
rect 13546 22822 13558 22874
rect 13558 22822 13580 22874
rect 13604 22822 13610 22874
rect 13610 22822 13622 22874
rect 13622 22822 13660 22874
rect 13684 22822 13686 22874
rect 13686 22822 13738 22874
rect 13738 22822 13740 22874
rect 13364 22820 13420 22822
rect 13444 22820 13500 22822
rect 13524 22820 13580 22822
rect 13604 22820 13660 22822
rect 13684 22820 13740 22822
rect 12530 21836 12532 21856
rect 12532 21836 12584 21856
rect 12584 21836 12586 21856
rect 11518 20848 11574 20904
rect 11426 20440 11482 20496
rect 12530 21800 12586 21836
rect 13818 21800 13874 21856
rect 13364 21786 13420 21788
rect 13444 21786 13500 21788
rect 13524 21786 13580 21788
rect 13604 21786 13660 21788
rect 13684 21786 13740 21788
rect 13364 21734 13366 21786
rect 13366 21734 13418 21786
rect 13418 21734 13420 21786
rect 13444 21734 13482 21786
rect 13482 21734 13494 21786
rect 13494 21734 13500 21786
rect 13524 21734 13546 21786
rect 13546 21734 13558 21786
rect 13558 21734 13580 21786
rect 13604 21734 13610 21786
rect 13610 21734 13622 21786
rect 13622 21734 13660 21786
rect 13684 21734 13686 21786
rect 13686 21734 13738 21786
rect 13738 21734 13740 21786
rect 13364 21732 13420 21734
rect 13444 21732 13500 21734
rect 13524 21732 13580 21734
rect 13604 21732 13660 21734
rect 13684 21732 13740 21734
rect 13910 21392 13966 21448
rect 12622 20848 12678 20904
rect 12530 20748 12532 20768
rect 12532 20748 12584 20768
rect 12584 20748 12586 20768
rect 12530 20712 12586 20748
rect 12806 20712 12862 20768
rect 13364 20698 13420 20700
rect 13444 20698 13500 20700
rect 13524 20698 13580 20700
rect 13604 20698 13660 20700
rect 13684 20698 13740 20700
rect 13364 20646 13366 20698
rect 13366 20646 13418 20698
rect 13418 20646 13420 20698
rect 13444 20646 13482 20698
rect 13482 20646 13494 20698
rect 13494 20646 13500 20698
rect 13524 20646 13546 20698
rect 13546 20646 13558 20698
rect 13558 20646 13580 20698
rect 13604 20646 13610 20698
rect 13610 20646 13622 20698
rect 13622 20646 13660 20698
rect 13684 20646 13686 20698
rect 13686 20646 13738 20698
rect 13738 20646 13740 20698
rect 13364 20644 13420 20646
rect 13444 20644 13500 20646
rect 13524 20644 13580 20646
rect 13604 20644 13660 20646
rect 13684 20644 13740 20646
rect 15106 22072 15162 22128
rect 10364 16890 10420 16892
rect 10444 16890 10500 16892
rect 10524 16890 10580 16892
rect 10604 16890 10660 16892
rect 10684 16890 10740 16892
rect 10364 16838 10366 16890
rect 10366 16838 10418 16890
rect 10418 16838 10420 16890
rect 10444 16838 10482 16890
rect 10482 16838 10494 16890
rect 10494 16838 10500 16890
rect 10524 16838 10546 16890
rect 10546 16838 10558 16890
rect 10558 16838 10580 16890
rect 10604 16838 10610 16890
rect 10610 16838 10622 16890
rect 10622 16838 10660 16890
rect 10684 16838 10686 16890
rect 10686 16838 10738 16890
rect 10738 16838 10740 16890
rect 10364 16836 10420 16838
rect 10444 16836 10500 16838
rect 10524 16836 10580 16838
rect 10604 16836 10660 16838
rect 10684 16836 10740 16838
rect 10598 16652 10654 16688
rect 10598 16632 10600 16652
rect 10600 16632 10652 16652
rect 10652 16632 10654 16652
rect 9034 14456 9090 14512
rect 8942 13504 8998 13560
rect 8574 12688 8630 12744
rect 7364 7642 7420 7644
rect 7444 7642 7500 7644
rect 7524 7642 7580 7644
rect 7604 7642 7660 7644
rect 7684 7642 7740 7644
rect 7364 7590 7366 7642
rect 7366 7590 7418 7642
rect 7418 7590 7420 7642
rect 7444 7590 7482 7642
rect 7482 7590 7494 7642
rect 7494 7590 7500 7642
rect 7524 7590 7546 7642
rect 7546 7590 7558 7642
rect 7558 7590 7580 7642
rect 7604 7590 7610 7642
rect 7610 7590 7622 7642
rect 7622 7590 7660 7642
rect 7684 7590 7686 7642
rect 7686 7590 7738 7642
rect 7738 7590 7740 7642
rect 7364 7588 7420 7590
rect 7444 7588 7500 7590
rect 7524 7588 7580 7590
rect 7604 7588 7660 7590
rect 7684 7588 7740 7590
rect 7194 6432 7250 6488
rect 7364 6554 7420 6556
rect 7444 6554 7500 6556
rect 7524 6554 7580 6556
rect 7604 6554 7660 6556
rect 7684 6554 7740 6556
rect 7364 6502 7366 6554
rect 7366 6502 7418 6554
rect 7418 6502 7420 6554
rect 7444 6502 7482 6554
rect 7482 6502 7494 6554
rect 7494 6502 7500 6554
rect 7524 6502 7546 6554
rect 7546 6502 7558 6554
rect 7558 6502 7580 6554
rect 7604 6502 7610 6554
rect 7610 6502 7622 6554
rect 7622 6502 7660 6554
rect 7684 6502 7686 6554
rect 7686 6502 7738 6554
rect 7738 6502 7740 6554
rect 7364 6500 7420 6502
rect 7444 6500 7500 6502
rect 7524 6500 7580 6502
rect 7604 6500 7660 6502
rect 7684 6500 7740 6502
rect 7746 6024 7802 6080
rect 7364 5466 7420 5468
rect 7444 5466 7500 5468
rect 7524 5466 7580 5468
rect 7604 5466 7660 5468
rect 7684 5466 7740 5468
rect 7364 5414 7366 5466
rect 7366 5414 7418 5466
rect 7418 5414 7420 5466
rect 7444 5414 7482 5466
rect 7482 5414 7494 5466
rect 7494 5414 7500 5466
rect 7524 5414 7546 5466
rect 7546 5414 7558 5466
rect 7558 5414 7580 5466
rect 7604 5414 7610 5466
rect 7610 5414 7622 5466
rect 7622 5414 7660 5466
rect 7684 5414 7686 5466
rect 7686 5414 7738 5466
rect 7738 5414 7740 5466
rect 7364 5412 7420 5414
rect 7444 5412 7500 5414
rect 7524 5412 7580 5414
rect 7604 5412 7660 5414
rect 7684 5412 7740 5414
rect 7364 4378 7420 4380
rect 7444 4378 7500 4380
rect 7524 4378 7580 4380
rect 7604 4378 7660 4380
rect 7684 4378 7740 4380
rect 7364 4326 7366 4378
rect 7366 4326 7418 4378
rect 7418 4326 7420 4378
rect 7444 4326 7482 4378
rect 7482 4326 7494 4378
rect 7494 4326 7500 4378
rect 7524 4326 7546 4378
rect 7546 4326 7558 4378
rect 7558 4326 7580 4378
rect 7604 4326 7610 4378
rect 7610 4326 7622 4378
rect 7622 4326 7660 4378
rect 7684 4326 7686 4378
rect 7686 4326 7738 4378
rect 7738 4326 7740 4378
rect 7364 4324 7420 4326
rect 7444 4324 7500 4326
rect 7524 4324 7580 4326
rect 7604 4324 7660 4326
rect 7684 4324 7740 4326
rect 8390 12144 8446 12200
rect 8298 11192 8354 11248
rect 8206 10648 8262 10704
rect 8206 9968 8262 10024
rect 8758 10512 8814 10568
rect 8114 8916 8116 8936
rect 8116 8916 8168 8936
rect 8168 8916 8170 8936
rect 8114 8880 8170 8916
rect 8390 7928 8446 7984
rect 8114 6160 8170 6216
rect 8390 7384 8446 7440
rect 8666 8472 8722 8528
rect 9218 14728 9274 14784
rect 9218 12180 9220 12200
rect 9220 12180 9272 12200
rect 9272 12180 9274 12200
rect 9218 12144 9274 12180
rect 9126 10784 9182 10840
rect 9034 10240 9090 10296
rect 9218 9968 9274 10024
rect 9126 9696 9182 9752
rect 9586 14592 9642 14648
rect 9770 14456 9826 14512
rect 9494 13640 9550 13696
rect 9310 9560 9366 9616
rect 8942 7928 8998 7984
rect 9770 12960 9826 13016
rect 9770 12824 9826 12880
rect 10364 15802 10420 15804
rect 10444 15802 10500 15804
rect 10524 15802 10580 15804
rect 10604 15802 10660 15804
rect 10684 15802 10740 15804
rect 10364 15750 10366 15802
rect 10366 15750 10418 15802
rect 10418 15750 10420 15802
rect 10444 15750 10482 15802
rect 10482 15750 10494 15802
rect 10494 15750 10500 15802
rect 10524 15750 10546 15802
rect 10546 15750 10558 15802
rect 10558 15750 10580 15802
rect 10604 15750 10610 15802
rect 10610 15750 10622 15802
rect 10622 15750 10660 15802
rect 10684 15750 10686 15802
rect 10686 15750 10738 15802
rect 10738 15750 10740 15802
rect 10364 15748 10420 15750
rect 10444 15748 10500 15750
rect 10524 15748 10580 15750
rect 10604 15748 10660 15750
rect 10684 15748 10740 15750
rect 10046 15000 10102 15056
rect 10138 14592 10194 14648
rect 10138 14340 10194 14376
rect 10138 14320 10140 14340
rect 10140 14320 10192 14340
rect 10192 14320 10194 14340
rect 10598 15000 10654 15056
rect 10364 14714 10420 14716
rect 10444 14714 10500 14716
rect 10524 14714 10580 14716
rect 10604 14714 10660 14716
rect 10684 14714 10740 14716
rect 10364 14662 10366 14714
rect 10366 14662 10418 14714
rect 10418 14662 10420 14714
rect 10444 14662 10482 14714
rect 10482 14662 10494 14714
rect 10494 14662 10500 14714
rect 10524 14662 10546 14714
rect 10546 14662 10558 14714
rect 10558 14662 10580 14714
rect 10604 14662 10610 14714
rect 10610 14662 10622 14714
rect 10622 14662 10660 14714
rect 10684 14662 10686 14714
rect 10686 14662 10738 14714
rect 10738 14662 10740 14714
rect 10364 14660 10420 14662
rect 10444 14660 10500 14662
rect 10524 14660 10580 14662
rect 10604 14660 10660 14662
rect 10684 14660 10740 14662
rect 10138 14048 10194 14104
rect 10322 13776 10378 13832
rect 10690 14184 10746 14240
rect 10364 13626 10420 13628
rect 10444 13626 10500 13628
rect 10524 13626 10580 13628
rect 10604 13626 10660 13628
rect 10684 13626 10740 13628
rect 10364 13574 10366 13626
rect 10366 13574 10418 13626
rect 10418 13574 10420 13626
rect 10444 13574 10482 13626
rect 10482 13574 10494 13626
rect 10494 13574 10500 13626
rect 10524 13574 10546 13626
rect 10546 13574 10558 13626
rect 10558 13574 10580 13626
rect 10604 13574 10610 13626
rect 10610 13574 10622 13626
rect 10622 13574 10660 13626
rect 10684 13574 10686 13626
rect 10686 13574 10738 13626
rect 10738 13574 10740 13626
rect 10364 13572 10420 13574
rect 10444 13572 10500 13574
rect 10524 13572 10580 13574
rect 10604 13572 10660 13574
rect 10684 13572 10740 13574
rect 10966 15136 11022 15192
rect 9862 9696 9918 9752
rect 9494 9424 9550 9480
rect 9586 8628 9642 8664
rect 9586 8608 9588 8628
rect 9588 8608 9640 8628
rect 9640 8608 9642 8628
rect 9310 8200 9366 8256
rect 8482 6568 8538 6624
rect 9126 7812 9182 7848
rect 9126 7792 9128 7812
rect 9128 7792 9180 7812
rect 9180 7792 9182 7812
rect 8114 5652 8116 5672
rect 8116 5652 8168 5672
rect 8168 5652 8170 5672
rect 8114 5616 8170 5652
rect 8114 5480 8170 5536
rect 9034 6568 9090 6624
rect 8022 4120 8078 4176
rect 7364 3290 7420 3292
rect 7444 3290 7500 3292
rect 7524 3290 7580 3292
rect 7604 3290 7660 3292
rect 7684 3290 7740 3292
rect 7364 3238 7366 3290
rect 7366 3238 7418 3290
rect 7418 3238 7420 3290
rect 7444 3238 7482 3290
rect 7482 3238 7494 3290
rect 7494 3238 7500 3290
rect 7524 3238 7546 3290
rect 7546 3238 7558 3290
rect 7558 3238 7580 3290
rect 7604 3238 7610 3290
rect 7610 3238 7622 3290
rect 7622 3238 7660 3290
rect 7684 3238 7686 3290
rect 7686 3238 7738 3290
rect 7738 3238 7740 3290
rect 7364 3236 7420 3238
rect 7444 3236 7500 3238
rect 7524 3236 7580 3238
rect 7604 3236 7660 3238
rect 7684 3236 7740 3238
rect 7746 3032 7802 3088
rect 6642 1980 6644 2000
rect 6644 1980 6696 2000
rect 6696 1980 6698 2000
rect 6642 1944 6698 1980
rect 7364 2202 7420 2204
rect 7444 2202 7500 2204
rect 7524 2202 7580 2204
rect 7604 2202 7660 2204
rect 7684 2202 7740 2204
rect 7364 2150 7366 2202
rect 7366 2150 7418 2202
rect 7418 2150 7420 2202
rect 7444 2150 7482 2202
rect 7482 2150 7494 2202
rect 7494 2150 7500 2202
rect 7524 2150 7546 2202
rect 7546 2150 7558 2202
rect 7558 2150 7580 2202
rect 7604 2150 7610 2202
rect 7610 2150 7622 2202
rect 7622 2150 7660 2202
rect 7684 2150 7686 2202
rect 7686 2150 7738 2202
rect 7738 2150 7740 2202
rect 7364 2148 7420 2150
rect 7444 2148 7500 2150
rect 7524 2148 7580 2150
rect 7604 2148 7660 2150
rect 7684 2148 7740 2150
rect 6734 1420 6790 1456
rect 6734 1400 6736 1420
rect 6736 1400 6788 1420
rect 6788 1400 6790 1420
rect 5262 720 5318 776
rect 7364 1114 7420 1116
rect 7444 1114 7500 1116
rect 7524 1114 7580 1116
rect 7604 1114 7660 1116
rect 7684 1114 7740 1116
rect 7364 1062 7366 1114
rect 7366 1062 7418 1114
rect 7418 1062 7420 1114
rect 7444 1062 7482 1114
rect 7482 1062 7494 1114
rect 7494 1062 7500 1114
rect 7524 1062 7546 1114
rect 7546 1062 7558 1114
rect 7558 1062 7580 1114
rect 7604 1062 7610 1114
rect 7610 1062 7622 1114
rect 7622 1062 7660 1114
rect 7684 1062 7686 1114
rect 7686 1062 7738 1114
rect 7738 1062 7740 1114
rect 7364 1060 7420 1062
rect 7444 1060 7500 1062
rect 7524 1060 7580 1062
rect 7604 1060 7660 1062
rect 7684 1060 7740 1062
rect 7102 892 7104 912
rect 7104 892 7156 912
rect 7156 892 7158 912
rect 7102 856 7158 892
rect 9770 8336 9826 8392
rect 9586 7928 9642 7984
rect 9218 6296 9274 6352
rect 9678 7248 9734 7304
rect 9034 3576 9090 3632
rect 9586 6296 9642 6352
rect 9586 2932 9588 2952
rect 9588 2932 9640 2952
rect 9640 2932 9642 2952
rect 9586 2896 9642 2932
rect 10364 12538 10420 12540
rect 10444 12538 10500 12540
rect 10524 12538 10580 12540
rect 10604 12538 10660 12540
rect 10684 12538 10740 12540
rect 10364 12486 10366 12538
rect 10366 12486 10418 12538
rect 10418 12486 10420 12538
rect 10444 12486 10482 12538
rect 10482 12486 10494 12538
rect 10494 12486 10500 12538
rect 10524 12486 10546 12538
rect 10546 12486 10558 12538
rect 10558 12486 10580 12538
rect 10604 12486 10610 12538
rect 10610 12486 10622 12538
rect 10622 12486 10660 12538
rect 10684 12486 10686 12538
rect 10686 12486 10738 12538
rect 10738 12486 10740 12538
rect 10364 12484 10420 12486
rect 10444 12484 10500 12486
rect 10524 12484 10580 12486
rect 10604 12484 10660 12486
rect 10684 12484 10740 12486
rect 11058 14048 11114 14104
rect 11242 17176 11298 17232
rect 11518 18128 11574 18184
rect 11334 16652 11390 16688
rect 11334 16632 11336 16652
rect 11336 16632 11388 16652
rect 11388 16632 11390 16652
rect 11702 16632 11758 16688
rect 10874 11872 10930 11928
rect 10364 11450 10420 11452
rect 10444 11450 10500 11452
rect 10524 11450 10580 11452
rect 10604 11450 10660 11452
rect 10684 11450 10740 11452
rect 10364 11398 10366 11450
rect 10366 11398 10418 11450
rect 10418 11398 10420 11450
rect 10444 11398 10482 11450
rect 10482 11398 10494 11450
rect 10494 11398 10500 11450
rect 10524 11398 10546 11450
rect 10546 11398 10558 11450
rect 10558 11398 10580 11450
rect 10604 11398 10610 11450
rect 10610 11398 10622 11450
rect 10622 11398 10660 11450
rect 10684 11398 10686 11450
rect 10686 11398 10738 11450
rect 10738 11398 10740 11450
rect 10364 11396 10420 11398
rect 10444 11396 10500 11398
rect 10524 11396 10580 11398
rect 10604 11396 10660 11398
rect 10684 11396 10740 11398
rect 10364 10362 10420 10364
rect 10444 10362 10500 10364
rect 10524 10362 10580 10364
rect 10604 10362 10660 10364
rect 10684 10362 10740 10364
rect 10364 10310 10366 10362
rect 10366 10310 10418 10362
rect 10418 10310 10420 10362
rect 10444 10310 10482 10362
rect 10482 10310 10494 10362
rect 10494 10310 10500 10362
rect 10524 10310 10546 10362
rect 10546 10310 10558 10362
rect 10558 10310 10580 10362
rect 10604 10310 10610 10362
rect 10610 10310 10622 10362
rect 10622 10310 10660 10362
rect 10684 10310 10686 10362
rect 10686 10310 10738 10362
rect 10738 10310 10740 10362
rect 10364 10308 10420 10310
rect 10444 10308 10500 10310
rect 10524 10308 10580 10310
rect 10604 10308 10660 10310
rect 10684 10308 10740 10310
rect 10046 9832 10102 9888
rect 11058 9696 11114 9752
rect 10322 9444 10378 9480
rect 10322 9424 10324 9444
rect 10324 9424 10376 9444
rect 10376 9424 10378 9444
rect 10874 9288 10930 9344
rect 10364 9274 10420 9276
rect 10444 9274 10500 9276
rect 10524 9274 10580 9276
rect 10604 9274 10660 9276
rect 10684 9274 10740 9276
rect 10364 9222 10366 9274
rect 10366 9222 10418 9274
rect 10418 9222 10420 9274
rect 10444 9222 10482 9274
rect 10482 9222 10494 9274
rect 10494 9222 10500 9274
rect 10524 9222 10546 9274
rect 10546 9222 10558 9274
rect 10558 9222 10580 9274
rect 10604 9222 10610 9274
rect 10610 9222 10622 9274
rect 10622 9222 10660 9274
rect 10684 9222 10686 9274
rect 10686 9222 10738 9274
rect 10738 9222 10740 9274
rect 10364 9220 10420 9222
rect 10444 9220 10500 9222
rect 10524 9220 10580 9222
rect 10604 9220 10660 9222
rect 10684 9220 10740 9222
rect 10322 8372 10324 8392
rect 10324 8372 10376 8392
rect 10376 8372 10378 8392
rect 10322 8336 10378 8372
rect 10364 8186 10420 8188
rect 10444 8186 10500 8188
rect 10524 8186 10580 8188
rect 10604 8186 10660 8188
rect 10684 8186 10740 8188
rect 10364 8134 10366 8186
rect 10366 8134 10418 8186
rect 10418 8134 10420 8186
rect 10444 8134 10482 8186
rect 10482 8134 10494 8186
rect 10494 8134 10500 8186
rect 10524 8134 10546 8186
rect 10546 8134 10558 8186
rect 10558 8134 10580 8186
rect 10604 8134 10610 8186
rect 10610 8134 10622 8186
rect 10622 8134 10660 8186
rect 10684 8134 10686 8186
rect 10686 8134 10738 8186
rect 10738 8134 10740 8186
rect 10364 8132 10420 8134
rect 10444 8132 10500 8134
rect 10524 8132 10580 8134
rect 10604 8132 10660 8134
rect 10684 8132 10740 8134
rect 10046 6024 10102 6080
rect 9954 5888 10010 5944
rect 10782 7928 10838 7984
rect 10364 7098 10420 7100
rect 10444 7098 10500 7100
rect 10524 7098 10580 7100
rect 10604 7098 10660 7100
rect 10684 7098 10740 7100
rect 10364 7046 10366 7098
rect 10366 7046 10418 7098
rect 10418 7046 10420 7098
rect 10444 7046 10482 7098
rect 10482 7046 10494 7098
rect 10494 7046 10500 7098
rect 10524 7046 10546 7098
rect 10546 7046 10558 7098
rect 10558 7046 10580 7098
rect 10604 7046 10610 7098
rect 10610 7046 10622 7098
rect 10622 7046 10660 7098
rect 10684 7046 10686 7098
rect 10686 7046 10738 7098
rect 10738 7046 10740 7098
rect 10364 7044 10420 7046
rect 10444 7044 10500 7046
rect 10524 7044 10580 7046
rect 10604 7044 10660 7046
rect 10684 7044 10740 7046
rect 10414 6860 10470 6896
rect 10414 6840 10416 6860
rect 10416 6840 10468 6860
rect 10468 6840 10470 6860
rect 10046 5480 10102 5536
rect 10138 5344 10194 5400
rect 10506 6568 10562 6624
rect 11150 9152 11206 9208
rect 10874 6296 10930 6352
rect 10364 6010 10420 6012
rect 10444 6010 10500 6012
rect 10524 6010 10580 6012
rect 10604 6010 10660 6012
rect 10684 6010 10740 6012
rect 10364 5958 10366 6010
rect 10366 5958 10418 6010
rect 10418 5958 10420 6010
rect 10444 5958 10482 6010
rect 10482 5958 10494 6010
rect 10494 5958 10500 6010
rect 10524 5958 10546 6010
rect 10546 5958 10558 6010
rect 10558 5958 10580 6010
rect 10604 5958 10610 6010
rect 10610 5958 10622 6010
rect 10622 5958 10660 6010
rect 10684 5958 10686 6010
rect 10686 5958 10738 6010
rect 10738 5958 10740 6010
rect 10364 5956 10420 5958
rect 10444 5956 10500 5958
rect 10524 5956 10580 5958
rect 10604 5956 10660 5958
rect 10684 5956 10740 5958
rect 10364 4922 10420 4924
rect 10444 4922 10500 4924
rect 10524 4922 10580 4924
rect 10604 4922 10660 4924
rect 10684 4922 10740 4924
rect 10364 4870 10366 4922
rect 10366 4870 10418 4922
rect 10418 4870 10420 4922
rect 10444 4870 10482 4922
rect 10482 4870 10494 4922
rect 10494 4870 10500 4922
rect 10524 4870 10546 4922
rect 10546 4870 10558 4922
rect 10558 4870 10580 4922
rect 10604 4870 10610 4922
rect 10610 4870 10622 4922
rect 10622 4870 10660 4922
rect 10684 4870 10686 4922
rect 10686 4870 10738 4922
rect 10738 4870 10740 4922
rect 10364 4868 10420 4870
rect 10444 4868 10500 4870
rect 10524 4868 10580 4870
rect 10604 4868 10660 4870
rect 10684 4868 10740 4870
rect 10046 3984 10102 4040
rect 10690 4020 10692 4040
rect 10692 4020 10744 4040
rect 10744 4020 10746 4040
rect 10690 3984 10746 4020
rect 10364 3834 10420 3836
rect 10444 3834 10500 3836
rect 10524 3834 10580 3836
rect 10604 3834 10660 3836
rect 10684 3834 10740 3836
rect 10364 3782 10366 3834
rect 10366 3782 10418 3834
rect 10418 3782 10420 3834
rect 10444 3782 10482 3834
rect 10482 3782 10494 3834
rect 10494 3782 10500 3834
rect 10524 3782 10546 3834
rect 10546 3782 10558 3834
rect 10558 3782 10580 3834
rect 10604 3782 10610 3834
rect 10610 3782 10622 3834
rect 10622 3782 10660 3834
rect 10684 3782 10686 3834
rect 10686 3782 10738 3834
rect 10738 3782 10740 3834
rect 10364 3780 10420 3782
rect 10444 3780 10500 3782
rect 10524 3780 10580 3782
rect 10604 3780 10660 3782
rect 10684 3780 10740 3782
rect 10506 3596 10562 3632
rect 11334 12280 11390 12336
rect 11610 15272 11666 15328
rect 11610 15136 11666 15192
rect 11518 11076 11574 11112
rect 11518 11056 11520 11076
rect 11520 11056 11572 11076
rect 11572 11056 11574 11076
rect 11610 10920 11666 10976
rect 12070 15544 12126 15600
rect 12438 15816 12494 15872
rect 12162 15000 12218 15056
rect 12070 14900 12072 14920
rect 12072 14900 12124 14920
rect 12124 14900 12126 14920
rect 12070 14864 12126 14900
rect 12070 14592 12126 14648
rect 12162 14320 12218 14376
rect 12254 13776 12310 13832
rect 11794 12300 11850 12336
rect 11794 12280 11796 12300
rect 11796 12280 11848 12300
rect 11848 12280 11850 12300
rect 11794 12008 11850 12064
rect 11794 11328 11850 11384
rect 12346 12824 12402 12880
rect 12346 12416 12402 12472
rect 12070 10920 12126 10976
rect 12714 17740 12770 17776
rect 12714 17720 12716 17740
rect 12716 17720 12768 17740
rect 12768 17720 12770 17740
rect 12806 16632 12862 16688
rect 13364 19610 13420 19612
rect 13444 19610 13500 19612
rect 13524 19610 13580 19612
rect 13604 19610 13660 19612
rect 13684 19610 13740 19612
rect 13364 19558 13366 19610
rect 13366 19558 13418 19610
rect 13418 19558 13420 19610
rect 13444 19558 13482 19610
rect 13482 19558 13494 19610
rect 13494 19558 13500 19610
rect 13524 19558 13546 19610
rect 13546 19558 13558 19610
rect 13558 19558 13580 19610
rect 13604 19558 13610 19610
rect 13610 19558 13622 19610
rect 13622 19558 13660 19610
rect 13684 19558 13686 19610
rect 13686 19558 13738 19610
rect 13738 19558 13740 19610
rect 13364 19556 13420 19558
rect 13444 19556 13500 19558
rect 13524 19556 13580 19558
rect 13604 19556 13660 19558
rect 13684 19556 13740 19558
rect 13266 18672 13322 18728
rect 13364 18522 13420 18524
rect 13444 18522 13500 18524
rect 13524 18522 13580 18524
rect 13604 18522 13660 18524
rect 13684 18522 13740 18524
rect 13364 18470 13366 18522
rect 13366 18470 13418 18522
rect 13418 18470 13420 18522
rect 13444 18470 13482 18522
rect 13482 18470 13494 18522
rect 13494 18470 13500 18522
rect 13524 18470 13546 18522
rect 13546 18470 13558 18522
rect 13558 18470 13580 18522
rect 13604 18470 13610 18522
rect 13610 18470 13622 18522
rect 13622 18470 13660 18522
rect 13684 18470 13686 18522
rect 13686 18470 13738 18522
rect 13738 18470 13740 18522
rect 13364 18468 13420 18470
rect 13444 18468 13500 18470
rect 13524 18468 13580 18470
rect 13604 18468 13660 18470
rect 13684 18468 13740 18470
rect 14370 18028 14372 18048
rect 14372 18028 14424 18048
rect 14424 18028 14426 18048
rect 14370 17992 14426 18028
rect 13364 17434 13420 17436
rect 13444 17434 13500 17436
rect 13524 17434 13580 17436
rect 13604 17434 13660 17436
rect 13684 17434 13740 17436
rect 13364 17382 13366 17434
rect 13366 17382 13418 17434
rect 13418 17382 13420 17434
rect 13444 17382 13482 17434
rect 13482 17382 13494 17434
rect 13494 17382 13500 17434
rect 13524 17382 13546 17434
rect 13546 17382 13558 17434
rect 13558 17382 13580 17434
rect 13604 17382 13610 17434
rect 13610 17382 13622 17434
rect 13622 17382 13660 17434
rect 13684 17382 13686 17434
rect 13686 17382 13738 17434
rect 13738 17382 13740 17434
rect 13364 17380 13420 17382
rect 13444 17380 13500 17382
rect 13524 17380 13580 17382
rect 13604 17380 13660 17382
rect 13684 17380 13740 17382
rect 13082 16632 13138 16688
rect 12898 15136 12954 15192
rect 12714 14592 12770 14648
rect 12622 14320 12678 14376
rect 12714 13504 12770 13560
rect 12806 13368 12862 13424
rect 12622 13096 12678 13152
rect 12622 12860 12624 12880
rect 12624 12860 12676 12880
rect 12676 12860 12678 12880
rect 12622 12824 12678 12860
rect 12622 11872 12678 11928
rect 11518 9152 11574 9208
rect 11702 9152 11758 9208
rect 11610 8336 11666 8392
rect 11702 6996 11758 7032
rect 11702 6976 11704 6996
rect 11704 6976 11756 6996
rect 11756 6976 11758 6996
rect 11702 6568 11758 6624
rect 11334 5208 11390 5264
rect 11334 4664 11390 4720
rect 10506 3576 10508 3596
rect 10508 3576 10560 3596
rect 10560 3576 10562 3596
rect 8298 2372 8354 2408
rect 8298 2352 8300 2372
rect 8300 2352 8352 2372
rect 8352 2352 8354 2372
rect 10230 3440 10286 3496
rect 10598 3304 10654 3360
rect 11334 3032 11390 3088
rect 11518 3304 11574 3360
rect 10966 2760 11022 2816
rect 10364 2746 10420 2748
rect 10444 2746 10500 2748
rect 10524 2746 10580 2748
rect 10604 2746 10660 2748
rect 10684 2746 10740 2748
rect 10364 2694 10366 2746
rect 10366 2694 10418 2746
rect 10418 2694 10420 2746
rect 10444 2694 10482 2746
rect 10482 2694 10494 2746
rect 10494 2694 10500 2746
rect 10524 2694 10546 2746
rect 10546 2694 10558 2746
rect 10558 2694 10580 2746
rect 10604 2694 10610 2746
rect 10610 2694 10622 2746
rect 10622 2694 10660 2746
rect 10684 2694 10686 2746
rect 10686 2694 10738 2746
rect 10738 2694 10740 2746
rect 10364 2692 10420 2694
rect 10444 2692 10500 2694
rect 10524 2692 10580 2694
rect 10604 2692 10660 2694
rect 10684 2692 10740 2694
rect 10230 2352 10286 2408
rect 8942 1420 8998 1456
rect 8942 1400 8944 1420
rect 8944 1400 8996 1420
rect 8996 1400 8998 1420
rect 9678 2216 9734 2272
rect 9954 2080 10010 2136
rect 9862 1944 9918 2000
rect 10046 1808 10102 1864
rect 11334 2644 11390 2680
rect 11610 2760 11666 2816
rect 12254 10548 12256 10568
rect 12256 10548 12308 10568
rect 12308 10548 12310 10568
rect 12254 10512 12310 10548
rect 12622 11600 12678 11656
rect 12530 11464 12586 11520
rect 13364 16346 13420 16348
rect 13444 16346 13500 16348
rect 13524 16346 13580 16348
rect 13604 16346 13660 16348
rect 13684 16346 13740 16348
rect 13364 16294 13366 16346
rect 13366 16294 13418 16346
rect 13418 16294 13420 16346
rect 13444 16294 13482 16346
rect 13482 16294 13494 16346
rect 13494 16294 13500 16346
rect 13524 16294 13546 16346
rect 13546 16294 13558 16346
rect 13558 16294 13580 16346
rect 13604 16294 13610 16346
rect 13610 16294 13622 16346
rect 13622 16294 13660 16346
rect 13684 16294 13686 16346
rect 13686 16294 13738 16346
rect 13738 16294 13740 16346
rect 13364 16292 13420 16294
rect 13444 16292 13500 16294
rect 13524 16292 13580 16294
rect 13604 16292 13660 16294
rect 13684 16292 13740 16294
rect 13364 15258 13420 15260
rect 13444 15258 13500 15260
rect 13524 15258 13580 15260
rect 13604 15258 13660 15260
rect 13684 15258 13740 15260
rect 13364 15206 13366 15258
rect 13366 15206 13418 15258
rect 13418 15206 13420 15258
rect 13444 15206 13482 15258
rect 13482 15206 13494 15258
rect 13494 15206 13500 15258
rect 13524 15206 13546 15258
rect 13546 15206 13558 15258
rect 13558 15206 13580 15258
rect 13604 15206 13610 15258
rect 13610 15206 13622 15258
rect 13622 15206 13660 15258
rect 13684 15206 13686 15258
rect 13686 15206 13738 15258
rect 13738 15206 13740 15258
rect 13364 15204 13420 15206
rect 13444 15204 13500 15206
rect 13524 15204 13580 15206
rect 13604 15204 13660 15206
rect 13684 15204 13740 15206
rect 13364 14170 13420 14172
rect 13444 14170 13500 14172
rect 13524 14170 13580 14172
rect 13604 14170 13660 14172
rect 13684 14170 13740 14172
rect 13364 14118 13366 14170
rect 13366 14118 13418 14170
rect 13418 14118 13420 14170
rect 13444 14118 13482 14170
rect 13482 14118 13494 14170
rect 13494 14118 13500 14170
rect 13524 14118 13546 14170
rect 13546 14118 13558 14170
rect 13558 14118 13580 14170
rect 13604 14118 13610 14170
rect 13610 14118 13622 14170
rect 13622 14118 13660 14170
rect 13684 14118 13686 14170
rect 13686 14118 13738 14170
rect 13738 14118 13740 14170
rect 13364 14116 13420 14118
rect 13444 14116 13500 14118
rect 13524 14116 13580 14118
rect 13604 14116 13660 14118
rect 13684 14116 13740 14118
rect 13266 13812 13268 13832
rect 13268 13812 13320 13832
rect 13320 13812 13322 13832
rect 13266 13776 13322 13812
rect 14094 14456 14150 14512
rect 13364 13082 13420 13084
rect 13444 13082 13500 13084
rect 13524 13082 13580 13084
rect 13604 13082 13660 13084
rect 13684 13082 13740 13084
rect 13364 13030 13366 13082
rect 13366 13030 13418 13082
rect 13418 13030 13420 13082
rect 13444 13030 13482 13082
rect 13482 13030 13494 13082
rect 13494 13030 13500 13082
rect 13524 13030 13546 13082
rect 13546 13030 13558 13082
rect 13558 13030 13580 13082
rect 13604 13030 13610 13082
rect 13610 13030 13622 13082
rect 13622 13030 13660 13082
rect 13684 13030 13686 13082
rect 13686 13030 13738 13082
rect 13738 13030 13740 13082
rect 13364 13028 13420 13030
rect 13444 13028 13500 13030
rect 13524 13028 13580 13030
rect 13604 13028 13660 13030
rect 13684 13028 13740 13030
rect 13910 12824 13966 12880
rect 13174 11736 13230 11792
rect 13364 11994 13420 11996
rect 13444 11994 13500 11996
rect 13524 11994 13580 11996
rect 13604 11994 13660 11996
rect 13684 11994 13740 11996
rect 13364 11942 13366 11994
rect 13366 11942 13418 11994
rect 13418 11942 13420 11994
rect 13444 11942 13482 11994
rect 13482 11942 13494 11994
rect 13494 11942 13500 11994
rect 13524 11942 13546 11994
rect 13546 11942 13558 11994
rect 13558 11942 13580 11994
rect 13604 11942 13610 11994
rect 13610 11942 13622 11994
rect 13622 11942 13660 11994
rect 13684 11942 13686 11994
rect 13686 11942 13738 11994
rect 13738 11942 13740 11994
rect 13364 11940 13420 11942
rect 13444 11940 13500 11942
rect 13524 11940 13580 11942
rect 13604 11940 13660 11942
rect 13684 11940 13740 11942
rect 13542 11600 13598 11656
rect 12714 11192 12770 11248
rect 12806 11056 12862 11112
rect 12806 10956 12808 10976
rect 12808 10956 12860 10976
rect 12860 10956 12862 10976
rect 12806 10920 12862 10956
rect 12254 10376 12310 10432
rect 12530 9696 12586 9752
rect 12530 9424 12586 9480
rect 13174 11212 13230 11248
rect 13174 11192 13176 11212
rect 13176 11192 13228 11212
rect 13228 11192 13230 11212
rect 13082 11056 13138 11112
rect 13082 10784 13138 10840
rect 12806 9152 12862 9208
rect 12714 8064 12770 8120
rect 12346 5072 12402 5128
rect 12254 4972 12256 4992
rect 12256 4972 12308 4992
rect 12308 4972 12310 4992
rect 12254 4936 12310 4972
rect 12254 4820 12310 4856
rect 12254 4800 12256 4820
rect 12256 4800 12308 4820
rect 12308 4800 12310 4820
rect 12622 4936 12678 4992
rect 12990 6024 13046 6080
rect 12898 5244 12900 5264
rect 12900 5244 12952 5264
rect 12952 5244 12954 5264
rect 12898 5208 12954 5244
rect 12898 4664 12954 4720
rect 13364 10906 13420 10908
rect 13444 10906 13500 10908
rect 13524 10906 13580 10908
rect 13604 10906 13660 10908
rect 13684 10906 13740 10908
rect 13364 10854 13366 10906
rect 13366 10854 13418 10906
rect 13418 10854 13420 10906
rect 13444 10854 13482 10906
rect 13482 10854 13494 10906
rect 13494 10854 13500 10906
rect 13524 10854 13546 10906
rect 13546 10854 13558 10906
rect 13558 10854 13580 10906
rect 13604 10854 13610 10906
rect 13610 10854 13622 10906
rect 13622 10854 13660 10906
rect 13684 10854 13686 10906
rect 13686 10854 13738 10906
rect 13738 10854 13740 10906
rect 13364 10852 13420 10854
rect 13444 10852 13500 10854
rect 13524 10852 13580 10854
rect 13604 10852 13660 10854
rect 13684 10852 13740 10854
rect 14738 16904 14794 16960
rect 14554 14220 14556 14240
rect 14556 14220 14608 14240
rect 14608 14220 14610 14240
rect 14554 14184 14610 14220
rect 14186 11872 14242 11928
rect 14186 11636 14188 11656
rect 14188 11636 14240 11656
rect 14240 11636 14242 11656
rect 14186 11600 14242 11636
rect 14370 11600 14426 11656
rect 14278 11192 14334 11248
rect 14186 11056 14242 11112
rect 13450 10512 13506 10568
rect 13634 10240 13690 10296
rect 13364 9818 13420 9820
rect 13444 9818 13500 9820
rect 13524 9818 13580 9820
rect 13604 9818 13660 9820
rect 13684 9818 13740 9820
rect 13364 9766 13366 9818
rect 13366 9766 13418 9818
rect 13418 9766 13420 9818
rect 13444 9766 13482 9818
rect 13482 9766 13494 9818
rect 13494 9766 13500 9818
rect 13524 9766 13546 9818
rect 13546 9766 13558 9818
rect 13558 9766 13580 9818
rect 13604 9766 13610 9818
rect 13610 9766 13622 9818
rect 13622 9766 13660 9818
rect 13684 9766 13686 9818
rect 13686 9766 13738 9818
rect 13738 9766 13740 9818
rect 13364 9764 13420 9766
rect 13444 9764 13500 9766
rect 13524 9764 13580 9766
rect 13604 9764 13660 9766
rect 13684 9764 13740 9766
rect 13818 9152 13874 9208
rect 13364 8730 13420 8732
rect 13444 8730 13500 8732
rect 13524 8730 13580 8732
rect 13604 8730 13660 8732
rect 13684 8730 13740 8732
rect 13364 8678 13366 8730
rect 13366 8678 13418 8730
rect 13418 8678 13420 8730
rect 13444 8678 13482 8730
rect 13482 8678 13494 8730
rect 13494 8678 13500 8730
rect 13524 8678 13546 8730
rect 13546 8678 13558 8730
rect 13558 8678 13580 8730
rect 13604 8678 13610 8730
rect 13610 8678 13622 8730
rect 13622 8678 13660 8730
rect 13684 8678 13686 8730
rect 13686 8678 13738 8730
rect 13738 8678 13740 8730
rect 13364 8676 13420 8678
rect 13444 8676 13500 8678
rect 13524 8676 13580 8678
rect 13604 8676 13660 8678
rect 13684 8676 13740 8678
rect 13364 7642 13420 7644
rect 13444 7642 13500 7644
rect 13524 7642 13580 7644
rect 13604 7642 13660 7644
rect 13684 7642 13740 7644
rect 13364 7590 13366 7642
rect 13366 7590 13418 7642
rect 13418 7590 13420 7642
rect 13444 7590 13482 7642
rect 13482 7590 13494 7642
rect 13494 7590 13500 7642
rect 13524 7590 13546 7642
rect 13546 7590 13558 7642
rect 13558 7590 13580 7642
rect 13604 7590 13610 7642
rect 13610 7590 13622 7642
rect 13622 7590 13660 7642
rect 13684 7590 13686 7642
rect 13686 7590 13738 7642
rect 13738 7590 13740 7642
rect 13364 7588 13420 7590
rect 13444 7588 13500 7590
rect 13524 7588 13580 7590
rect 13604 7588 13660 7590
rect 13684 7588 13740 7590
rect 13634 7284 13636 7304
rect 13636 7284 13688 7304
rect 13688 7284 13690 7304
rect 13634 7248 13690 7284
rect 13910 7248 13966 7304
rect 13910 6740 13912 6760
rect 13912 6740 13964 6760
rect 13964 6740 13966 6760
rect 13910 6704 13966 6740
rect 13364 6554 13420 6556
rect 13444 6554 13500 6556
rect 13524 6554 13580 6556
rect 13604 6554 13660 6556
rect 13684 6554 13740 6556
rect 13364 6502 13366 6554
rect 13366 6502 13418 6554
rect 13418 6502 13420 6554
rect 13444 6502 13482 6554
rect 13482 6502 13494 6554
rect 13494 6502 13500 6554
rect 13524 6502 13546 6554
rect 13546 6502 13558 6554
rect 13558 6502 13580 6554
rect 13604 6502 13610 6554
rect 13610 6502 13622 6554
rect 13622 6502 13660 6554
rect 13684 6502 13686 6554
rect 13686 6502 13738 6554
rect 13738 6502 13740 6554
rect 13364 6500 13420 6502
rect 13444 6500 13500 6502
rect 13524 6500 13580 6502
rect 13604 6500 13660 6502
rect 13684 6500 13740 6502
rect 14278 9968 14334 10024
rect 13364 5466 13420 5468
rect 13444 5466 13500 5468
rect 13524 5466 13580 5468
rect 13604 5466 13660 5468
rect 13684 5466 13740 5468
rect 13364 5414 13366 5466
rect 13366 5414 13418 5466
rect 13418 5414 13420 5466
rect 13444 5414 13482 5466
rect 13482 5414 13494 5466
rect 13494 5414 13500 5466
rect 13524 5414 13546 5466
rect 13546 5414 13558 5466
rect 13558 5414 13580 5466
rect 13604 5414 13610 5466
rect 13610 5414 13622 5466
rect 13622 5414 13660 5466
rect 13684 5414 13686 5466
rect 13686 5414 13738 5466
rect 13738 5414 13740 5466
rect 13364 5412 13420 5414
rect 13444 5412 13500 5414
rect 13524 5412 13580 5414
rect 13604 5412 13660 5414
rect 13684 5412 13740 5414
rect 12898 4564 12900 4584
rect 12900 4564 12952 4584
rect 12952 4564 12954 4584
rect 12898 4528 12954 4564
rect 11334 2624 11336 2644
rect 11336 2624 11388 2644
rect 11388 2624 11390 2644
rect 10966 2352 11022 2408
rect 10364 1658 10420 1660
rect 10444 1658 10500 1660
rect 10524 1658 10580 1660
rect 10604 1658 10660 1660
rect 10684 1658 10740 1660
rect 10364 1606 10366 1658
rect 10366 1606 10418 1658
rect 10418 1606 10420 1658
rect 10444 1606 10482 1658
rect 10482 1606 10494 1658
rect 10494 1606 10500 1658
rect 10524 1606 10546 1658
rect 10546 1606 10558 1658
rect 10558 1606 10580 1658
rect 10604 1606 10610 1658
rect 10610 1606 10622 1658
rect 10622 1606 10660 1658
rect 10684 1606 10686 1658
rect 10686 1606 10738 1658
rect 10738 1606 10740 1658
rect 10364 1604 10420 1606
rect 10444 1604 10500 1606
rect 10524 1604 10580 1606
rect 10604 1604 10660 1606
rect 10684 1604 10740 1606
rect 9862 1284 9918 1320
rect 9862 1264 9864 1284
rect 9864 1264 9916 1284
rect 9916 1264 9918 1284
rect 10966 1400 11022 1456
rect 10364 570 10420 572
rect 10444 570 10500 572
rect 10524 570 10580 572
rect 10604 570 10660 572
rect 10684 570 10740 572
rect 10364 518 10366 570
rect 10366 518 10418 570
rect 10418 518 10420 570
rect 10444 518 10482 570
rect 10482 518 10494 570
rect 10494 518 10500 570
rect 10524 518 10546 570
rect 10546 518 10558 570
rect 10558 518 10580 570
rect 10604 518 10610 570
rect 10610 518 10622 570
rect 10622 518 10660 570
rect 10684 518 10686 570
rect 10686 518 10738 570
rect 10738 518 10740 570
rect 10364 516 10420 518
rect 10444 516 10500 518
rect 10524 516 10580 518
rect 10604 516 10660 518
rect 10684 516 10740 518
rect 11242 2388 11244 2408
rect 11244 2388 11296 2408
rect 11296 2388 11298 2408
rect 11242 2352 11298 2388
rect 11886 2644 11942 2680
rect 11886 2624 11888 2644
rect 11888 2624 11940 2644
rect 11940 2624 11942 2644
rect 11886 2216 11942 2272
rect 12162 2080 12218 2136
rect 12438 2524 12440 2544
rect 12440 2524 12492 2544
rect 12492 2524 12494 2544
rect 12438 2488 12494 2524
rect 12622 2796 12624 2816
rect 12624 2796 12676 2816
rect 12676 2796 12678 2816
rect 12622 2760 12678 2796
rect 12438 2216 12494 2272
rect 12438 1808 12494 1864
rect 12070 1536 12126 1592
rect 12622 1808 12678 1864
rect 10046 176 10102 232
rect 12070 76 12072 96
rect 12072 76 12124 96
rect 12124 76 12126 96
rect 12070 40 12126 76
rect 12806 1808 12862 1864
rect 13364 4378 13420 4380
rect 13444 4378 13500 4380
rect 13524 4378 13580 4380
rect 13604 4378 13660 4380
rect 13684 4378 13740 4380
rect 13364 4326 13366 4378
rect 13366 4326 13418 4378
rect 13418 4326 13420 4378
rect 13444 4326 13482 4378
rect 13482 4326 13494 4378
rect 13494 4326 13500 4378
rect 13524 4326 13546 4378
rect 13546 4326 13558 4378
rect 13558 4326 13580 4378
rect 13604 4326 13610 4378
rect 13610 4326 13622 4378
rect 13622 4326 13660 4378
rect 13684 4326 13686 4378
rect 13686 4326 13738 4378
rect 13738 4326 13740 4378
rect 13364 4324 13420 4326
rect 13444 4324 13500 4326
rect 13524 4324 13580 4326
rect 13604 4324 13660 4326
rect 13684 4324 13740 4326
rect 15106 20848 15162 20904
rect 16364 22330 16420 22332
rect 16444 22330 16500 22332
rect 16524 22330 16580 22332
rect 16604 22330 16660 22332
rect 16684 22330 16740 22332
rect 16364 22278 16366 22330
rect 16366 22278 16418 22330
rect 16418 22278 16420 22330
rect 16444 22278 16482 22330
rect 16482 22278 16494 22330
rect 16494 22278 16500 22330
rect 16524 22278 16546 22330
rect 16546 22278 16558 22330
rect 16558 22278 16580 22330
rect 16604 22278 16610 22330
rect 16610 22278 16622 22330
rect 16622 22278 16660 22330
rect 16684 22278 16686 22330
rect 16686 22278 16738 22330
rect 16738 22278 16740 22330
rect 16364 22276 16420 22278
rect 16444 22276 16500 22278
rect 16524 22276 16580 22278
rect 16604 22276 16660 22278
rect 16684 22276 16740 22278
rect 16118 21664 16174 21720
rect 15934 21528 15990 21584
rect 16364 21242 16420 21244
rect 16444 21242 16500 21244
rect 16524 21242 16580 21244
rect 16604 21242 16660 21244
rect 16684 21242 16740 21244
rect 16364 21190 16366 21242
rect 16366 21190 16418 21242
rect 16418 21190 16420 21242
rect 16444 21190 16482 21242
rect 16482 21190 16494 21242
rect 16494 21190 16500 21242
rect 16524 21190 16546 21242
rect 16546 21190 16558 21242
rect 16558 21190 16580 21242
rect 16604 21190 16610 21242
rect 16610 21190 16622 21242
rect 16622 21190 16660 21242
rect 16684 21190 16686 21242
rect 16686 21190 16738 21242
rect 16738 21190 16740 21242
rect 16364 21188 16420 21190
rect 16444 21188 16500 21190
rect 16524 21188 16580 21190
rect 16604 21188 16660 21190
rect 16684 21188 16740 21190
rect 16210 20460 16266 20496
rect 16210 20440 16212 20460
rect 16212 20440 16264 20460
rect 16264 20440 16266 20460
rect 16364 20154 16420 20156
rect 16444 20154 16500 20156
rect 16524 20154 16580 20156
rect 16604 20154 16660 20156
rect 16684 20154 16740 20156
rect 16364 20102 16366 20154
rect 16366 20102 16418 20154
rect 16418 20102 16420 20154
rect 16444 20102 16482 20154
rect 16482 20102 16494 20154
rect 16494 20102 16500 20154
rect 16524 20102 16546 20154
rect 16546 20102 16558 20154
rect 16558 20102 16580 20154
rect 16604 20102 16610 20154
rect 16610 20102 16622 20154
rect 16622 20102 16660 20154
rect 16684 20102 16686 20154
rect 16686 20102 16738 20154
rect 16738 20102 16740 20154
rect 16364 20100 16420 20102
rect 16444 20100 16500 20102
rect 16524 20100 16580 20102
rect 16604 20100 16660 20102
rect 16684 20100 16740 20102
rect 16854 20340 16856 20360
rect 16856 20340 16908 20360
rect 16908 20340 16910 20360
rect 16854 20304 16910 20340
rect 17222 20576 17278 20632
rect 16302 19352 16358 19408
rect 16364 19066 16420 19068
rect 16444 19066 16500 19068
rect 16524 19066 16580 19068
rect 16604 19066 16660 19068
rect 16684 19066 16740 19068
rect 16364 19014 16366 19066
rect 16366 19014 16418 19066
rect 16418 19014 16420 19066
rect 16444 19014 16482 19066
rect 16482 19014 16494 19066
rect 16494 19014 16500 19066
rect 16524 19014 16546 19066
rect 16546 19014 16558 19066
rect 16558 19014 16580 19066
rect 16604 19014 16610 19066
rect 16610 19014 16622 19066
rect 16622 19014 16660 19066
rect 16684 19014 16686 19066
rect 16686 19014 16738 19066
rect 16738 19014 16740 19066
rect 16364 19012 16420 19014
rect 16444 19012 16500 19014
rect 16524 19012 16580 19014
rect 16604 19012 16660 19014
rect 16684 19012 16740 19014
rect 16364 17978 16420 17980
rect 16444 17978 16500 17980
rect 16524 17978 16580 17980
rect 16604 17978 16660 17980
rect 16684 17978 16740 17980
rect 16364 17926 16366 17978
rect 16366 17926 16418 17978
rect 16418 17926 16420 17978
rect 16444 17926 16482 17978
rect 16482 17926 16494 17978
rect 16494 17926 16500 17978
rect 16524 17926 16546 17978
rect 16546 17926 16558 17978
rect 16558 17926 16580 17978
rect 16604 17926 16610 17978
rect 16610 17926 16622 17978
rect 16622 17926 16660 17978
rect 16684 17926 16686 17978
rect 16686 17926 16738 17978
rect 16738 17926 16740 17978
rect 16364 17924 16420 17926
rect 16444 17924 16500 17926
rect 16524 17924 16580 17926
rect 16604 17924 16660 17926
rect 16684 17924 16740 17926
rect 15842 17740 15898 17776
rect 15842 17720 15844 17740
rect 15844 17720 15896 17740
rect 15896 17720 15898 17740
rect 15750 16904 15806 16960
rect 15658 15816 15714 15872
rect 15198 14320 15254 14376
rect 15842 13912 15898 13968
rect 15750 13640 15806 13696
rect 15474 12416 15530 12472
rect 15382 12008 15438 12064
rect 15382 11212 15438 11248
rect 15382 11192 15384 11212
rect 15384 11192 15436 11212
rect 15436 11192 15438 11212
rect 14830 10512 14886 10568
rect 14646 10376 14702 10432
rect 14830 9832 14886 9888
rect 14462 9016 14518 9072
rect 14554 7692 14556 7712
rect 14556 7692 14608 7712
rect 14608 7692 14610 7712
rect 14554 7656 14610 7692
rect 15106 9288 15162 9344
rect 15106 9036 15162 9072
rect 15106 9016 15108 9036
rect 15108 9016 15160 9036
rect 15160 9016 15162 9036
rect 14922 8472 14978 8528
rect 15106 8780 15108 8800
rect 15108 8780 15160 8800
rect 15160 8780 15162 8800
rect 15106 8744 15162 8780
rect 15106 8472 15162 8528
rect 14186 4276 14242 4312
rect 14186 4256 14188 4276
rect 14188 4256 14240 4276
rect 14240 4256 14242 4276
rect 14094 3596 14150 3632
rect 14094 3576 14096 3596
rect 14096 3576 14148 3596
rect 14148 3576 14150 3596
rect 13364 3290 13420 3292
rect 13444 3290 13500 3292
rect 13524 3290 13580 3292
rect 13604 3290 13660 3292
rect 13684 3290 13740 3292
rect 13364 3238 13366 3290
rect 13366 3238 13418 3290
rect 13418 3238 13420 3290
rect 13444 3238 13482 3290
rect 13482 3238 13494 3290
rect 13494 3238 13500 3290
rect 13524 3238 13546 3290
rect 13546 3238 13558 3290
rect 13558 3238 13580 3290
rect 13604 3238 13610 3290
rect 13610 3238 13622 3290
rect 13622 3238 13660 3290
rect 13684 3238 13686 3290
rect 13686 3238 13738 3290
rect 13738 3238 13740 3290
rect 13364 3236 13420 3238
rect 13444 3236 13500 3238
rect 13524 3236 13580 3238
rect 13604 3236 13660 3238
rect 13684 3236 13740 3238
rect 13726 2760 13782 2816
rect 14094 2932 14096 2952
rect 14096 2932 14148 2952
rect 14148 2932 14150 2952
rect 14094 2896 14150 2932
rect 13082 2080 13138 2136
rect 15290 9696 15346 9752
rect 15290 9152 15346 9208
rect 15474 8336 15530 8392
rect 17314 19760 17370 19816
rect 16364 16890 16420 16892
rect 16444 16890 16500 16892
rect 16524 16890 16580 16892
rect 16604 16890 16660 16892
rect 16684 16890 16740 16892
rect 16364 16838 16366 16890
rect 16366 16838 16418 16890
rect 16418 16838 16420 16890
rect 16444 16838 16482 16890
rect 16482 16838 16494 16890
rect 16494 16838 16500 16890
rect 16524 16838 16546 16890
rect 16546 16838 16558 16890
rect 16558 16838 16580 16890
rect 16604 16838 16610 16890
rect 16610 16838 16622 16890
rect 16622 16838 16660 16890
rect 16684 16838 16686 16890
rect 16686 16838 16738 16890
rect 16738 16838 16740 16890
rect 16364 16836 16420 16838
rect 16444 16836 16500 16838
rect 16524 16836 16580 16838
rect 16604 16836 16660 16838
rect 16684 16836 16740 16838
rect 16026 15680 16082 15736
rect 16364 15802 16420 15804
rect 16444 15802 16500 15804
rect 16524 15802 16580 15804
rect 16604 15802 16660 15804
rect 16684 15802 16740 15804
rect 16364 15750 16366 15802
rect 16366 15750 16418 15802
rect 16418 15750 16420 15802
rect 16444 15750 16482 15802
rect 16482 15750 16494 15802
rect 16494 15750 16500 15802
rect 16524 15750 16546 15802
rect 16546 15750 16558 15802
rect 16558 15750 16580 15802
rect 16604 15750 16610 15802
rect 16610 15750 16622 15802
rect 16622 15750 16660 15802
rect 16684 15750 16686 15802
rect 16686 15750 16738 15802
rect 16738 15750 16740 15802
rect 16364 15748 16420 15750
rect 16444 15748 16500 15750
rect 16524 15748 16580 15750
rect 16604 15748 16660 15750
rect 16684 15748 16740 15750
rect 15934 9696 15990 9752
rect 15658 8608 15714 8664
rect 15566 7520 15622 7576
rect 15566 7112 15622 7168
rect 15382 6976 15438 7032
rect 15198 6024 15254 6080
rect 14922 4800 14978 4856
rect 15382 6024 15438 6080
rect 16364 14714 16420 14716
rect 16444 14714 16500 14716
rect 16524 14714 16580 14716
rect 16604 14714 16660 14716
rect 16684 14714 16740 14716
rect 16364 14662 16366 14714
rect 16366 14662 16418 14714
rect 16418 14662 16420 14714
rect 16444 14662 16482 14714
rect 16482 14662 16494 14714
rect 16494 14662 16500 14714
rect 16524 14662 16546 14714
rect 16546 14662 16558 14714
rect 16558 14662 16580 14714
rect 16604 14662 16610 14714
rect 16610 14662 16622 14714
rect 16622 14662 16660 14714
rect 16684 14662 16686 14714
rect 16686 14662 16738 14714
rect 16738 14662 16740 14714
rect 16364 14660 16420 14662
rect 16444 14660 16500 14662
rect 16524 14660 16580 14662
rect 16604 14660 16660 14662
rect 16684 14660 16740 14662
rect 16364 13626 16420 13628
rect 16444 13626 16500 13628
rect 16524 13626 16580 13628
rect 16604 13626 16660 13628
rect 16684 13626 16740 13628
rect 16364 13574 16366 13626
rect 16366 13574 16418 13626
rect 16418 13574 16420 13626
rect 16444 13574 16482 13626
rect 16482 13574 16494 13626
rect 16494 13574 16500 13626
rect 16524 13574 16546 13626
rect 16546 13574 16558 13626
rect 16558 13574 16580 13626
rect 16604 13574 16610 13626
rect 16610 13574 16622 13626
rect 16622 13574 16660 13626
rect 16684 13574 16686 13626
rect 16686 13574 16738 13626
rect 16738 13574 16740 13626
rect 16364 13572 16420 13574
rect 16444 13572 16500 13574
rect 16524 13572 16580 13574
rect 16604 13572 16660 13574
rect 16684 13572 16740 13574
rect 16364 12538 16420 12540
rect 16444 12538 16500 12540
rect 16524 12538 16580 12540
rect 16604 12538 16660 12540
rect 16684 12538 16740 12540
rect 16364 12486 16366 12538
rect 16366 12486 16418 12538
rect 16418 12486 16420 12538
rect 16444 12486 16482 12538
rect 16482 12486 16494 12538
rect 16494 12486 16500 12538
rect 16524 12486 16546 12538
rect 16546 12486 16558 12538
rect 16558 12486 16580 12538
rect 16604 12486 16610 12538
rect 16610 12486 16622 12538
rect 16622 12486 16660 12538
rect 16684 12486 16686 12538
rect 16686 12486 16738 12538
rect 16738 12486 16740 12538
rect 16364 12484 16420 12486
rect 16444 12484 16500 12486
rect 16524 12484 16580 12486
rect 16604 12484 16660 12486
rect 16684 12484 16740 12486
rect 16670 12144 16726 12200
rect 16578 11636 16580 11656
rect 16580 11636 16632 11656
rect 16632 11636 16634 11656
rect 16578 11600 16634 11636
rect 16364 11450 16420 11452
rect 16444 11450 16500 11452
rect 16524 11450 16580 11452
rect 16604 11450 16660 11452
rect 16684 11450 16740 11452
rect 16364 11398 16366 11450
rect 16366 11398 16418 11450
rect 16418 11398 16420 11450
rect 16444 11398 16482 11450
rect 16482 11398 16494 11450
rect 16494 11398 16500 11450
rect 16524 11398 16546 11450
rect 16546 11398 16558 11450
rect 16558 11398 16580 11450
rect 16604 11398 16610 11450
rect 16610 11398 16622 11450
rect 16622 11398 16660 11450
rect 16684 11398 16686 11450
rect 16686 11398 16738 11450
rect 16738 11398 16740 11450
rect 16364 11396 16420 11398
rect 16444 11396 16500 11398
rect 16524 11396 16580 11398
rect 16604 11396 16660 11398
rect 16684 11396 16740 11398
rect 16302 11212 16358 11248
rect 16302 11192 16304 11212
rect 16304 11192 16356 11212
rect 16356 11192 16358 11212
rect 16118 10124 16174 10160
rect 16118 10104 16120 10124
rect 16120 10104 16172 10124
rect 16172 10104 16174 10124
rect 16026 8064 16082 8120
rect 15750 4120 15806 4176
rect 14186 2352 14242 2408
rect 13364 2202 13420 2204
rect 13444 2202 13500 2204
rect 13524 2202 13580 2204
rect 13604 2202 13660 2204
rect 13684 2202 13740 2204
rect 13364 2150 13366 2202
rect 13366 2150 13418 2202
rect 13418 2150 13420 2202
rect 13444 2150 13482 2202
rect 13482 2150 13494 2202
rect 13494 2150 13500 2202
rect 13524 2150 13546 2202
rect 13546 2150 13558 2202
rect 13558 2150 13580 2202
rect 13604 2150 13610 2202
rect 13610 2150 13622 2202
rect 13622 2150 13660 2202
rect 13684 2150 13686 2202
rect 13686 2150 13738 2202
rect 13738 2150 13740 2202
rect 13364 2148 13420 2150
rect 13444 2148 13500 2150
rect 13524 2148 13580 2150
rect 13604 2148 13660 2150
rect 13684 2148 13740 2150
rect 13818 2080 13874 2136
rect 14278 2216 14334 2272
rect 13358 1400 13414 1456
rect 13364 1114 13420 1116
rect 13444 1114 13500 1116
rect 13524 1114 13580 1116
rect 13604 1114 13660 1116
rect 13684 1114 13740 1116
rect 13364 1062 13366 1114
rect 13366 1062 13418 1114
rect 13418 1062 13420 1114
rect 13444 1062 13482 1114
rect 13482 1062 13494 1114
rect 13494 1062 13500 1114
rect 13524 1062 13546 1114
rect 13546 1062 13558 1114
rect 13558 1062 13580 1114
rect 13604 1062 13610 1114
rect 13610 1062 13622 1114
rect 13622 1062 13660 1114
rect 13684 1062 13686 1114
rect 13686 1062 13738 1114
rect 13738 1062 13740 1114
rect 13364 1060 13420 1062
rect 13444 1060 13500 1062
rect 13524 1060 13580 1062
rect 13604 1060 13660 1062
rect 13684 1060 13740 1062
rect 14186 1012 14242 1048
rect 14186 992 14188 1012
rect 14188 992 14240 1012
rect 14240 992 14242 1012
rect 14554 1808 14610 1864
rect 14554 1128 14610 1184
rect 15014 1672 15070 1728
rect 16364 10362 16420 10364
rect 16444 10362 16500 10364
rect 16524 10362 16580 10364
rect 16604 10362 16660 10364
rect 16684 10362 16740 10364
rect 16364 10310 16366 10362
rect 16366 10310 16418 10362
rect 16418 10310 16420 10362
rect 16444 10310 16482 10362
rect 16482 10310 16494 10362
rect 16494 10310 16500 10362
rect 16524 10310 16546 10362
rect 16546 10310 16558 10362
rect 16558 10310 16580 10362
rect 16604 10310 16610 10362
rect 16610 10310 16622 10362
rect 16622 10310 16660 10362
rect 16684 10310 16686 10362
rect 16686 10310 16738 10362
rect 16738 10310 16740 10362
rect 16364 10308 16420 10310
rect 16444 10308 16500 10310
rect 16524 10308 16580 10310
rect 16604 10308 16660 10310
rect 16684 10308 16740 10310
rect 16394 9988 16450 10024
rect 16394 9968 16396 9988
rect 16396 9968 16448 9988
rect 16448 9968 16450 9988
rect 16762 9696 16818 9752
rect 16394 9580 16450 9616
rect 16394 9560 16396 9580
rect 16396 9560 16448 9580
rect 16448 9560 16450 9580
rect 16762 9560 16818 9616
rect 16670 9460 16672 9480
rect 16672 9460 16724 9480
rect 16724 9460 16726 9480
rect 16670 9424 16726 9460
rect 16364 9274 16420 9276
rect 16444 9274 16500 9276
rect 16524 9274 16580 9276
rect 16604 9274 16660 9276
rect 16684 9274 16740 9276
rect 16364 9222 16366 9274
rect 16366 9222 16418 9274
rect 16418 9222 16420 9274
rect 16444 9222 16482 9274
rect 16482 9222 16494 9274
rect 16494 9222 16500 9274
rect 16524 9222 16546 9274
rect 16546 9222 16558 9274
rect 16558 9222 16580 9274
rect 16604 9222 16610 9274
rect 16610 9222 16622 9274
rect 16622 9222 16660 9274
rect 16684 9222 16686 9274
rect 16686 9222 16738 9274
rect 16738 9222 16740 9274
rect 16364 9220 16420 9222
rect 16444 9220 16500 9222
rect 16524 9220 16580 9222
rect 16604 9220 16660 9222
rect 16684 9220 16740 9222
rect 16946 10920 17002 10976
rect 16364 8186 16420 8188
rect 16444 8186 16500 8188
rect 16524 8186 16580 8188
rect 16604 8186 16660 8188
rect 16684 8186 16740 8188
rect 16364 8134 16366 8186
rect 16366 8134 16418 8186
rect 16418 8134 16420 8186
rect 16444 8134 16482 8186
rect 16482 8134 16494 8186
rect 16494 8134 16500 8186
rect 16524 8134 16546 8186
rect 16546 8134 16558 8186
rect 16558 8134 16580 8186
rect 16604 8134 16610 8186
rect 16610 8134 16622 8186
rect 16622 8134 16660 8186
rect 16684 8134 16686 8186
rect 16686 8134 16738 8186
rect 16738 8134 16740 8186
rect 16364 8132 16420 8134
rect 16444 8132 16500 8134
rect 16524 8132 16580 8134
rect 16604 8132 16660 8134
rect 16684 8132 16740 8134
rect 16364 7098 16420 7100
rect 16444 7098 16500 7100
rect 16524 7098 16580 7100
rect 16604 7098 16660 7100
rect 16684 7098 16740 7100
rect 16364 7046 16366 7098
rect 16366 7046 16418 7098
rect 16418 7046 16420 7098
rect 16444 7046 16482 7098
rect 16482 7046 16494 7098
rect 16494 7046 16500 7098
rect 16524 7046 16546 7098
rect 16546 7046 16558 7098
rect 16558 7046 16580 7098
rect 16604 7046 16610 7098
rect 16610 7046 16622 7098
rect 16622 7046 16660 7098
rect 16684 7046 16686 7098
rect 16686 7046 16738 7098
rect 16738 7046 16740 7098
rect 16364 7044 16420 7046
rect 16444 7044 16500 7046
rect 16524 7044 16580 7046
rect 16604 7044 16660 7046
rect 16684 7044 16740 7046
rect 16302 6196 16304 6216
rect 16304 6196 16356 6216
rect 16356 6196 16358 6216
rect 16302 6160 16358 6196
rect 16364 6010 16420 6012
rect 16444 6010 16500 6012
rect 16524 6010 16580 6012
rect 16604 6010 16660 6012
rect 16684 6010 16740 6012
rect 16364 5958 16366 6010
rect 16366 5958 16418 6010
rect 16418 5958 16420 6010
rect 16444 5958 16482 6010
rect 16482 5958 16494 6010
rect 16494 5958 16500 6010
rect 16524 5958 16546 6010
rect 16546 5958 16558 6010
rect 16558 5958 16580 6010
rect 16604 5958 16610 6010
rect 16610 5958 16622 6010
rect 16622 5958 16660 6010
rect 16684 5958 16686 6010
rect 16686 5958 16738 6010
rect 16738 5958 16740 6010
rect 16364 5956 16420 5958
rect 16444 5956 16500 5958
rect 16524 5956 16580 5958
rect 16604 5956 16660 5958
rect 16684 5956 16740 5958
rect 17130 10920 17186 10976
rect 17130 9052 17132 9072
rect 17132 9052 17184 9072
rect 17184 9052 17186 9072
rect 17130 9016 17186 9052
rect 17958 21664 18014 21720
rect 19364 22874 19420 22876
rect 19444 22874 19500 22876
rect 19524 22874 19580 22876
rect 19604 22874 19660 22876
rect 19684 22874 19740 22876
rect 19364 22822 19366 22874
rect 19366 22822 19418 22874
rect 19418 22822 19420 22874
rect 19444 22822 19482 22874
rect 19482 22822 19494 22874
rect 19494 22822 19500 22874
rect 19524 22822 19546 22874
rect 19546 22822 19558 22874
rect 19558 22822 19580 22874
rect 19604 22822 19610 22874
rect 19610 22822 19622 22874
rect 19622 22822 19660 22874
rect 19684 22822 19686 22874
rect 19686 22822 19738 22874
rect 19738 22822 19740 22874
rect 19364 22820 19420 22822
rect 19444 22820 19500 22822
rect 19524 22820 19580 22822
rect 19604 22820 19660 22822
rect 19684 22820 19740 22822
rect 19246 22072 19302 22128
rect 18602 19896 18658 19952
rect 18694 19624 18750 19680
rect 18878 20984 18934 21040
rect 17590 15952 17646 16008
rect 17498 12008 17554 12064
rect 17314 9152 17370 9208
rect 17590 10648 17646 10704
rect 18050 12300 18106 12336
rect 18050 12280 18052 12300
rect 18052 12280 18104 12300
rect 18104 12280 18106 12300
rect 18142 11600 18198 11656
rect 17774 10784 17830 10840
rect 17774 10240 17830 10296
rect 17682 9152 17738 9208
rect 17866 9460 17868 9480
rect 17868 9460 17920 9480
rect 17920 9460 17922 9480
rect 17866 9424 17922 9460
rect 17590 8608 17646 8664
rect 17498 8064 17554 8120
rect 17498 7248 17554 7304
rect 16364 4922 16420 4924
rect 16444 4922 16500 4924
rect 16524 4922 16580 4924
rect 16604 4922 16660 4924
rect 16684 4922 16740 4924
rect 16364 4870 16366 4922
rect 16366 4870 16418 4922
rect 16418 4870 16420 4922
rect 16444 4870 16482 4922
rect 16482 4870 16494 4922
rect 16494 4870 16500 4922
rect 16524 4870 16546 4922
rect 16546 4870 16558 4922
rect 16558 4870 16580 4922
rect 16604 4870 16610 4922
rect 16610 4870 16622 4922
rect 16622 4870 16660 4922
rect 16684 4870 16686 4922
rect 16686 4870 16738 4922
rect 16738 4870 16740 4922
rect 16364 4868 16420 4870
rect 16444 4868 16500 4870
rect 16524 4868 16580 4870
rect 16604 4868 16660 4870
rect 16684 4868 16740 4870
rect 16302 4140 16358 4176
rect 16302 4120 16304 4140
rect 16304 4120 16356 4140
rect 16356 4120 16358 4140
rect 16364 3834 16420 3836
rect 16444 3834 16500 3836
rect 16524 3834 16580 3836
rect 16604 3834 16660 3836
rect 16684 3834 16740 3836
rect 16364 3782 16366 3834
rect 16366 3782 16418 3834
rect 16418 3782 16420 3834
rect 16444 3782 16482 3834
rect 16482 3782 16494 3834
rect 16494 3782 16500 3834
rect 16524 3782 16546 3834
rect 16546 3782 16558 3834
rect 16558 3782 16580 3834
rect 16604 3782 16610 3834
rect 16610 3782 16622 3834
rect 16622 3782 16660 3834
rect 16684 3782 16686 3834
rect 16686 3782 16738 3834
rect 16738 3782 16740 3834
rect 16364 3780 16420 3782
rect 16444 3780 16500 3782
rect 16524 3780 16580 3782
rect 16604 3780 16660 3782
rect 16684 3780 16740 3782
rect 15198 2508 15254 2544
rect 15198 2488 15200 2508
rect 15200 2488 15252 2508
rect 15252 2488 15254 2508
rect 15198 1536 15254 1592
rect 16364 2746 16420 2748
rect 16444 2746 16500 2748
rect 16524 2746 16580 2748
rect 16604 2746 16660 2748
rect 16684 2746 16740 2748
rect 16364 2694 16366 2746
rect 16366 2694 16418 2746
rect 16418 2694 16420 2746
rect 16444 2694 16482 2746
rect 16482 2694 16494 2746
rect 16494 2694 16500 2746
rect 16524 2694 16546 2746
rect 16546 2694 16558 2746
rect 16558 2694 16580 2746
rect 16604 2694 16610 2746
rect 16610 2694 16622 2746
rect 16622 2694 16660 2746
rect 16684 2694 16686 2746
rect 16686 2694 16738 2746
rect 16738 2694 16740 2746
rect 16364 2692 16420 2694
rect 16444 2692 16500 2694
rect 16524 2692 16580 2694
rect 16604 2692 16660 2694
rect 16684 2692 16740 2694
rect 16302 2508 16358 2544
rect 16302 2488 16304 2508
rect 16304 2488 16356 2508
rect 16356 2488 16358 2508
rect 15934 1536 15990 1592
rect 16364 1658 16420 1660
rect 16444 1658 16500 1660
rect 16524 1658 16580 1660
rect 16604 1658 16660 1660
rect 16684 1658 16740 1660
rect 16364 1606 16366 1658
rect 16366 1606 16418 1658
rect 16418 1606 16420 1658
rect 16444 1606 16482 1658
rect 16482 1606 16494 1658
rect 16494 1606 16500 1658
rect 16524 1606 16546 1658
rect 16546 1606 16558 1658
rect 16558 1606 16580 1658
rect 16604 1606 16610 1658
rect 16610 1606 16622 1658
rect 16622 1606 16660 1658
rect 16684 1606 16686 1658
rect 16686 1606 16738 1658
rect 16738 1606 16740 1658
rect 16364 1604 16420 1606
rect 16444 1604 16500 1606
rect 16524 1604 16580 1606
rect 16604 1604 16660 1606
rect 16684 1604 16740 1606
rect 17406 5208 17462 5264
rect 17866 8608 17922 8664
rect 17958 8200 18014 8256
rect 17774 7792 17830 7848
rect 18510 15000 18566 15056
rect 19338 21936 19394 21992
rect 19364 21786 19420 21788
rect 19444 21786 19500 21788
rect 19524 21786 19580 21788
rect 19604 21786 19660 21788
rect 19684 21786 19740 21788
rect 19364 21734 19366 21786
rect 19366 21734 19418 21786
rect 19418 21734 19420 21786
rect 19444 21734 19482 21786
rect 19482 21734 19494 21786
rect 19494 21734 19500 21786
rect 19524 21734 19546 21786
rect 19546 21734 19558 21786
rect 19558 21734 19580 21786
rect 19604 21734 19610 21786
rect 19610 21734 19622 21786
rect 19622 21734 19660 21786
rect 19684 21734 19686 21786
rect 19686 21734 19738 21786
rect 19738 21734 19740 21786
rect 19364 21732 19420 21734
rect 19444 21732 19500 21734
rect 19524 21732 19580 21734
rect 19604 21732 19660 21734
rect 19684 21732 19740 21734
rect 19982 21664 20038 21720
rect 20074 21528 20130 21584
rect 20074 21256 20130 21312
rect 19430 20848 19486 20904
rect 19364 20698 19420 20700
rect 19444 20698 19500 20700
rect 19524 20698 19580 20700
rect 19604 20698 19660 20700
rect 19684 20698 19740 20700
rect 19364 20646 19366 20698
rect 19366 20646 19418 20698
rect 19418 20646 19420 20698
rect 19444 20646 19482 20698
rect 19482 20646 19494 20698
rect 19494 20646 19500 20698
rect 19524 20646 19546 20698
rect 19546 20646 19558 20698
rect 19558 20646 19580 20698
rect 19604 20646 19610 20698
rect 19610 20646 19622 20698
rect 19622 20646 19660 20698
rect 19684 20646 19686 20698
rect 19686 20646 19738 20698
rect 19738 20646 19740 20698
rect 19364 20644 19420 20646
rect 19444 20644 19500 20646
rect 19524 20644 19580 20646
rect 19604 20644 19660 20646
rect 19684 20644 19740 20646
rect 19890 20304 19946 20360
rect 18970 19352 19026 19408
rect 19364 19610 19420 19612
rect 19444 19610 19500 19612
rect 19524 19610 19580 19612
rect 19604 19610 19660 19612
rect 19684 19610 19740 19612
rect 19364 19558 19366 19610
rect 19366 19558 19418 19610
rect 19418 19558 19420 19610
rect 19444 19558 19482 19610
rect 19482 19558 19494 19610
rect 19494 19558 19500 19610
rect 19524 19558 19546 19610
rect 19546 19558 19558 19610
rect 19558 19558 19580 19610
rect 19604 19558 19610 19610
rect 19610 19558 19622 19610
rect 19622 19558 19660 19610
rect 19684 19558 19686 19610
rect 19686 19558 19738 19610
rect 19738 19558 19740 19610
rect 19364 19556 19420 19558
rect 19444 19556 19500 19558
rect 19524 19556 19580 19558
rect 19604 19556 19660 19558
rect 19684 19556 19740 19558
rect 20074 19624 20130 19680
rect 19364 18522 19420 18524
rect 19444 18522 19500 18524
rect 19524 18522 19580 18524
rect 19604 18522 19660 18524
rect 19684 18522 19740 18524
rect 19364 18470 19366 18522
rect 19366 18470 19418 18522
rect 19418 18470 19420 18522
rect 19444 18470 19482 18522
rect 19482 18470 19494 18522
rect 19494 18470 19500 18522
rect 19524 18470 19546 18522
rect 19546 18470 19558 18522
rect 19558 18470 19580 18522
rect 19604 18470 19610 18522
rect 19610 18470 19622 18522
rect 19622 18470 19660 18522
rect 19684 18470 19686 18522
rect 19686 18470 19738 18522
rect 19738 18470 19740 18522
rect 19364 18468 19420 18470
rect 19444 18468 19500 18470
rect 19524 18468 19580 18470
rect 19604 18468 19660 18470
rect 19684 18468 19740 18470
rect 19364 17434 19420 17436
rect 19444 17434 19500 17436
rect 19524 17434 19580 17436
rect 19604 17434 19660 17436
rect 19684 17434 19740 17436
rect 19364 17382 19366 17434
rect 19366 17382 19418 17434
rect 19418 17382 19420 17434
rect 19444 17382 19482 17434
rect 19482 17382 19494 17434
rect 19494 17382 19500 17434
rect 19524 17382 19546 17434
rect 19546 17382 19558 17434
rect 19558 17382 19580 17434
rect 19604 17382 19610 17434
rect 19610 17382 19622 17434
rect 19622 17382 19660 17434
rect 19684 17382 19686 17434
rect 19686 17382 19738 17434
rect 19738 17382 19740 17434
rect 19364 17380 19420 17382
rect 19444 17380 19500 17382
rect 19524 17380 19580 17382
rect 19604 17380 19660 17382
rect 19684 17380 19740 17382
rect 19364 16346 19420 16348
rect 19444 16346 19500 16348
rect 19524 16346 19580 16348
rect 19604 16346 19660 16348
rect 19684 16346 19740 16348
rect 19364 16294 19366 16346
rect 19366 16294 19418 16346
rect 19418 16294 19420 16346
rect 19444 16294 19482 16346
rect 19482 16294 19494 16346
rect 19494 16294 19500 16346
rect 19524 16294 19546 16346
rect 19546 16294 19558 16346
rect 19558 16294 19580 16346
rect 19604 16294 19610 16346
rect 19610 16294 19622 16346
rect 19622 16294 19660 16346
rect 19684 16294 19686 16346
rect 19686 16294 19738 16346
rect 19738 16294 19740 16346
rect 19364 16292 19420 16294
rect 19444 16292 19500 16294
rect 19524 16292 19580 16294
rect 19604 16292 19660 16294
rect 19684 16292 19740 16294
rect 18694 15544 18750 15600
rect 18694 14184 18750 14240
rect 18326 11872 18382 11928
rect 18326 11076 18382 11112
rect 18326 11056 18328 11076
rect 18328 11056 18380 11076
rect 18380 11056 18382 11076
rect 18234 10512 18290 10568
rect 18234 9696 18290 9752
rect 18142 9172 18198 9208
rect 18142 9152 18144 9172
rect 18144 9152 18196 9172
rect 18196 9152 18198 9172
rect 18142 9016 18198 9072
rect 18234 8880 18290 8936
rect 18142 7520 18198 7576
rect 18418 9832 18474 9888
rect 18694 11464 18750 11520
rect 18602 9968 18658 10024
rect 19338 15408 19394 15464
rect 19364 15258 19420 15260
rect 19444 15258 19500 15260
rect 19524 15258 19580 15260
rect 19604 15258 19660 15260
rect 19684 15258 19740 15260
rect 19364 15206 19366 15258
rect 19366 15206 19418 15258
rect 19418 15206 19420 15258
rect 19444 15206 19482 15258
rect 19482 15206 19494 15258
rect 19494 15206 19500 15258
rect 19524 15206 19546 15258
rect 19546 15206 19558 15258
rect 19558 15206 19580 15258
rect 19604 15206 19610 15258
rect 19610 15206 19622 15258
rect 19622 15206 19660 15258
rect 19684 15206 19686 15258
rect 19686 15206 19738 15258
rect 19738 15206 19740 15258
rect 19364 15204 19420 15206
rect 19444 15204 19500 15206
rect 19524 15204 19580 15206
rect 19604 15204 19660 15206
rect 19684 15204 19740 15206
rect 21638 22924 21640 22944
rect 21640 22924 21692 22944
rect 21692 22924 21694 22944
rect 21086 22208 21142 22264
rect 20718 20848 20774 20904
rect 20810 20476 20812 20496
rect 20812 20476 20864 20496
rect 20864 20476 20866 20496
rect 20810 20440 20866 20476
rect 20626 20304 20682 20360
rect 19890 18536 19946 18592
rect 19890 16496 19946 16552
rect 19338 14456 19394 14512
rect 20626 19916 20682 19952
rect 20626 19896 20628 19916
rect 20628 19896 20680 19916
rect 20680 19896 20682 19916
rect 20626 19624 20682 19680
rect 20810 19780 20866 19816
rect 20810 19760 20812 19780
rect 20812 19760 20864 19780
rect 20864 19760 20866 19780
rect 20626 19252 20628 19272
rect 20628 19252 20680 19272
rect 20680 19252 20682 19272
rect 20626 19216 20682 19252
rect 20534 17992 20590 18048
rect 19364 14170 19420 14172
rect 19444 14170 19500 14172
rect 19524 14170 19580 14172
rect 19604 14170 19660 14172
rect 19684 14170 19740 14172
rect 19364 14118 19366 14170
rect 19366 14118 19418 14170
rect 19418 14118 19420 14170
rect 19444 14118 19482 14170
rect 19482 14118 19494 14170
rect 19494 14118 19500 14170
rect 19524 14118 19546 14170
rect 19546 14118 19558 14170
rect 19558 14118 19580 14170
rect 19604 14118 19610 14170
rect 19610 14118 19622 14170
rect 19622 14118 19660 14170
rect 19684 14118 19686 14170
rect 19686 14118 19738 14170
rect 19738 14118 19740 14170
rect 19364 14116 19420 14118
rect 19444 14116 19500 14118
rect 19524 14116 19580 14118
rect 19604 14116 19660 14118
rect 19684 14116 19740 14118
rect 19364 13082 19420 13084
rect 19444 13082 19500 13084
rect 19524 13082 19580 13084
rect 19604 13082 19660 13084
rect 19684 13082 19740 13084
rect 19364 13030 19366 13082
rect 19366 13030 19418 13082
rect 19418 13030 19420 13082
rect 19444 13030 19482 13082
rect 19482 13030 19494 13082
rect 19494 13030 19500 13082
rect 19524 13030 19546 13082
rect 19546 13030 19558 13082
rect 19558 13030 19580 13082
rect 19604 13030 19610 13082
rect 19610 13030 19622 13082
rect 19622 13030 19660 13082
rect 19684 13030 19686 13082
rect 19686 13030 19738 13082
rect 19738 13030 19740 13082
rect 19364 13028 19420 13030
rect 19444 13028 19500 13030
rect 19524 13028 19580 13030
rect 19604 13028 19660 13030
rect 19684 13028 19740 13030
rect 19338 12824 19394 12880
rect 19522 12824 19578 12880
rect 19522 12164 19578 12200
rect 19522 12144 19524 12164
rect 19524 12144 19576 12164
rect 19576 12144 19578 12164
rect 19364 11994 19420 11996
rect 19444 11994 19500 11996
rect 19524 11994 19580 11996
rect 19604 11994 19660 11996
rect 19684 11994 19740 11996
rect 19364 11942 19366 11994
rect 19366 11942 19418 11994
rect 19418 11942 19420 11994
rect 19444 11942 19482 11994
rect 19482 11942 19494 11994
rect 19494 11942 19500 11994
rect 19524 11942 19546 11994
rect 19546 11942 19558 11994
rect 19558 11942 19580 11994
rect 19604 11942 19610 11994
rect 19610 11942 19622 11994
rect 19622 11942 19660 11994
rect 19684 11942 19686 11994
rect 19686 11942 19738 11994
rect 19738 11942 19740 11994
rect 19364 11940 19420 11942
rect 19444 11940 19500 11942
rect 19524 11940 19580 11942
rect 19604 11940 19660 11942
rect 19684 11940 19740 11942
rect 19522 11736 19578 11792
rect 19062 11500 19064 11520
rect 19064 11500 19116 11520
rect 19116 11500 19118 11520
rect 19062 11464 19118 11500
rect 18878 11192 18934 11248
rect 18786 9288 18842 9344
rect 19338 11092 19340 11112
rect 19340 11092 19392 11112
rect 19392 11092 19394 11112
rect 19338 11056 19394 11092
rect 19364 10906 19420 10908
rect 19444 10906 19500 10908
rect 19524 10906 19580 10908
rect 19604 10906 19660 10908
rect 19684 10906 19740 10908
rect 19364 10854 19366 10906
rect 19366 10854 19418 10906
rect 19418 10854 19420 10906
rect 19444 10854 19482 10906
rect 19482 10854 19494 10906
rect 19494 10854 19500 10906
rect 19524 10854 19546 10906
rect 19546 10854 19558 10906
rect 19558 10854 19580 10906
rect 19604 10854 19610 10906
rect 19610 10854 19622 10906
rect 19622 10854 19660 10906
rect 19684 10854 19686 10906
rect 19686 10854 19738 10906
rect 19738 10854 19740 10906
rect 19364 10852 19420 10854
rect 19444 10852 19500 10854
rect 19524 10852 19580 10854
rect 19604 10852 19660 10854
rect 19684 10852 19740 10854
rect 19246 10648 19302 10704
rect 19614 10512 19670 10568
rect 19364 9818 19420 9820
rect 19444 9818 19500 9820
rect 19524 9818 19580 9820
rect 19604 9818 19660 9820
rect 19684 9818 19740 9820
rect 19364 9766 19366 9818
rect 19366 9766 19418 9818
rect 19418 9766 19420 9818
rect 19444 9766 19482 9818
rect 19482 9766 19494 9818
rect 19494 9766 19500 9818
rect 19524 9766 19546 9818
rect 19546 9766 19558 9818
rect 19558 9766 19580 9818
rect 19604 9766 19610 9818
rect 19610 9766 19622 9818
rect 19622 9766 19660 9818
rect 19684 9766 19686 9818
rect 19686 9766 19738 9818
rect 19738 9766 19740 9818
rect 19364 9764 19420 9766
rect 19444 9764 19500 9766
rect 19524 9764 19580 9766
rect 19604 9764 19660 9766
rect 19684 9764 19740 9766
rect 19430 9460 19432 9480
rect 19432 9460 19484 9480
rect 19484 9460 19486 9480
rect 19430 9424 19486 9460
rect 18418 8608 18474 8664
rect 18418 7928 18474 7984
rect 18694 8608 18750 8664
rect 18694 7792 18750 7848
rect 19338 9152 19394 9208
rect 19062 9036 19118 9072
rect 19062 9016 19064 9036
rect 19064 9016 19116 9036
rect 19116 9016 19118 9036
rect 20166 12824 20222 12880
rect 21638 22888 21694 22924
rect 21454 21664 21510 21720
rect 21546 21392 21602 21448
rect 21822 21392 21878 21448
rect 21454 21292 21456 21312
rect 21456 21292 21508 21312
rect 21508 21292 21510 21312
rect 21454 21256 21510 21292
rect 21362 19760 21418 19816
rect 21270 19352 21326 19408
rect 20718 17584 20774 17640
rect 20810 17040 20866 17096
rect 20718 16652 20774 16688
rect 20718 16632 20720 16652
rect 20720 16632 20772 16652
rect 20772 16632 20774 16652
rect 20258 11192 20314 11248
rect 19890 9424 19946 9480
rect 19246 8880 19302 8936
rect 19706 8880 19762 8936
rect 20074 9460 20076 9480
rect 20076 9460 20128 9480
rect 20128 9460 20130 9480
rect 20074 9424 20130 9460
rect 18970 8744 19026 8800
rect 19154 8200 19210 8256
rect 18970 7656 19026 7712
rect 18050 4564 18052 4584
rect 18052 4564 18104 4584
rect 18104 4564 18106 4584
rect 18050 4528 18106 4564
rect 17682 2352 17738 2408
rect 17866 2372 17922 2408
rect 17866 2352 17868 2372
rect 17868 2352 17920 2372
rect 17920 2352 17922 2372
rect 19364 8730 19420 8732
rect 19444 8730 19500 8732
rect 19524 8730 19580 8732
rect 19604 8730 19660 8732
rect 19684 8730 19740 8732
rect 19364 8678 19366 8730
rect 19366 8678 19418 8730
rect 19418 8678 19420 8730
rect 19444 8678 19482 8730
rect 19482 8678 19494 8730
rect 19494 8678 19500 8730
rect 19524 8678 19546 8730
rect 19546 8678 19558 8730
rect 19558 8678 19580 8730
rect 19604 8678 19610 8730
rect 19610 8678 19622 8730
rect 19622 8678 19660 8730
rect 19684 8678 19686 8730
rect 19686 8678 19738 8730
rect 19738 8678 19740 8730
rect 19364 8676 19420 8678
rect 19444 8676 19500 8678
rect 19524 8676 19580 8678
rect 19604 8676 19660 8678
rect 19684 8676 19740 8678
rect 19364 7642 19420 7644
rect 19444 7642 19500 7644
rect 19524 7642 19580 7644
rect 19604 7642 19660 7644
rect 19684 7642 19740 7644
rect 19364 7590 19366 7642
rect 19366 7590 19418 7642
rect 19418 7590 19420 7642
rect 19444 7590 19482 7642
rect 19482 7590 19494 7642
rect 19494 7590 19500 7642
rect 19524 7590 19546 7642
rect 19546 7590 19558 7642
rect 19558 7590 19580 7642
rect 19604 7590 19610 7642
rect 19610 7590 19622 7642
rect 19622 7590 19660 7642
rect 19684 7590 19686 7642
rect 19686 7590 19738 7642
rect 19738 7590 19740 7642
rect 19364 7588 19420 7590
rect 19444 7588 19500 7590
rect 19524 7588 19580 7590
rect 19604 7588 19660 7590
rect 19684 7588 19740 7590
rect 19246 7384 19302 7440
rect 19614 7384 19670 7440
rect 19798 6840 19854 6896
rect 19706 6704 19762 6760
rect 19364 6554 19420 6556
rect 19444 6554 19500 6556
rect 19524 6554 19580 6556
rect 19604 6554 19660 6556
rect 19684 6554 19740 6556
rect 19364 6502 19366 6554
rect 19366 6502 19418 6554
rect 19418 6502 19420 6554
rect 19444 6502 19482 6554
rect 19482 6502 19494 6554
rect 19494 6502 19500 6554
rect 19524 6502 19546 6554
rect 19546 6502 19558 6554
rect 19558 6502 19580 6554
rect 19604 6502 19610 6554
rect 19610 6502 19622 6554
rect 19622 6502 19660 6554
rect 19684 6502 19686 6554
rect 19686 6502 19738 6554
rect 19738 6502 19740 6554
rect 19364 6500 19420 6502
rect 19444 6500 19500 6502
rect 19524 6500 19580 6502
rect 19604 6500 19660 6502
rect 19684 6500 19740 6502
rect 19430 6296 19486 6352
rect 19522 5772 19578 5808
rect 19522 5752 19524 5772
rect 19524 5752 19576 5772
rect 19576 5752 19578 5772
rect 19364 5466 19420 5468
rect 19444 5466 19500 5468
rect 19524 5466 19580 5468
rect 19604 5466 19660 5468
rect 19684 5466 19740 5468
rect 19364 5414 19366 5466
rect 19366 5414 19418 5466
rect 19418 5414 19420 5466
rect 19444 5414 19482 5466
rect 19482 5414 19494 5466
rect 19494 5414 19500 5466
rect 19524 5414 19546 5466
rect 19546 5414 19558 5466
rect 19558 5414 19580 5466
rect 19604 5414 19610 5466
rect 19610 5414 19622 5466
rect 19622 5414 19660 5466
rect 19684 5414 19686 5466
rect 19686 5414 19738 5466
rect 19738 5414 19740 5466
rect 19364 5412 19420 5414
rect 19444 5412 19500 5414
rect 19524 5412 19580 5414
rect 19604 5412 19660 5414
rect 19684 5412 19740 5414
rect 19706 5208 19762 5264
rect 19154 5072 19210 5128
rect 18510 2624 18566 2680
rect 18050 2216 18106 2272
rect 17774 1944 17830 2000
rect 16854 1128 16910 1184
rect 16364 570 16420 572
rect 16444 570 16500 572
rect 16524 570 16580 572
rect 16604 570 16660 572
rect 16684 570 16740 572
rect 16364 518 16366 570
rect 16366 518 16418 570
rect 16418 518 16420 570
rect 16444 518 16482 570
rect 16482 518 16494 570
rect 16494 518 16500 570
rect 16524 518 16546 570
rect 16546 518 16558 570
rect 16558 518 16580 570
rect 16604 518 16610 570
rect 16610 518 16622 570
rect 16622 518 16660 570
rect 16684 518 16686 570
rect 16686 518 16738 570
rect 16738 518 16740 570
rect 16364 516 16420 518
rect 16444 516 16500 518
rect 16524 516 16580 518
rect 16604 516 16660 518
rect 16684 516 16740 518
rect 19062 4256 19118 4312
rect 18878 3476 18880 3496
rect 18880 3476 18932 3496
rect 18932 3476 18934 3496
rect 18878 3440 18934 3476
rect 20810 12824 20866 12880
rect 20626 12180 20628 12200
rect 20628 12180 20680 12200
rect 20680 12180 20682 12200
rect 20626 12144 20682 12180
rect 20350 9288 20406 9344
rect 20258 6860 20314 6896
rect 20258 6840 20260 6860
rect 20260 6840 20312 6860
rect 20312 6840 20314 6860
rect 20074 5616 20130 5672
rect 19364 4378 19420 4380
rect 19444 4378 19500 4380
rect 19524 4378 19580 4380
rect 19604 4378 19660 4380
rect 19684 4378 19740 4380
rect 19364 4326 19366 4378
rect 19366 4326 19418 4378
rect 19418 4326 19420 4378
rect 19444 4326 19482 4378
rect 19482 4326 19494 4378
rect 19494 4326 19500 4378
rect 19524 4326 19546 4378
rect 19546 4326 19558 4378
rect 19558 4326 19580 4378
rect 19604 4326 19610 4378
rect 19610 4326 19622 4378
rect 19622 4326 19660 4378
rect 19684 4326 19686 4378
rect 19686 4326 19738 4378
rect 19738 4326 19740 4378
rect 19364 4324 19420 4326
rect 19444 4324 19500 4326
rect 19524 4324 19580 4326
rect 19604 4324 19660 4326
rect 19684 4324 19740 4326
rect 19982 3984 20038 4040
rect 19522 3596 19578 3632
rect 19522 3576 19524 3596
rect 19524 3576 19576 3596
rect 19576 3576 19578 3596
rect 19890 3596 19946 3632
rect 19890 3576 19892 3596
rect 19892 3576 19944 3596
rect 19944 3576 19946 3596
rect 19338 3476 19340 3496
rect 19340 3476 19392 3496
rect 19392 3476 19394 3496
rect 19338 3440 19394 3476
rect 19364 3290 19420 3292
rect 19444 3290 19500 3292
rect 19524 3290 19580 3292
rect 19604 3290 19660 3292
rect 19684 3290 19740 3292
rect 19364 3238 19366 3290
rect 19366 3238 19418 3290
rect 19418 3238 19420 3290
rect 19444 3238 19482 3290
rect 19482 3238 19494 3290
rect 19494 3238 19500 3290
rect 19524 3238 19546 3290
rect 19546 3238 19558 3290
rect 19558 3238 19580 3290
rect 19604 3238 19610 3290
rect 19610 3238 19622 3290
rect 19622 3238 19660 3290
rect 19684 3238 19686 3290
rect 19686 3238 19738 3290
rect 19738 3238 19740 3290
rect 19364 3236 19420 3238
rect 19444 3236 19500 3238
rect 19524 3236 19580 3238
rect 19604 3236 19660 3238
rect 19684 3236 19740 3238
rect 20258 4020 20260 4040
rect 20260 4020 20312 4040
rect 20312 4020 20314 4040
rect 20258 3984 20314 4020
rect 18694 1944 18750 2000
rect 17866 992 17922 1048
rect 18602 720 18658 776
rect 17866 176 17922 232
rect 17590 40 17646 96
rect 19364 2202 19420 2204
rect 19444 2202 19500 2204
rect 19524 2202 19580 2204
rect 19604 2202 19660 2204
rect 19684 2202 19740 2204
rect 19364 2150 19366 2202
rect 19366 2150 19418 2202
rect 19418 2150 19420 2202
rect 19444 2150 19482 2202
rect 19482 2150 19494 2202
rect 19494 2150 19500 2202
rect 19524 2150 19546 2202
rect 19546 2150 19558 2202
rect 19558 2150 19580 2202
rect 19604 2150 19610 2202
rect 19610 2150 19622 2202
rect 19622 2150 19660 2202
rect 19684 2150 19686 2202
rect 19686 2150 19738 2202
rect 19738 2150 19740 2202
rect 19364 2148 19420 2150
rect 19444 2148 19500 2150
rect 19524 2148 19580 2150
rect 19604 2148 19660 2150
rect 19684 2148 19740 2150
rect 19338 1708 19340 1728
rect 19340 1708 19392 1728
rect 19392 1708 19394 1728
rect 19338 1672 19394 1708
rect 19706 1420 19762 1456
rect 19890 2216 19946 2272
rect 20074 2352 20130 2408
rect 19706 1400 19708 1420
rect 19708 1400 19760 1420
rect 19760 1400 19762 1420
rect 19798 1264 19854 1320
rect 19364 1114 19420 1116
rect 19444 1114 19500 1116
rect 19524 1114 19580 1116
rect 19604 1114 19660 1116
rect 19684 1114 19740 1116
rect 19364 1062 19366 1114
rect 19366 1062 19418 1114
rect 19418 1062 19420 1114
rect 19444 1062 19482 1114
rect 19482 1062 19494 1114
rect 19494 1062 19500 1114
rect 19524 1062 19546 1114
rect 19546 1062 19558 1114
rect 19558 1062 19580 1114
rect 19604 1062 19610 1114
rect 19610 1062 19622 1114
rect 19622 1062 19660 1114
rect 19684 1062 19686 1114
rect 19686 1062 19738 1114
rect 19738 1062 19740 1114
rect 19364 1060 19420 1062
rect 19444 1060 19500 1062
rect 19524 1060 19580 1062
rect 19604 1060 19660 1062
rect 19684 1060 19740 1062
rect 19890 992 19946 1048
rect 20074 1400 20130 1456
rect 21546 18028 21548 18048
rect 21548 18028 21600 18048
rect 21600 18028 21602 18048
rect 21546 17992 21602 18028
rect 21822 18536 21878 18592
rect 22364 23418 22420 23420
rect 22444 23418 22500 23420
rect 22524 23418 22580 23420
rect 22604 23418 22660 23420
rect 22684 23418 22740 23420
rect 22364 23366 22366 23418
rect 22366 23366 22418 23418
rect 22418 23366 22420 23418
rect 22444 23366 22482 23418
rect 22482 23366 22494 23418
rect 22494 23366 22500 23418
rect 22524 23366 22546 23418
rect 22546 23366 22558 23418
rect 22558 23366 22580 23418
rect 22604 23366 22610 23418
rect 22610 23366 22622 23418
rect 22622 23366 22660 23418
rect 22684 23366 22686 23418
rect 22686 23366 22738 23418
rect 22738 23366 22740 23418
rect 22364 23364 22420 23366
rect 22444 23364 22500 23366
rect 22524 23364 22580 23366
rect 22604 23364 22660 23366
rect 22684 23364 22740 23366
rect 22364 22330 22420 22332
rect 22444 22330 22500 22332
rect 22524 22330 22580 22332
rect 22604 22330 22660 22332
rect 22684 22330 22740 22332
rect 22364 22278 22366 22330
rect 22366 22278 22418 22330
rect 22418 22278 22420 22330
rect 22444 22278 22482 22330
rect 22482 22278 22494 22330
rect 22494 22278 22500 22330
rect 22524 22278 22546 22330
rect 22546 22278 22558 22330
rect 22558 22278 22580 22330
rect 22604 22278 22610 22330
rect 22610 22278 22622 22330
rect 22622 22278 22660 22330
rect 22684 22278 22686 22330
rect 22686 22278 22738 22330
rect 22738 22278 22740 22330
rect 22364 22276 22420 22278
rect 22444 22276 22500 22278
rect 22524 22276 22580 22278
rect 22604 22276 22660 22278
rect 22684 22276 22740 22278
rect 22006 19352 22062 19408
rect 22364 21242 22420 21244
rect 22444 21242 22500 21244
rect 22524 21242 22580 21244
rect 22604 21242 22660 21244
rect 22684 21242 22740 21244
rect 22364 21190 22366 21242
rect 22366 21190 22418 21242
rect 22418 21190 22420 21242
rect 22444 21190 22482 21242
rect 22482 21190 22494 21242
rect 22494 21190 22500 21242
rect 22524 21190 22546 21242
rect 22546 21190 22558 21242
rect 22558 21190 22580 21242
rect 22604 21190 22610 21242
rect 22610 21190 22622 21242
rect 22622 21190 22660 21242
rect 22684 21190 22686 21242
rect 22686 21190 22738 21242
rect 22738 21190 22740 21242
rect 22364 21188 22420 21190
rect 22444 21188 22500 21190
rect 22524 21188 22580 21190
rect 22604 21188 22660 21190
rect 22684 21188 22740 21190
rect 22190 19896 22246 19952
rect 22374 20340 22376 20360
rect 22376 20340 22428 20360
rect 22428 20340 22430 20360
rect 22374 20304 22430 20340
rect 22364 20154 22420 20156
rect 22444 20154 22500 20156
rect 22524 20154 22580 20156
rect 22604 20154 22660 20156
rect 22684 20154 22740 20156
rect 22364 20102 22366 20154
rect 22366 20102 22418 20154
rect 22418 20102 22420 20154
rect 22444 20102 22482 20154
rect 22482 20102 22494 20154
rect 22494 20102 22500 20154
rect 22524 20102 22546 20154
rect 22546 20102 22558 20154
rect 22558 20102 22580 20154
rect 22604 20102 22610 20154
rect 22610 20102 22622 20154
rect 22622 20102 22660 20154
rect 22684 20102 22686 20154
rect 22686 20102 22738 20154
rect 22738 20102 22740 20154
rect 22364 20100 22420 20102
rect 22444 20100 22500 20102
rect 22524 20100 22580 20102
rect 22604 20100 22660 20102
rect 22684 20100 22740 20102
rect 22364 19066 22420 19068
rect 22444 19066 22500 19068
rect 22524 19066 22580 19068
rect 22604 19066 22660 19068
rect 22684 19066 22740 19068
rect 22364 19014 22366 19066
rect 22366 19014 22418 19066
rect 22418 19014 22420 19066
rect 22444 19014 22482 19066
rect 22482 19014 22494 19066
rect 22494 19014 22500 19066
rect 22524 19014 22546 19066
rect 22546 19014 22558 19066
rect 22558 19014 22580 19066
rect 22604 19014 22610 19066
rect 22610 19014 22622 19066
rect 22622 19014 22660 19066
rect 22684 19014 22686 19066
rect 22686 19014 22738 19066
rect 22738 19014 22740 19066
rect 22364 19012 22420 19014
rect 22444 19012 22500 19014
rect 22524 19012 22580 19014
rect 22604 19012 22660 19014
rect 22684 19012 22740 19014
rect 22006 18536 22062 18592
rect 22364 17978 22420 17980
rect 22444 17978 22500 17980
rect 22524 17978 22580 17980
rect 22604 17978 22660 17980
rect 22684 17978 22740 17980
rect 22364 17926 22366 17978
rect 22366 17926 22418 17978
rect 22418 17926 22420 17978
rect 22444 17926 22482 17978
rect 22482 17926 22494 17978
rect 22494 17926 22500 17978
rect 22524 17926 22546 17978
rect 22546 17926 22558 17978
rect 22558 17926 22580 17978
rect 22604 17926 22610 17978
rect 22610 17926 22622 17978
rect 22622 17926 22660 17978
rect 22684 17926 22686 17978
rect 22686 17926 22738 17978
rect 22738 17926 22740 17978
rect 22364 17924 22420 17926
rect 22444 17924 22500 17926
rect 22524 17924 22580 17926
rect 22604 17924 22660 17926
rect 22684 17924 22740 17926
rect 22364 16890 22420 16892
rect 22444 16890 22500 16892
rect 22524 16890 22580 16892
rect 22604 16890 22660 16892
rect 22684 16890 22740 16892
rect 22364 16838 22366 16890
rect 22366 16838 22418 16890
rect 22418 16838 22420 16890
rect 22444 16838 22482 16890
rect 22482 16838 22494 16890
rect 22494 16838 22500 16890
rect 22524 16838 22546 16890
rect 22546 16838 22558 16890
rect 22558 16838 22580 16890
rect 22604 16838 22610 16890
rect 22610 16838 22622 16890
rect 22622 16838 22660 16890
rect 22684 16838 22686 16890
rect 22686 16838 22738 16890
rect 22738 16838 22740 16890
rect 22364 16836 22420 16838
rect 22444 16836 22500 16838
rect 22524 16836 22580 16838
rect 22604 16836 22660 16838
rect 22684 16836 22740 16838
rect 22364 15802 22420 15804
rect 22444 15802 22500 15804
rect 22524 15802 22580 15804
rect 22604 15802 22660 15804
rect 22684 15802 22740 15804
rect 22364 15750 22366 15802
rect 22366 15750 22418 15802
rect 22418 15750 22420 15802
rect 22444 15750 22482 15802
rect 22482 15750 22494 15802
rect 22494 15750 22500 15802
rect 22524 15750 22546 15802
rect 22546 15750 22558 15802
rect 22558 15750 22580 15802
rect 22604 15750 22610 15802
rect 22610 15750 22622 15802
rect 22622 15750 22660 15802
rect 22684 15750 22686 15802
rect 22686 15750 22738 15802
rect 22738 15750 22740 15802
rect 22364 15748 22420 15750
rect 22444 15748 22500 15750
rect 22524 15748 22580 15750
rect 22604 15748 22660 15750
rect 22684 15748 22740 15750
rect 23202 18672 23258 18728
rect 22364 14714 22420 14716
rect 22444 14714 22500 14716
rect 22524 14714 22580 14716
rect 22604 14714 22660 14716
rect 22684 14714 22740 14716
rect 22364 14662 22366 14714
rect 22366 14662 22418 14714
rect 22418 14662 22420 14714
rect 22444 14662 22482 14714
rect 22482 14662 22494 14714
rect 22494 14662 22500 14714
rect 22524 14662 22546 14714
rect 22546 14662 22558 14714
rect 22558 14662 22580 14714
rect 22604 14662 22610 14714
rect 22610 14662 22622 14714
rect 22622 14662 22660 14714
rect 22684 14662 22686 14714
rect 22686 14662 22738 14714
rect 22738 14662 22740 14714
rect 22364 14660 22420 14662
rect 22444 14660 22500 14662
rect 22524 14660 22580 14662
rect 22604 14660 22660 14662
rect 22684 14660 22740 14662
rect 21086 9596 21088 9616
rect 21088 9596 21140 9616
rect 21140 9596 21142 9616
rect 21086 9560 21142 9596
rect 21730 10240 21786 10296
rect 21454 10104 21510 10160
rect 21086 8472 21142 8528
rect 22364 13626 22420 13628
rect 22444 13626 22500 13628
rect 22524 13626 22580 13628
rect 22604 13626 22660 13628
rect 22684 13626 22740 13628
rect 22364 13574 22366 13626
rect 22366 13574 22418 13626
rect 22418 13574 22420 13626
rect 22444 13574 22482 13626
rect 22482 13574 22494 13626
rect 22494 13574 22500 13626
rect 22524 13574 22546 13626
rect 22546 13574 22558 13626
rect 22558 13574 22580 13626
rect 22604 13574 22610 13626
rect 22610 13574 22622 13626
rect 22622 13574 22660 13626
rect 22684 13574 22686 13626
rect 22686 13574 22738 13626
rect 22738 13574 22740 13626
rect 22364 13572 22420 13574
rect 22444 13572 22500 13574
rect 22524 13572 22580 13574
rect 22604 13572 22660 13574
rect 22684 13572 22740 13574
rect 22364 12538 22420 12540
rect 22444 12538 22500 12540
rect 22524 12538 22580 12540
rect 22604 12538 22660 12540
rect 22684 12538 22740 12540
rect 22364 12486 22366 12538
rect 22366 12486 22418 12538
rect 22418 12486 22420 12538
rect 22444 12486 22482 12538
rect 22482 12486 22494 12538
rect 22494 12486 22500 12538
rect 22524 12486 22546 12538
rect 22546 12486 22558 12538
rect 22558 12486 22580 12538
rect 22604 12486 22610 12538
rect 22610 12486 22622 12538
rect 22622 12486 22660 12538
rect 22684 12486 22686 12538
rect 22686 12486 22738 12538
rect 22738 12486 22740 12538
rect 22364 12484 22420 12486
rect 22444 12484 22500 12486
rect 22524 12484 22580 12486
rect 22604 12484 22660 12486
rect 22684 12484 22740 12486
rect 22364 11450 22420 11452
rect 22444 11450 22500 11452
rect 22524 11450 22580 11452
rect 22604 11450 22660 11452
rect 22684 11450 22740 11452
rect 22364 11398 22366 11450
rect 22366 11398 22418 11450
rect 22418 11398 22420 11450
rect 22444 11398 22482 11450
rect 22482 11398 22494 11450
rect 22494 11398 22500 11450
rect 22524 11398 22546 11450
rect 22546 11398 22558 11450
rect 22558 11398 22580 11450
rect 22604 11398 22610 11450
rect 22610 11398 22622 11450
rect 22622 11398 22660 11450
rect 22684 11398 22686 11450
rect 22686 11398 22738 11450
rect 22738 11398 22740 11450
rect 22364 11396 22420 11398
rect 22444 11396 22500 11398
rect 22524 11396 22580 11398
rect 22604 11396 22660 11398
rect 22684 11396 22740 11398
rect 22364 10362 22420 10364
rect 22444 10362 22500 10364
rect 22524 10362 22580 10364
rect 22604 10362 22660 10364
rect 22684 10362 22740 10364
rect 22364 10310 22366 10362
rect 22366 10310 22418 10362
rect 22418 10310 22420 10362
rect 22444 10310 22482 10362
rect 22482 10310 22494 10362
rect 22494 10310 22500 10362
rect 22524 10310 22546 10362
rect 22546 10310 22558 10362
rect 22558 10310 22580 10362
rect 22604 10310 22610 10362
rect 22610 10310 22622 10362
rect 22622 10310 22660 10362
rect 22684 10310 22686 10362
rect 22686 10310 22738 10362
rect 22738 10310 22740 10362
rect 22364 10308 22420 10310
rect 22444 10308 22500 10310
rect 22524 10308 22580 10310
rect 22604 10308 22660 10310
rect 22684 10308 22740 10310
rect 21454 9036 21510 9072
rect 21454 9016 21456 9036
rect 21456 9016 21508 9036
rect 21508 9016 21510 9036
rect 21546 7384 21602 7440
rect 21362 6160 21418 6216
rect 21086 4140 21142 4176
rect 21086 4120 21088 4140
rect 21088 4120 21140 4140
rect 21140 4120 21142 4140
rect 20350 3032 20406 3088
rect 21086 3576 21142 3632
rect 21178 3440 21234 3496
rect 22364 9274 22420 9276
rect 22444 9274 22500 9276
rect 22524 9274 22580 9276
rect 22604 9274 22660 9276
rect 22684 9274 22740 9276
rect 22364 9222 22366 9274
rect 22366 9222 22418 9274
rect 22418 9222 22420 9274
rect 22444 9222 22482 9274
rect 22482 9222 22494 9274
rect 22494 9222 22500 9274
rect 22524 9222 22546 9274
rect 22546 9222 22558 9274
rect 22558 9222 22580 9274
rect 22604 9222 22610 9274
rect 22610 9222 22622 9274
rect 22622 9222 22660 9274
rect 22684 9222 22686 9274
rect 22686 9222 22738 9274
rect 22738 9222 22740 9274
rect 22364 9220 22420 9222
rect 22444 9220 22500 9222
rect 22524 9220 22580 9222
rect 22604 9220 22660 9222
rect 22684 9220 22740 9222
rect 21914 6840 21970 6896
rect 22834 8336 22890 8392
rect 22364 8186 22420 8188
rect 22444 8186 22500 8188
rect 22524 8186 22580 8188
rect 22604 8186 22660 8188
rect 22684 8186 22740 8188
rect 22364 8134 22366 8186
rect 22366 8134 22418 8186
rect 22418 8134 22420 8186
rect 22444 8134 22482 8186
rect 22482 8134 22494 8186
rect 22494 8134 22500 8186
rect 22524 8134 22546 8186
rect 22546 8134 22558 8186
rect 22558 8134 22580 8186
rect 22604 8134 22610 8186
rect 22610 8134 22622 8186
rect 22622 8134 22660 8186
rect 22684 8134 22686 8186
rect 22686 8134 22738 8186
rect 22738 8134 22740 8186
rect 22364 8132 22420 8134
rect 22444 8132 22500 8134
rect 22524 8132 22580 8134
rect 22604 8132 22660 8134
rect 22684 8132 22740 8134
rect 22364 7098 22420 7100
rect 22444 7098 22500 7100
rect 22524 7098 22580 7100
rect 22604 7098 22660 7100
rect 22684 7098 22740 7100
rect 22364 7046 22366 7098
rect 22366 7046 22418 7098
rect 22418 7046 22420 7098
rect 22444 7046 22482 7098
rect 22482 7046 22494 7098
rect 22494 7046 22500 7098
rect 22524 7046 22546 7098
rect 22546 7046 22558 7098
rect 22558 7046 22580 7098
rect 22604 7046 22610 7098
rect 22610 7046 22622 7098
rect 22622 7046 22660 7098
rect 22684 7046 22686 7098
rect 22686 7046 22738 7098
rect 22738 7046 22740 7098
rect 22364 7044 22420 7046
rect 22444 7044 22500 7046
rect 22524 7044 22580 7046
rect 22604 7044 22660 7046
rect 22684 7044 22740 7046
rect 22098 6840 22154 6896
rect 21914 6568 21970 6624
rect 22364 6010 22420 6012
rect 22444 6010 22500 6012
rect 22524 6010 22580 6012
rect 22604 6010 22660 6012
rect 22684 6010 22740 6012
rect 22364 5958 22366 6010
rect 22366 5958 22418 6010
rect 22418 5958 22420 6010
rect 22444 5958 22482 6010
rect 22482 5958 22494 6010
rect 22494 5958 22500 6010
rect 22524 5958 22546 6010
rect 22546 5958 22558 6010
rect 22558 5958 22580 6010
rect 22604 5958 22610 6010
rect 22610 5958 22622 6010
rect 22622 5958 22660 6010
rect 22684 5958 22686 6010
rect 22686 5958 22738 6010
rect 22738 5958 22740 6010
rect 22364 5956 22420 5958
rect 22444 5956 22500 5958
rect 22524 5956 22580 5958
rect 22604 5956 22660 5958
rect 22684 5956 22740 5958
rect 20442 1808 20498 1864
rect 20350 1672 20406 1728
rect 20166 1264 20222 1320
rect 20626 1300 20628 1320
rect 20628 1300 20680 1320
rect 20680 1300 20682 1320
rect 21822 2624 21878 2680
rect 22364 4922 22420 4924
rect 22444 4922 22500 4924
rect 22524 4922 22580 4924
rect 22604 4922 22660 4924
rect 22684 4922 22740 4924
rect 22364 4870 22366 4922
rect 22366 4870 22418 4922
rect 22418 4870 22420 4922
rect 22444 4870 22482 4922
rect 22482 4870 22494 4922
rect 22494 4870 22500 4922
rect 22524 4870 22546 4922
rect 22546 4870 22558 4922
rect 22558 4870 22580 4922
rect 22604 4870 22610 4922
rect 22610 4870 22622 4922
rect 22622 4870 22660 4922
rect 22684 4870 22686 4922
rect 22686 4870 22738 4922
rect 22738 4870 22740 4922
rect 22364 4868 22420 4870
rect 22444 4868 22500 4870
rect 22524 4868 22580 4870
rect 22604 4868 22660 4870
rect 22684 4868 22740 4870
rect 22364 3834 22420 3836
rect 22444 3834 22500 3836
rect 22524 3834 22580 3836
rect 22604 3834 22660 3836
rect 22684 3834 22740 3836
rect 22364 3782 22366 3834
rect 22366 3782 22418 3834
rect 22418 3782 22420 3834
rect 22444 3782 22482 3834
rect 22482 3782 22494 3834
rect 22494 3782 22500 3834
rect 22524 3782 22546 3834
rect 22546 3782 22558 3834
rect 22558 3782 22580 3834
rect 22604 3782 22610 3834
rect 22610 3782 22622 3834
rect 22622 3782 22660 3834
rect 22684 3782 22686 3834
rect 22686 3782 22738 3834
rect 22738 3782 22740 3834
rect 22364 3780 22420 3782
rect 22444 3780 22500 3782
rect 22524 3780 22580 3782
rect 22604 3780 22660 3782
rect 22684 3780 22740 3782
rect 22190 2352 22246 2408
rect 20626 1264 20682 1300
rect 20442 1164 20444 1184
rect 20444 1164 20496 1184
rect 20496 1164 20498 1184
rect 20442 1128 20498 1164
rect 20718 992 20774 1048
rect 20626 448 20682 504
rect 21638 856 21694 912
rect 21822 448 21878 504
rect 22364 2746 22420 2748
rect 22444 2746 22500 2748
rect 22524 2746 22580 2748
rect 22604 2746 22660 2748
rect 22684 2746 22740 2748
rect 22364 2694 22366 2746
rect 22366 2694 22418 2746
rect 22418 2694 22420 2746
rect 22444 2694 22482 2746
rect 22482 2694 22494 2746
rect 22494 2694 22500 2746
rect 22524 2694 22546 2746
rect 22546 2694 22558 2746
rect 22558 2694 22580 2746
rect 22604 2694 22610 2746
rect 22610 2694 22622 2746
rect 22622 2694 22660 2746
rect 22684 2694 22686 2746
rect 22686 2694 22738 2746
rect 22738 2694 22740 2746
rect 22364 2692 22420 2694
rect 22444 2692 22500 2694
rect 22524 2692 22580 2694
rect 22604 2692 22660 2694
rect 22684 2692 22740 2694
rect 22466 2216 22522 2272
rect 22558 1844 22560 1864
rect 22560 1844 22612 1864
rect 22612 1844 22614 1864
rect 22558 1808 22614 1844
rect 22364 1658 22420 1660
rect 22444 1658 22500 1660
rect 22524 1658 22580 1660
rect 22604 1658 22660 1660
rect 22684 1658 22740 1660
rect 22364 1606 22366 1658
rect 22366 1606 22418 1658
rect 22418 1606 22420 1658
rect 22444 1606 22482 1658
rect 22482 1606 22494 1658
rect 22494 1606 22500 1658
rect 22524 1606 22546 1658
rect 22546 1606 22558 1658
rect 22558 1606 22580 1658
rect 22604 1606 22610 1658
rect 22610 1606 22622 1658
rect 22622 1606 22660 1658
rect 22684 1606 22686 1658
rect 22686 1606 22738 1658
rect 22738 1606 22740 1658
rect 22364 1604 22420 1606
rect 22444 1604 22500 1606
rect 22524 1604 22580 1606
rect 22604 1604 22660 1606
rect 22684 1604 22740 1606
rect 22364 570 22420 572
rect 22444 570 22500 572
rect 22524 570 22580 572
rect 22604 570 22660 572
rect 22684 570 22740 572
rect 22364 518 22366 570
rect 22366 518 22418 570
rect 22418 518 22420 570
rect 22444 518 22482 570
rect 22482 518 22494 570
rect 22494 518 22500 570
rect 22524 518 22546 570
rect 22546 518 22558 570
rect 22558 518 22580 570
rect 22604 518 22610 570
rect 22610 518 22622 570
rect 22622 518 22660 570
rect 22684 518 22686 570
rect 22686 518 22738 570
rect 22738 518 22740 570
rect 22364 516 22420 518
rect 22444 516 22500 518
rect 22524 516 22580 518
rect 22604 516 22660 518
rect 22684 516 22740 518
<< metal3 >>
rect 4354 23424 4750 23425
rect 4354 23360 4360 23424
rect 4424 23360 4440 23424
rect 4504 23360 4520 23424
rect 4584 23360 4600 23424
rect 4664 23360 4680 23424
rect 4744 23360 4750 23424
rect 4354 23359 4750 23360
rect 10354 23424 10750 23425
rect 10354 23360 10360 23424
rect 10424 23360 10440 23424
rect 10504 23360 10520 23424
rect 10584 23360 10600 23424
rect 10664 23360 10680 23424
rect 10744 23360 10750 23424
rect 10354 23359 10750 23360
rect 16354 23424 16750 23425
rect 16354 23360 16360 23424
rect 16424 23360 16440 23424
rect 16504 23360 16520 23424
rect 16584 23360 16600 23424
rect 16664 23360 16680 23424
rect 16744 23360 16750 23424
rect 16354 23359 16750 23360
rect 22354 23424 22750 23425
rect 22354 23360 22360 23424
rect 22424 23360 22440 23424
rect 22504 23360 22520 23424
rect 22584 23360 22600 23424
rect 22664 23360 22680 23424
rect 22744 23360 22750 23424
rect 22354 23359 22750 23360
rect 21633 22948 21699 22949
rect 21582 22884 21588 22948
rect 21652 22946 21699 22948
rect 21652 22944 21744 22946
rect 21694 22888 21744 22944
rect 21652 22886 21744 22888
rect 21652 22884 21699 22886
rect 21633 22883 21699 22884
rect 1354 22880 1750 22881
rect 1354 22816 1360 22880
rect 1424 22816 1440 22880
rect 1504 22816 1520 22880
rect 1584 22816 1600 22880
rect 1664 22816 1680 22880
rect 1744 22816 1750 22880
rect 1354 22815 1750 22816
rect 7354 22880 7750 22881
rect 7354 22816 7360 22880
rect 7424 22816 7440 22880
rect 7504 22816 7520 22880
rect 7584 22816 7600 22880
rect 7664 22816 7680 22880
rect 7744 22816 7750 22880
rect 7354 22815 7750 22816
rect 13354 22880 13750 22881
rect 13354 22816 13360 22880
rect 13424 22816 13440 22880
rect 13504 22816 13520 22880
rect 13584 22816 13600 22880
rect 13664 22816 13680 22880
rect 13744 22816 13750 22880
rect 13354 22815 13750 22816
rect 19354 22880 19750 22881
rect 19354 22816 19360 22880
rect 19424 22816 19440 22880
rect 19504 22816 19520 22880
rect 19584 22816 19600 22880
rect 19664 22816 19680 22880
rect 19744 22816 19750 22880
rect 19354 22815 19750 22816
rect 10777 22674 10843 22677
rect 11646 22674 11652 22676
rect 10777 22672 11652 22674
rect 10777 22616 10782 22672
rect 10838 22616 11652 22672
rect 10777 22614 11652 22616
rect 10777 22611 10843 22614
rect 11646 22612 11652 22614
rect 11716 22612 11722 22676
rect 10041 22540 10107 22541
rect 9990 22538 9996 22540
rect 9950 22478 9996 22538
rect 10060 22536 10107 22540
rect 10102 22480 10107 22536
rect 9990 22476 9996 22478
rect 10060 22476 10107 22480
rect 10041 22475 10107 22476
rect 2957 22402 3023 22405
rect 3182 22402 3188 22404
rect 2957 22400 3188 22402
rect 2957 22344 2962 22400
rect 3018 22344 3188 22400
rect 2957 22342 3188 22344
rect 2957 22339 3023 22342
rect 3182 22340 3188 22342
rect 3252 22340 3258 22404
rect 6494 22340 6500 22404
rect 6564 22402 6570 22404
rect 9673 22402 9739 22405
rect 6564 22400 9739 22402
rect 6564 22344 9678 22400
rect 9734 22344 9739 22400
rect 6564 22342 9739 22344
rect 6564 22340 6570 22342
rect 9673 22339 9739 22342
rect 4354 22336 4750 22337
rect 4354 22272 4360 22336
rect 4424 22272 4440 22336
rect 4504 22272 4520 22336
rect 4584 22272 4600 22336
rect 4664 22272 4680 22336
rect 4744 22272 4750 22336
rect 4354 22271 4750 22272
rect 10354 22336 10750 22337
rect 10354 22272 10360 22336
rect 10424 22272 10440 22336
rect 10504 22272 10520 22336
rect 10584 22272 10600 22336
rect 10664 22272 10680 22336
rect 10744 22272 10750 22336
rect 10354 22271 10750 22272
rect 16354 22336 16750 22337
rect 16354 22272 16360 22336
rect 16424 22272 16440 22336
rect 16504 22272 16520 22336
rect 16584 22272 16600 22336
rect 16664 22272 16680 22336
rect 16744 22272 16750 22336
rect 16354 22271 16750 22272
rect 22354 22336 22750 22337
rect 22354 22272 22360 22336
rect 22424 22272 22440 22336
rect 22504 22272 22520 22336
rect 22584 22272 22600 22336
rect 22664 22272 22680 22336
rect 22744 22272 22750 22336
rect 22354 22271 22750 22272
rect 21081 22266 21147 22269
rect 21214 22266 21220 22268
rect 21081 22264 21220 22266
rect 21081 22208 21086 22264
rect 21142 22208 21220 22264
rect 21081 22206 21220 22208
rect 21081 22203 21147 22206
rect 21214 22204 21220 22206
rect 21284 22204 21290 22268
rect 3918 22068 3924 22132
rect 3988 22130 3994 22132
rect 5349 22130 5415 22133
rect 3988 22128 5415 22130
rect 3988 22072 5354 22128
rect 5410 22072 5415 22128
rect 3988 22070 5415 22072
rect 3988 22068 3994 22070
rect 5349 22067 5415 22070
rect 15101 22130 15167 22133
rect 19241 22130 19307 22133
rect 15101 22128 19307 22130
rect 15101 22072 15106 22128
rect 15162 22072 19246 22128
rect 19302 22072 19307 22128
rect 15101 22070 19307 22072
rect 15101 22067 15167 22070
rect 19241 22067 19307 22070
rect 8017 21994 8083 21997
rect 9397 21994 9463 21997
rect 8017 21992 9463 21994
rect 8017 21936 8022 21992
rect 8078 21936 9402 21992
rect 9458 21936 9463 21992
rect 8017 21934 9463 21936
rect 8017 21931 8083 21934
rect 9397 21931 9463 21934
rect 13169 21994 13235 21997
rect 19333 21994 19399 21997
rect 13169 21992 19399 21994
rect 13169 21936 13174 21992
rect 13230 21936 19338 21992
rect 19394 21936 19399 21992
rect 13169 21934 19399 21936
rect 13169 21931 13235 21934
rect 19333 21931 19399 21934
rect 9806 21796 9812 21860
rect 9876 21858 9882 21860
rect 12525 21858 12591 21861
rect 9876 21856 12591 21858
rect 9876 21800 12530 21856
rect 12586 21800 12591 21856
rect 9876 21798 12591 21800
rect 9876 21796 9882 21798
rect 12525 21795 12591 21798
rect 13813 21858 13879 21861
rect 14406 21858 14412 21860
rect 13813 21856 14412 21858
rect 13813 21800 13818 21856
rect 13874 21800 14412 21856
rect 13813 21798 14412 21800
rect 13813 21795 13879 21798
rect 14406 21796 14412 21798
rect 14476 21796 14482 21860
rect 1354 21792 1750 21793
rect 1354 21728 1360 21792
rect 1424 21728 1440 21792
rect 1504 21728 1520 21792
rect 1584 21728 1600 21792
rect 1664 21728 1680 21792
rect 1744 21728 1750 21792
rect 1354 21727 1750 21728
rect 7354 21792 7750 21793
rect 7354 21728 7360 21792
rect 7424 21728 7440 21792
rect 7504 21728 7520 21792
rect 7584 21728 7600 21792
rect 7664 21728 7680 21792
rect 7744 21728 7750 21792
rect 7354 21727 7750 21728
rect 13354 21792 13750 21793
rect 13354 21728 13360 21792
rect 13424 21728 13440 21792
rect 13504 21728 13520 21792
rect 13584 21728 13600 21792
rect 13664 21728 13680 21792
rect 13744 21728 13750 21792
rect 13354 21727 13750 21728
rect 19354 21792 19750 21793
rect 19354 21728 19360 21792
rect 19424 21728 19440 21792
rect 19504 21728 19520 21792
rect 19584 21728 19600 21792
rect 19664 21728 19680 21792
rect 19744 21728 19750 21792
rect 19354 21727 19750 21728
rect 16113 21722 16179 21725
rect 17953 21722 18019 21725
rect 16113 21720 18019 21722
rect 16113 21664 16118 21720
rect 16174 21664 17958 21720
rect 18014 21664 18019 21720
rect 16113 21662 18019 21664
rect 16113 21659 16179 21662
rect 17953 21659 18019 21662
rect 19977 21722 20043 21725
rect 21449 21722 21515 21725
rect 19977 21720 21515 21722
rect 19977 21664 19982 21720
rect 20038 21664 21454 21720
rect 21510 21664 21515 21720
rect 19977 21662 21515 21664
rect 19977 21659 20043 21662
rect 21449 21659 21515 21662
rect 3877 21586 3943 21589
rect 8569 21586 8635 21589
rect 3877 21584 8635 21586
rect 3877 21528 3882 21584
rect 3938 21528 8574 21584
rect 8630 21528 8635 21584
rect 3877 21526 8635 21528
rect 3877 21523 3943 21526
rect 8569 21523 8635 21526
rect 11145 21586 11211 21589
rect 15929 21586 15995 21589
rect 20069 21586 20135 21589
rect 11145 21584 20135 21586
rect 11145 21528 11150 21584
rect 11206 21528 15934 21584
rect 15990 21528 20074 21584
rect 20130 21528 20135 21584
rect 11145 21526 20135 21528
rect 11145 21523 11211 21526
rect 15929 21523 15995 21526
rect 20069 21523 20135 21526
rect 2773 21450 2839 21453
rect 10041 21450 10107 21453
rect 2773 21448 10107 21450
rect 2773 21392 2778 21448
rect 2834 21392 10046 21448
rect 10102 21392 10107 21448
rect 2773 21390 10107 21392
rect 2773 21387 2839 21390
rect 10041 21387 10107 21390
rect 13905 21450 13971 21453
rect 21541 21450 21607 21453
rect 21817 21450 21883 21453
rect 13905 21448 21883 21450
rect 13905 21392 13910 21448
rect 13966 21392 21546 21448
rect 21602 21392 21822 21448
rect 21878 21392 21883 21448
rect 13905 21390 21883 21392
rect 13905 21387 13971 21390
rect 21541 21387 21607 21390
rect 21817 21387 21883 21390
rect 7097 21314 7163 21317
rect 8753 21314 8819 21317
rect 7097 21312 8819 21314
rect 7097 21256 7102 21312
rect 7158 21256 8758 21312
rect 8814 21256 8819 21312
rect 7097 21254 8819 21256
rect 7097 21251 7163 21254
rect 8753 21251 8819 21254
rect 20069 21314 20135 21317
rect 21449 21314 21515 21317
rect 20069 21312 21515 21314
rect 20069 21256 20074 21312
rect 20130 21256 21454 21312
rect 21510 21256 21515 21312
rect 20069 21254 21515 21256
rect 20069 21251 20135 21254
rect 21449 21251 21515 21254
rect 4354 21248 4750 21249
rect 4354 21184 4360 21248
rect 4424 21184 4440 21248
rect 4504 21184 4520 21248
rect 4584 21184 4600 21248
rect 4664 21184 4680 21248
rect 4744 21184 4750 21248
rect 4354 21183 4750 21184
rect 10354 21248 10750 21249
rect 10354 21184 10360 21248
rect 10424 21184 10440 21248
rect 10504 21184 10520 21248
rect 10584 21184 10600 21248
rect 10664 21184 10680 21248
rect 10744 21184 10750 21248
rect 10354 21183 10750 21184
rect 16354 21248 16750 21249
rect 16354 21184 16360 21248
rect 16424 21184 16440 21248
rect 16504 21184 16520 21248
rect 16584 21184 16600 21248
rect 16664 21184 16680 21248
rect 16744 21184 16750 21248
rect 16354 21183 16750 21184
rect 22354 21248 22750 21249
rect 22354 21184 22360 21248
rect 22424 21184 22440 21248
rect 22504 21184 22520 21248
rect 22584 21184 22600 21248
rect 22664 21184 22680 21248
rect 22744 21184 22750 21248
rect 22354 21183 22750 21184
rect 4981 21178 5047 21181
rect 8937 21178 9003 21181
rect 4981 21176 9003 21178
rect 4981 21120 4986 21176
rect 5042 21120 8942 21176
rect 8998 21120 9003 21176
rect 4981 21118 9003 21120
rect 4981 21115 5047 21118
rect 8937 21115 9003 21118
rect 3509 21042 3575 21045
rect 6085 21042 6151 21045
rect 7373 21042 7439 21045
rect 3509 21040 7439 21042
rect 3509 20984 3514 21040
rect 3570 20984 6090 21040
rect 6146 20984 7378 21040
rect 7434 20984 7439 21040
rect 3509 20982 7439 20984
rect 3509 20979 3575 20982
rect 6085 20979 6151 20982
rect 7373 20979 7439 20982
rect 9029 21042 9095 21045
rect 18873 21042 18939 21045
rect 9029 21040 18939 21042
rect 9029 20984 9034 21040
rect 9090 20984 18878 21040
rect 18934 20984 18939 21040
rect 9029 20982 18939 20984
rect 9029 20979 9095 20982
rect 18873 20979 18939 20982
rect 4061 20906 4127 20909
rect 4705 20906 4771 20909
rect 4061 20904 4771 20906
rect 4061 20848 4066 20904
rect 4122 20848 4710 20904
rect 4766 20848 4771 20904
rect 4061 20846 4771 20848
rect 4061 20843 4127 20846
rect 4705 20843 4771 20846
rect 6269 20906 6335 20909
rect 9857 20906 9923 20909
rect 6269 20904 9923 20906
rect 6269 20848 6274 20904
rect 6330 20848 9862 20904
rect 9918 20848 9923 20904
rect 6269 20846 9923 20848
rect 6269 20843 6335 20846
rect 9857 20843 9923 20846
rect 11513 20906 11579 20909
rect 12617 20906 12683 20909
rect 15101 20906 15167 20909
rect 19425 20906 19491 20909
rect 11513 20904 12683 20906
rect 11513 20848 11518 20904
rect 11574 20848 12622 20904
rect 12678 20848 12683 20904
rect 11513 20846 12683 20848
rect 11513 20843 11579 20846
rect 12617 20843 12683 20846
rect 13172 20904 15167 20906
rect 13172 20848 15106 20904
rect 15162 20848 15167 20904
rect 13172 20846 15167 20848
rect 6545 20770 6611 20773
rect 6678 20770 6684 20772
rect 6545 20768 6684 20770
rect 6545 20712 6550 20768
rect 6606 20712 6684 20768
rect 6545 20710 6684 20712
rect 6545 20707 6611 20710
rect 6678 20708 6684 20710
rect 6748 20708 6754 20772
rect 8753 20770 8819 20773
rect 9581 20770 9647 20773
rect 12525 20770 12591 20773
rect 12801 20772 12867 20773
rect 8753 20768 12591 20770
rect 8753 20712 8758 20768
rect 8814 20712 9586 20768
rect 9642 20712 12530 20768
rect 12586 20712 12591 20768
rect 8753 20710 12591 20712
rect 8753 20707 8819 20710
rect 9581 20707 9647 20710
rect 12525 20707 12591 20710
rect 12750 20708 12756 20772
rect 12820 20770 12867 20772
rect 12820 20768 12912 20770
rect 12862 20712 12912 20768
rect 12820 20710 12912 20712
rect 12820 20708 12867 20710
rect 12801 20707 12867 20708
rect 1354 20704 1750 20705
rect 1354 20640 1360 20704
rect 1424 20640 1440 20704
rect 1504 20640 1520 20704
rect 1584 20640 1600 20704
rect 1664 20640 1680 20704
rect 1744 20640 1750 20704
rect 1354 20639 1750 20640
rect 7354 20704 7750 20705
rect 7354 20640 7360 20704
rect 7424 20640 7440 20704
rect 7504 20640 7520 20704
rect 7584 20640 7600 20704
rect 7664 20640 7680 20704
rect 7744 20640 7750 20704
rect 7354 20639 7750 20640
rect 9949 20634 10015 20637
rect 13172 20634 13232 20846
rect 15101 20843 15167 20846
rect 17910 20904 19491 20906
rect 17910 20848 19430 20904
rect 19486 20848 19491 20904
rect 17910 20846 19491 20848
rect 13354 20704 13750 20705
rect 13354 20640 13360 20704
rect 13424 20640 13440 20704
rect 13504 20640 13520 20704
rect 13584 20640 13600 20704
rect 13664 20640 13680 20704
rect 13744 20640 13750 20704
rect 13354 20639 13750 20640
rect 17217 20634 17283 20637
rect 17910 20634 17970 20846
rect 19425 20843 19491 20846
rect 20713 20906 20779 20909
rect 21030 20906 21036 20908
rect 20713 20904 21036 20906
rect 20713 20848 20718 20904
rect 20774 20848 21036 20904
rect 20713 20846 21036 20848
rect 20713 20843 20779 20846
rect 21030 20844 21036 20846
rect 21100 20844 21106 20908
rect 19354 20704 19750 20705
rect 19354 20640 19360 20704
rect 19424 20640 19440 20704
rect 19504 20640 19520 20704
rect 19584 20640 19600 20704
rect 19664 20640 19680 20704
rect 19744 20640 19750 20704
rect 19354 20639 19750 20640
rect 9949 20632 13232 20634
rect 9949 20576 9954 20632
rect 10010 20576 13232 20632
rect 9949 20574 13232 20576
rect 16070 20632 17970 20634
rect 16070 20576 17222 20632
rect 17278 20576 17970 20632
rect 16070 20574 17970 20576
rect 9949 20571 10015 20574
rect 2129 20498 2195 20501
rect 11421 20498 11487 20501
rect 16070 20498 16130 20574
rect 17217 20571 17283 20574
rect 2129 20496 11487 20498
rect 2129 20440 2134 20496
rect 2190 20440 11426 20496
rect 11482 20440 11487 20496
rect 2129 20438 11487 20440
rect 2129 20435 2195 20438
rect 11421 20435 11487 20438
rect 12390 20438 16130 20498
rect 16205 20498 16271 20501
rect 20805 20498 20871 20501
rect 16205 20496 20871 20498
rect 16205 20440 16210 20496
rect 16266 20440 20810 20496
rect 20866 20440 20871 20496
rect 16205 20438 20871 20440
rect 2037 20362 2103 20365
rect 12390 20362 12450 20438
rect 16205 20435 16271 20438
rect 20805 20435 20871 20438
rect 16849 20362 16915 20365
rect 2037 20360 12450 20362
rect 2037 20304 2042 20360
rect 2098 20304 12450 20360
rect 2037 20302 12450 20304
rect 14598 20360 16915 20362
rect 14598 20304 16854 20360
rect 16910 20304 16915 20360
rect 14598 20302 16915 20304
rect 2037 20299 2103 20302
rect 6913 20226 6979 20229
rect 8569 20226 8635 20229
rect 6913 20224 8635 20226
rect 6913 20168 6918 20224
rect 6974 20168 8574 20224
rect 8630 20168 8635 20224
rect 6913 20166 8635 20168
rect 6913 20163 6979 20166
rect 8569 20163 8635 20166
rect 10961 20226 11027 20229
rect 14598 20226 14658 20302
rect 16849 20299 16915 20302
rect 19885 20362 19951 20365
rect 20621 20362 20687 20365
rect 22369 20362 22435 20365
rect 19885 20360 22435 20362
rect 19885 20304 19890 20360
rect 19946 20304 20626 20360
rect 20682 20304 22374 20360
rect 22430 20304 22435 20360
rect 19885 20302 22435 20304
rect 19885 20299 19951 20302
rect 20621 20299 20687 20302
rect 22369 20299 22435 20302
rect 10961 20224 14658 20226
rect 10961 20168 10966 20224
rect 11022 20168 14658 20224
rect 10961 20166 14658 20168
rect 10961 20163 11027 20166
rect 4354 20160 4750 20161
rect 4354 20096 4360 20160
rect 4424 20096 4440 20160
rect 4504 20096 4520 20160
rect 4584 20096 4600 20160
rect 4664 20096 4680 20160
rect 4744 20096 4750 20160
rect 4354 20095 4750 20096
rect 10354 20160 10750 20161
rect 10354 20096 10360 20160
rect 10424 20096 10440 20160
rect 10504 20096 10520 20160
rect 10584 20096 10600 20160
rect 10664 20096 10680 20160
rect 10744 20096 10750 20160
rect 10354 20095 10750 20096
rect 16354 20160 16750 20161
rect 16354 20096 16360 20160
rect 16424 20096 16440 20160
rect 16504 20096 16520 20160
rect 16584 20096 16600 20160
rect 16664 20096 16680 20160
rect 16744 20096 16750 20160
rect 16354 20095 16750 20096
rect 22354 20160 22750 20161
rect 22354 20096 22360 20160
rect 22424 20096 22440 20160
rect 22504 20096 22520 20160
rect 22584 20096 22600 20160
rect 22664 20096 22680 20160
rect 22744 20096 22750 20160
rect 22354 20095 22750 20096
rect 6545 20090 6611 20093
rect 8201 20090 8267 20093
rect 6545 20088 8770 20090
rect 6545 20032 6550 20088
rect 6606 20032 8206 20088
rect 8262 20032 8770 20088
rect 6545 20030 8770 20032
rect 6545 20027 6611 20030
rect 8201 20027 8267 20030
rect 5441 19954 5507 19957
rect 8017 19954 8083 19957
rect 5441 19952 8083 19954
rect 5441 19896 5446 19952
rect 5502 19896 8022 19952
rect 8078 19896 8083 19952
rect 5441 19894 8083 19896
rect 8710 19954 8770 20030
rect 18597 19954 18663 19957
rect 8710 19952 18663 19954
rect 8710 19896 18602 19952
rect 18658 19896 18663 19952
rect 8710 19894 18663 19896
rect 5441 19891 5507 19894
rect 8017 19891 8083 19894
rect 18597 19891 18663 19894
rect 20621 19954 20687 19957
rect 22185 19954 22251 19957
rect 20621 19952 22251 19954
rect 20621 19896 20626 19952
rect 20682 19896 22190 19952
rect 22246 19896 22251 19952
rect 20621 19894 22251 19896
rect 20621 19891 20687 19894
rect 22185 19891 22251 19894
rect 7373 19818 7439 19821
rect 7925 19818 7991 19821
rect 17309 19818 17375 19821
rect 20805 19818 20871 19821
rect 21357 19818 21423 19821
rect 7373 19816 21423 19818
rect 7373 19760 7378 19816
rect 7434 19760 7930 19816
rect 7986 19760 17314 19816
rect 17370 19760 20810 19816
rect 20866 19760 21362 19816
rect 21418 19760 21423 19816
rect 7373 19758 21423 19760
rect 7373 19755 7439 19758
rect 7925 19755 7991 19758
rect 17309 19755 17375 19758
rect 20805 19755 20871 19758
rect 21357 19755 21423 19758
rect 10501 19682 10567 19685
rect 9676 19680 10567 19682
rect 9676 19624 10506 19680
rect 10562 19624 10567 19680
rect 9676 19622 10567 19624
rect 1354 19616 1750 19617
rect 1354 19552 1360 19616
rect 1424 19552 1440 19616
rect 1504 19552 1520 19616
rect 1584 19552 1600 19616
rect 1664 19552 1680 19616
rect 1744 19552 1750 19616
rect 1354 19551 1750 19552
rect 7354 19616 7750 19617
rect 7354 19552 7360 19616
rect 7424 19552 7440 19616
rect 7504 19552 7520 19616
rect 7584 19552 7600 19616
rect 7664 19552 7680 19616
rect 7744 19552 7750 19616
rect 7354 19551 7750 19552
rect 9676 19549 9736 19622
rect 10501 19619 10567 19622
rect 18689 19682 18755 19685
rect 18822 19682 18828 19684
rect 18689 19680 18828 19682
rect 18689 19624 18694 19680
rect 18750 19624 18828 19680
rect 18689 19622 18828 19624
rect 18689 19619 18755 19622
rect 18822 19620 18828 19622
rect 18892 19620 18898 19684
rect 20069 19682 20135 19685
rect 20621 19682 20687 19685
rect 20069 19680 20687 19682
rect 20069 19624 20074 19680
rect 20130 19624 20626 19680
rect 20682 19624 20687 19680
rect 20069 19622 20687 19624
rect 20069 19619 20135 19622
rect 20621 19619 20687 19622
rect 13354 19616 13750 19617
rect 13354 19552 13360 19616
rect 13424 19552 13440 19616
rect 13504 19552 13520 19616
rect 13584 19552 13600 19616
rect 13664 19552 13680 19616
rect 13744 19552 13750 19616
rect 13354 19551 13750 19552
rect 19354 19616 19750 19617
rect 19354 19552 19360 19616
rect 19424 19552 19440 19616
rect 19504 19552 19520 19616
rect 19584 19552 19600 19616
rect 19664 19552 19680 19616
rect 19744 19552 19750 19616
rect 19354 19551 19750 19552
rect 9673 19544 9739 19549
rect 9673 19488 9678 19544
rect 9734 19488 9739 19544
rect 9673 19483 9739 19488
rect 3417 19410 3483 19413
rect 16297 19410 16363 19413
rect 3417 19408 16363 19410
rect 3417 19352 3422 19408
rect 3478 19352 16302 19408
rect 16358 19352 16363 19408
rect 3417 19350 16363 19352
rect 3417 19347 3483 19350
rect 16297 19347 16363 19350
rect 18965 19412 19031 19413
rect 18965 19408 19012 19412
rect 19076 19410 19082 19412
rect 21265 19410 21331 19413
rect 22001 19410 22067 19413
rect 18965 19352 18970 19408
rect 18965 19348 19012 19352
rect 19076 19350 19122 19410
rect 21265 19408 22067 19410
rect 21265 19352 21270 19408
rect 21326 19352 22006 19408
rect 22062 19352 22067 19408
rect 21265 19350 22067 19352
rect 19076 19348 19082 19350
rect 18965 19347 19031 19348
rect 21265 19347 21331 19350
rect 22001 19347 22067 19350
rect 1945 19274 2011 19277
rect 4061 19274 4127 19277
rect 1945 19272 4127 19274
rect 1945 19216 1950 19272
rect 2006 19216 4066 19272
rect 4122 19216 4127 19272
rect 1945 19214 4127 19216
rect 1945 19211 2011 19214
rect 4061 19211 4127 19214
rect 6913 19274 6979 19277
rect 8661 19274 8727 19277
rect 6913 19272 8727 19274
rect 6913 19216 6918 19272
rect 6974 19216 8666 19272
rect 8722 19216 8727 19272
rect 6913 19214 8727 19216
rect 6913 19211 6979 19214
rect 8661 19211 8727 19214
rect 9121 19274 9187 19277
rect 15694 19274 15700 19276
rect 9121 19272 15700 19274
rect 9121 19216 9126 19272
rect 9182 19216 15700 19272
rect 9121 19214 15700 19216
rect 9121 19211 9187 19214
rect 15694 19212 15700 19214
rect 15764 19212 15770 19276
rect 20621 19274 20687 19277
rect 21214 19274 21220 19276
rect 20621 19272 21220 19274
rect 20621 19216 20626 19272
rect 20682 19216 21220 19272
rect 20621 19214 21220 19216
rect 20621 19211 20687 19214
rect 21214 19212 21220 19214
rect 21284 19212 21290 19276
rect 2221 19138 2287 19141
rect 3785 19138 3851 19141
rect 2221 19136 3851 19138
rect 2221 19080 2226 19136
rect 2282 19080 3790 19136
rect 3846 19080 3851 19136
rect 2221 19078 3851 19080
rect 2221 19075 2287 19078
rect 3785 19075 3851 19078
rect 6821 19138 6887 19141
rect 9213 19138 9279 19141
rect 6821 19136 9279 19138
rect 6821 19080 6826 19136
rect 6882 19080 9218 19136
rect 9274 19080 9279 19136
rect 6821 19078 9279 19080
rect 6821 19075 6887 19078
rect 9213 19075 9279 19078
rect 9857 19138 9923 19141
rect 10174 19138 10180 19140
rect 9857 19136 10180 19138
rect 9857 19080 9862 19136
rect 9918 19080 10180 19136
rect 9857 19078 10180 19080
rect 9857 19075 9923 19078
rect 10174 19076 10180 19078
rect 10244 19076 10250 19140
rect 4354 19072 4750 19073
rect 4354 19008 4360 19072
rect 4424 19008 4440 19072
rect 4504 19008 4520 19072
rect 4584 19008 4600 19072
rect 4664 19008 4680 19072
rect 4744 19008 4750 19072
rect 4354 19007 4750 19008
rect 10354 19072 10750 19073
rect 10354 19008 10360 19072
rect 10424 19008 10440 19072
rect 10504 19008 10520 19072
rect 10584 19008 10600 19072
rect 10664 19008 10680 19072
rect 10744 19008 10750 19072
rect 10354 19007 10750 19008
rect 16354 19072 16750 19073
rect 16354 19008 16360 19072
rect 16424 19008 16440 19072
rect 16504 19008 16520 19072
rect 16584 19008 16600 19072
rect 16664 19008 16680 19072
rect 16744 19008 16750 19072
rect 16354 19007 16750 19008
rect 22354 19072 22750 19073
rect 22354 19008 22360 19072
rect 22424 19008 22440 19072
rect 22504 19008 22520 19072
rect 22584 19008 22600 19072
rect 22664 19008 22680 19072
rect 22744 19008 22750 19072
rect 22354 19007 22750 19008
rect 13261 18730 13327 18733
rect 23197 18730 23263 18733
rect 13261 18728 23263 18730
rect 13261 18672 13266 18728
rect 13322 18672 23202 18728
rect 23258 18672 23263 18728
rect 13261 18670 23263 18672
rect 13261 18667 13327 18670
rect 23197 18667 23263 18670
rect 5717 18594 5783 18597
rect 7005 18594 7071 18597
rect 5717 18592 7071 18594
rect 5717 18536 5722 18592
rect 5778 18536 7010 18592
rect 7066 18536 7071 18592
rect 5717 18534 7071 18536
rect 5717 18531 5783 18534
rect 7005 18531 7071 18534
rect 19885 18596 19951 18597
rect 19885 18592 19932 18596
rect 19996 18594 20002 18596
rect 21817 18594 21883 18597
rect 22001 18594 22067 18597
rect 19885 18536 19890 18592
rect 19885 18532 19932 18536
rect 19996 18534 20042 18594
rect 21817 18592 22067 18594
rect 21817 18536 21822 18592
rect 21878 18536 22006 18592
rect 22062 18536 22067 18592
rect 21817 18534 22067 18536
rect 19996 18532 20002 18534
rect 19885 18531 19951 18532
rect 21817 18531 21883 18534
rect 22001 18531 22067 18534
rect 1354 18528 1750 18529
rect 1354 18464 1360 18528
rect 1424 18464 1440 18528
rect 1504 18464 1520 18528
rect 1584 18464 1600 18528
rect 1664 18464 1680 18528
rect 1744 18464 1750 18528
rect 1354 18463 1750 18464
rect 7354 18528 7750 18529
rect 7354 18464 7360 18528
rect 7424 18464 7440 18528
rect 7504 18464 7520 18528
rect 7584 18464 7600 18528
rect 7664 18464 7680 18528
rect 7744 18464 7750 18528
rect 7354 18463 7750 18464
rect 13354 18528 13750 18529
rect 13354 18464 13360 18528
rect 13424 18464 13440 18528
rect 13504 18464 13520 18528
rect 13584 18464 13600 18528
rect 13664 18464 13680 18528
rect 13744 18464 13750 18528
rect 13354 18463 13750 18464
rect 19354 18528 19750 18529
rect 19354 18464 19360 18528
rect 19424 18464 19440 18528
rect 19504 18464 19520 18528
rect 19584 18464 19600 18528
rect 19664 18464 19680 18528
rect 19744 18464 19750 18528
rect 19354 18463 19750 18464
rect 5073 18322 5139 18325
rect 9305 18322 9371 18325
rect 10225 18322 10291 18325
rect 5073 18320 10291 18322
rect 5073 18264 5078 18320
rect 5134 18264 9310 18320
rect 9366 18264 10230 18320
rect 10286 18264 10291 18320
rect 5073 18262 10291 18264
rect 5073 18259 5139 18262
rect 9305 18259 9371 18262
rect 10225 18259 10291 18262
rect 4061 18186 4127 18189
rect 9305 18186 9371 18189
rect 4061 18184 9371 18186
rect 4061 18128 4066 18184
rect 4122 18128 9310 18184
rect 9366 18128 9371 18184
rect 4061 18126 9371 18128
rect 4061 18123 4127 18126
rect 9305 18123 9371 18126
rect 9438 18124 9444 18188
rect 9508 18186 9514 18188
rect 11513 18186 11579 18189
rect 9508 18184 11579 18186
rect 9508 18128 11518 18184
rect 11574 18128 11579 18184
rect 9508 18126 11579 18128
rect 9508 18124 9514 18126
rect 11513 18123 11579 18126
rect 7649 18050 7715 18053
rect 9213 18050 9279 18053
rect 7649 18048 9279 18050
rect 7649 17992 7654 18048
rect 7710 17992 9218 18048
rect 9274 17992 9279 18048
rect 7649 17990 9279 17992
rect 7649 17987 7715 17990
rect 9213 17987 9279 17990
rect 14365 18050 14431 18053
rect 14958 18050 14964 18052
rect 14365 18048 14964 18050
rect 14365 17992 14370 18048
rect 14426 17992 14964 18048
rect 14365 17990 14964 17992
rect 14365 17987 14431 17990
rect 14958 17988 14964 17990
rect 15028 17988 15034 18052
rect 20529 18050 20595 18053
rect 21541 18052 21607 18053
rect 20662 18050 20668 18052
rect 20529 18048 20668 18050
rect 20529 17992 20534 18048
rect 20590 17992 20668 18048
rect 20529 17990 20668 17992
rect 20529 17987 20595 17990
rect 20662 17988 20668 17990
rect 20732 17988 20738 18052
rect 21541 18050 21588 18052
rect 21496 18048 21588 18050
rect 21496 17992 21546 18048
rect 21496 17990 21588 17992
rect 21541 17988 21588 17990
rect 21652 17988 21658 18052
rect 21541 17987 21607 17988
rect 4354 17984 4750 17985
rect 4354 17920 4360 17984
rect 4424 17920 4440 17984
rect 4504 17920 4520 17984
rect 4584 17920 4600 17984
rect 4664 17920 4680 17984
rect 4744 17920 4750 17984
rect 4354 17919 4750 17920
rect 10354 17984 10750 17985
rect 10354 17920 10360 17984
rect 10424 17920 10440 17984
rect 10504 17920 10520 17984
rect 10584 17920 10600 17984
rect 10664 17920 10680 17984
rect 10744 17920 10750 17984
rect 10354 17919 10750 17920
rect 16354 17984 16750 17985
rect 16354 17920 16360 17984
rect 16424 17920 16440 17984
rect 16504 17920 16520 17984
rect 16584 17920 16600 17984
rect 16664 17920 16680 17984
rect 16744 17920 16750 17984
rect 16354 17919 16750 17920
rect 22354 17984 22750 17985
rect 22354 17920 22360 17984
rect 22424 17920 22440 17984
rect 22504 17920 22520 17984
rect 22584 17920 22600 17984
rect 22664 17920 22680 17984
rect 22744 17920 22750 17984
rect 22354 17919 22750 17920
rect 6637 17914 6703 17917
rect 7373 17914 7439 17917
rect 7966 17914 7972 17916
rect 6637 17912 7972 17914
rect 6637 17856 6642 17912
rect 6698 17856 7378 17912
rect 7434 17856 7972 17912
rect 6637 17854 7972 17856
rect 6637 17851 6703 17854
rect 7373 17851 7439 17854
rect 7966 17852 7972 17854
rect 8036 17852 8042 17916
rect 9305 17778 9371 17781
rect 6364 17776 9371 17778
rect 6364 17720 9310 17776
rect 9366 17720 9371 17776
rect 6364 17718 9371 17720
rect 6364 17645 6424 17718
rect 9305 17715 9371 17718
rect 12709 17778 12775 17781
rect 15837 17778 15903 17781
rect 12709 17776 15903 17778
rect 12709 17720 12714 17776
rect 12770 17720 15842 17776
rect 15898 17720 15903 17776
rect 12709 17718 15903 17720
rect 12709 17715 12775 17718
rect 15837 17715 15903 17718
rect 2681 17642 2747 17645
rect 5809 17642 5875 17645
rect 6361 17642 6427 17645
rect 2681 17640 6427 17642
rect 2681 17584 2686 17640
rect 2742 17584 5814 17640
rect 5870 17584 6366 17640
rect 6422 17584 6427 17640
rect 2681 17582 6427 17584
rect 2681 17579 2747 17582
rect 5809 17579 5875 17582
rect 6361 17579 6427 17582
rect 6913 17642 6979 17645
rect 11830 17642 11836 17644
rect 6913 17640 11836 17642
rect 6913 17584 6918 17640
rect 6974 17584 11836 17640
rect 6913 17582 11836 17584
rect 6913 17579 6979 17582
rect 11830 17580 11836 17582
rect 11900 17580 11906 17644
rect 20713 17642 20779 17645
rect 21030 17642 21036 17644
rect 20713 17640 21036 17642
rect 20713 17584 20718 17640
rect 20774 17584 21036 17640
rect 20713 17582 21036 17584
rect 20713 17579 20779 17582
rect 21030 17580 21036 17582
rect 21100 17580 21106 17644
rect 1354 17440 1750 17441
rect 1354 17376 1360 17440
rect 1424 17376 1440 17440
rect 1504 17376 1520 17440
rect 1584 17376 1600 17440
rect 1664 17376 1680 17440
rect 1744 17376 1750 17440
rect 1354 17375 1750 17376
rect 7354 17440 7750 17441
rect 7354 17376 7360 17440
rect 7424 17376 7440 17440
rect 7504 17376 7520 17440
rect 7584 17376 7600 17440
rect 7664 17376 7680 17440
rect 7744 17376 7750 17440
rect 7354 17375 7750 17376
rect 13354 17440 13750 17441
rect 13354 17376 13360 17440
rect 13424 17376 13440 17440
rect 13504 17376 13520 17440
rect 13584 17376 13600 17440
rect 13664 17376 13680 17440
rect 13744 17376 13750 17440
rect 13354 17375 13750 17376
rect 19354 17440 19750 17441
rect 19354 17376 19360 17440
rect 19424 17376 19440 17440
rect 19504 17376 19520 17440
rect 19584 17376 19600 17440
rect 19664 17376 19680 17440
rect 19744 17376 19750 17440
rect 19354 17375 19750 17376
rect 3785 17234 3851 17237
rect 5073 17234 5139 17237
rect 3785 17232 5139 17234
rect 3785 17176 3790 17232
rect 3846 17176 5078 17232
rect 5134 17176 5139 17232
rect 3785 17174 5139 17176
rect 3785 17171 3851 17174
rect 5073 17171 5139 17174
rect 9438 17172 9444 17236
rect 9508 17234 9514 17236
rect 11237 17234 11303 17237
rect 9508 17232 11303 17234
rect 9508 17176 11242 17232
rect 11298 17176 11303 17232
rect 9508 17174 11303 17176
rect 9508 17172 9514 17174
rect 11237 17171 11303 17174
rect 3049 17098 3115 17101
rect 5257 17098 5323 17101
rect 5809 17100 5875 17101
rect 3049 17096 5323 17098
rect 3049 17040 3054 17096
rect 3110 17040 5262 17096
rect 5318 17040 5323 17096
rect 3049 17038 5323 17040
rect 3049 17035 3115 17038
rect 5257 17035 5323 17038
rect 5758 17036 5764 17100
rect 5828 17098 5875 17100
rect 7005 17098 7071 17101
rect 20805 17098 20871 17101
rect 5828 17096 7071 17098
rect 5870 17040 7010 17096
rect 7066 17040 7071 17096
rect 5828 17038 7071 17040
rect 5828 17036 5875 17038
rect 5809 17035 5875 17036
rect 7005 17035 7071 17038
rect 9630 17096 20871 17098
rect 9630 17040 20810 17096
rect 20866 17040 20871 17096
rect 9630 17038 20871 17040
rect 6269 16962 6335 16965
rect 9630 16962 9690 17038
rect 20805 17035 20871 17038
rect 6269 16960 9690 16962
rect 6269 16904 6274 16960
rect 6330 16904 9690 16960
rect 6269 16902 9690 16904
rect 14733 16962 14799 16965
rect 15745 16962 15811 16965
rect 14733 16960 15811 16962
rect 14733 16904 14738 16960
rect 14794 16904 15750 16960
rect 15806 16904 15811 16960
rect 14733 16902 15811 16904
rect 6269 16899 6335 16902
rect 14733 16899 14799 16902
rect 15745 16899 15811 16902
rect 4354 16896 4750 16897
rect 4354 16832 4360 16896
rect 4424 16832 4440 16896
rect 4504 16832 4520 16896
rect 4584 16832 4600 16896
rect 4664 16832 4680 16896
rect 4744 16832 4750 16896
rect 4354 16831 4750 16832
rect 10354 16896 10750 16897
rect 10354 16832 10360 16896
rect 10424 16832 10440 16896
rect 10504 16832 10520 16896
rect 10584 16832 10600 16896
rect 10664 16832 10680 16896
rect 10744 16832 10750 16896
rect 10354 16831 10750 16832
rect 16354 16896 16750 16897
rect 16354 16832 16360 16896
rect 16424 16832 16440 16896
rect 16504 16832 16520 16896
rect 16584 16832 16600 16896
rect 16664 16832 16680 16896
rect 16744 16832 16750 16896
rect 16354 16831 16750 16832
rect 22354 16896 22750 16897
rect 22354 16832 22360 16896
rect 22424 16832 22440 16896
rect 22504 16832 22520 16896
rect 22584 16832 22600 16896
rect 22664 16832 22680 16896
rect 22744 16832 22750 16896
rect 22354 16831 22750 16832
rect 2405 16690 2471 16693
rect 3785 16690 3851 16693
rect 2405 16688 3851 16690
rect 2405 16632 2410 16688
rect 2466 16632 3790 16688
rect 3846 16632 3851 16688
rect 2405 16630 3851 16632
rect 2405 16627 2471 16630
rect 3785 16627 3851 16630
rect 6361 16690 6427 16693
rect 8661 16690 8727 16693
rect 8937 16690 9003 16693
rect 6361 16688 9003 16690
rect 6361 16632 6366 16688
rect 6422 16632 8666 16688
rect 8722 16632 8942 16688
rect 8998 16632 9003 16688
rect 6361 16630 9003 16632
rect 6361 16627 6427 16630
rect 8661 16627 8727 16630
rect 8937 16627 9003 16630
rect 10593 16690 10659 16693
rect 11329 16690 11395 16693
rect 10593 16688 11395 16690
rect 10593 16632 10598 16688
rect 10654 16632 11334 16688
rect 11390 16632 11395 16688
rect 10593 16630 11395 16632
rect 10593 16627 10659 16630
rect 11329 16627 11395 16630
rect 11697 16690 11763 16693
rect 12801 16690 12867 16693
rect 13077 16690 13143 16693
rect 20713 16690 20779 16693
rect 11697 16688 20779 16690
rect 11697 16632 11702 16688
rect 11758 16632 12806 16688
rect 12862 16632 13082 16688
rect 13138 16632 20718 16688
rect 20774 16632 20779 16688
rect 11697 16630 20779 16632
rect 11697 16627 11763 16630
rect 12801 16627 12867 16630
rect 13077 16627 13143 16630
rect 19888 16557 19948 16630
rect 20713 16627 20779 16630
rect 2497 16554 2563 16557
rect 2957 16554 3023 16557
rect 3509 16554 3575 16557
rect 2497 16552 3575 16554
rect 2497 16496 2502 16552
rect 2558 16496 2962 16552
rect 3018 16496 3514 16552
rect 3570 16496 3575 16552
rect 2497 16494 3575 16496
rect 2497 16491 2563 16494
rect 2957 16491 3023 16494
rect 3509 16491 3575 16494
rect 4797 16554 4863 16557
rect 7281 16554 7347 16557
rect 7465 16554 7531 16557
rect 4797 16552 7531 16554
rect 4797 16496 4802 16552
rect 4858 16496 7286 16552
rect 7342 16496 7470 16552
rect 7526 16496 7531 16552
rect 4797 16494 7531 16496
rect 4797 16491 4863 16494
rect 7281 16491 7347 16494
rect 7465 16491 7531 16494
rect 19885 16552 19951 16557
rect 19885 16496 19890 16552
rect 19946 16496 19951 16552
rect 19885 16491 19951 16496
rect 1354 16352 1750 16353
rect 1354 16288 1360 16352
rect 1424 16288 1440 16352
rect 1504 16288 1520 16352
rect 1584 16288 1600 16352
rect 1664 16288 1680 16352
rect 1744 16288 1750 16352
rect 1354 16287 1750 16288
rect 7354 16352 7750 16353
rect 7354 16288 7360 16352
rect 7424 16288 7440 16352
rect 7504 16288 7520 16352
rect 7584 16288 7600 16352
rect 7664 16288 7680 16352
rect 7744 16288 7750 16352
rect 7354 16287 7750 16288
rect 13354 16352 13750 16353
rect 13354 16288 13360 16352
rect 13424 16288 13440 16352
rect 13504 16288 13520 16352
rect 13584 16288 13600 16352
rect 13664 16288 13680 16352
rect 13744 16288 13750 16352
rect 13354 16287 13750 16288
rect 19354 16352 19750 16353
rect 19354 16288 19360 16352
rect 19424 16288 19440 16352
rect 19504 16288 19520 16352
rect 19584 16288 19600 16352
rect 19664 16288 19680 16352
rect 19744 16288 19750 16352
rect 19354 16287 19750 16288
rect 2589 16146 2655 16149
rect 6729 16146 6795 16149
rect 2589 16144 6795 16146
rect 2589 16088 2594 16144
rect 2650 16088 6734 16144
rect 6790 16088 6795 16144
rect 2589 16086 6795 16088
rect 2589 16083 2655 16086
rect 6729 16083 6795 16086
rect 1209 16010 1275 16013
rect 17585 16010 17651 16013
rect 1209 16008 17651 16010
rect 1209 15952 1214 16008
rect 1270 15952 17590 16008
rect 17646 15952 17651 16008
rect 1209 15950 17651 15952
rect 1209 15947 1275 15950
rect 17585 15947 17651 15950
rect 5349 15874 5415 15877
rect 8293 15874 8359 15877
rect 9489 15874 9555 15877
rect 5349 15872 9555 15874
rect 5349 15816 5354 15872
rect 5410 15816 8298 15872
rect 8354 15816 9494 15872
rect 9550 15816 9555 15872
rect 5349 15814 9555 15816
rect 5349 15811 5415 15814
rect 8293 15811 8359 15814
rect 9489 15811 9555 15814
rect 12433 15874 12499 15877
rect 15653 15874 15719 15877
rect 12433 15872 15719 15874
rect 12433 15816 12438 15872
rect 12494 15816 15658 15872
rect 15714 15816 15719 15872
rect 12433 15814 15719 15816
rect 12433 15811 12499 15814
rect 15653 15811 15719 15814
rect 4354 15808 4750 15809
rect 4354 15744 4360 15808
rect 4424 15744 4440 15808
rect 4504 15744 4520 15808
rect 4584 15744 4600 15808
rect 4664 15744 4680 15808
rect 4744 15744 4750 15808
rect 4354 15743 4750 15744
rect 10354 15808 10750 15809
rect 10354 15744 10360 15808
rect 10424 15744 10440 15808
rect 10504 15744 10520 15808
rect 10584 15744 10600 15808
rect 10664 15744 10680 15808
rect 10744 15744 10750 15808
rect 10354 15743 10750 15744
rect 16354 15808 16750 15809
rect 16354 15744 16360 15808
rect 16424 15744 16440 15808
rect 16504 15744 16520 15808
rect 16584 15744 16600 15808
rect 16664 15744 16680 15808
rect 16744 15744 16750 15808
rect 16354 15743 16750 15744
rect 22354 15808 22750 15809
rect 22354 15744 22360 15808
rect 22424 15744 22440 15808
rect 22504 15744 22520 15808
rect 22584 15744 22600 15808
rect 22664 15744 22680 15808
rect 22744 15744 22750 15808
rect 22354 15743 22750 15744
rect 5993 15738 6059 15741
rect 8753 15738 8819 15741
rect 16021 15738 16087 15741
rect 5993 15736 8819 15738
rect 5993 15680 5998 15736
rect 6054 15680 8758 15736
rect 8814 15680 8819 15736
rect 5993 15678 8819 15680
rect 5993 15675 6059 15678
rect 8753 15675 8819 15678
rect 12390 15736 16087 15738
rect 12390 15680 16026 15736
rect 16082 15680 16087 15736
rect 12390 15678 16087 15680
rect 5441 15602 5507 15605
rect 6637 15602 6703 15605
rect 5441 15600 6703 15602
rect 5441 15544 5446 15600
rect 5502 15544 6642 15600
rect 6698 15544 6703 15600
rect 5441 15542 6703 15544
rect 5441 15539 5507 15542
rect 6637 15539 6703 15542
rect 7373 15602 7439 15605
rect 12065 15602 12131 15605
rect 12390 15602 12450 15678
rect 16021 15675 16087 15678
rect 7373 15600 9000 15602
rect 7373 15544 7378 15600
rect 7434 15544 9000 15600
rect 7373 15542 9000 15544
rect 7373 15539 7439 15542
rect 2865 15466 2931 15469
rect 3325 15466 3391 15469
rect 3734 15466 3740 15468
rect 2865 15464 3740 15466
rect 2865 15408 2870 15464
rect 2926 15408 3330 15464
rect 3386 15408 3740 15464
rect 2865 15406 3740 15408
rect 2865 15403 2931 15406
rect 3325 15403 3391 15406
rect 3734 15404 3740 15406
rect 3804 15404 3810 15468
rect 4981 15466 5047 15469
rect 8293 15466 8359 15469
rect 4294 15464 8359 15466
rect 4294 15408 4986 15464
rect 5042 15408 8298 15464
rect 8354 15408 8359 15464
rect 4294 15406 8359 15408
rect 1354 15264 1750 15265
rect 1354 15200 1360 15264
rect 1424 15200 1440 15264
rect 1504 15200 1520 15264
rect 1584 15200 1600 15264
rect 1664 15200 1680 15264
rect 1744 15200 1750 15264
rect 1354 15199 1750 15200
rect 4294 15197 4354 15406
rect 4981 15403 5047 15406
rect 8293 15403 8359 15406
rect 8940 15466 9000 15542
rect 12065 15600 12450 15602
rect 12065 15544 12070 15600
rect 12126 15544 12450 15600
rect 12065 15542 12450 15544
rect 12065 15539 12131 15542
rect 18086 15540 18092 15604
rect 18156 15602 18162 15604
rect 18689 15602 18755 15605
rect 18156 15600 18755 15602
rect 18156 15544 18694 15600
rect 18750 15544 18755 15600
rect 18156 15542 18755 15544
rect 18156 15540 18162 15542
rect 18689 15539 18755 15542
rect 19333 15466 19399 15469
rect 8940 15464 19399 15466
rect 8940 15408 19338 15464
rect 19394 15408 19399 15464
rect 8940 15406 19399 15408
rect 8940 15333 9000 15406
rect 19333 15403 19399 15406
rect 8937 15328 9003 15333
rect 8937 15272 8942 15328
rect 8998 15272 9003 15328
rect 8937 15267 9003 15272
rect 11278 15268 11284 15332
rect 11348 15330 11354 15332
rect 11605 15330 11671 15333
rect 11348 15328 11671 15330
rect 11348 15272 11610 15328
rect 11666 15272 11671 15328
rect 11348 15270 11671 15272
rect 11348 15268 11354 15270
rect 11605 15267 11671 15270
rect 7354 15264 7750 15265
rect 7354 15200 7360 15264
rect 7424 15200 7440 15264
rect 7504 15200 7520 15264
rect 7584 15200 7600 15264
rect 7664 15200 7680 15264
rect 7744 15200 7750 15264
rect 7354 15199 7750 15200
rect 13354 15264 13750 15265
rect 13354 15200 13360 15264
rect 13424 15200 13440 15264
rect 13504 15200 13520 15264
rect 13584 15200 13600 15264
rect 13664 15200 13680 15264
rect 13744 15200 13750 15264
rect 13354 15199 13750 15200
rect 19354 15264 19750 15265
rect 19354 15200 19360 15264
rect 19424 15200 19440 15264
rect 19504 15200 19520 15264
rect 19584 15200 19600 15264
rect 19664 15200 19680 15264
rect 19744 15200 19750 15264
rect 19354 15199 19750 15200
rect 4245 15192 4354 15197
rect 4245 15136 4250 15192
rect 4306 15136 4354 15192
rect 4245 15134 4354 15136
rect 10961 15194 11027 15197
rect 11605 15194 11671 15197
rect 12893 15194 12959 15197
rect 10961 15192 12959 15194
rect 10961 15136 10966 15192
rect 11022 15136 11610 15192
rect 11666 15136 12898 15192
rect 12954 15136 12959 15192
rect 10961 15134 12959 15136
rect 4245 15131 4311 15134
rect 10961 15131 11027 15134
rect 11605 15131 11671 15134
rect 12893 15131 12959 15134
rect 4429 15058 4495 15061
rect 6453 15058 6519 15061
rect 4429 15056 6519 15058
rect 4429 15000 4434 15056
rect 4490 15000 6458 15056
rect 6514 15000 6519 15056
rect 4429 14998 6519 15000
rect 4429 14995 4495 14998
rect 6453 14995 6519 14998
rect 10041 15058 10107 15061
rect 10593 15058 10659 15061
rect 10910 15058 10916 15060
rect 10041 15056 10916 15058
rect 10041 15000 10046 15056
rect 10102 15000 10598 15056
rect 10654 15000 10916 15056
rect 10041 14998 10916 15000
rect 10041 14995 10107 14998
rect 10593 14995 10659 14998
rect 10910 14996 10916 14998
rect 10980 14996 10986 15060
rect 12157 15058 12223 15061
rect 18505 15058 18571 15061
rect 12157 15056 18571 15058
rect 12157 15000 12162 15056
rect 12218 15000 18510 15056
rect 18566 15000 18571 15056
rect 12157 14998 18571 15000
rect 12157 14995 12223 14998
rect 18505 14995 18571 14998
rect 4705 14922 4771 14925
rect 5257 14922 5323 14925
rect 4705 14920 5323 14922
rect 4705 14864 4710 14920
rect 4766 14864 5262 14920
rect 5318 14864 5323 14920
rect 4705 14862 5323 14864
rect 4705 14859 4771 14862
rect 5257 14859 5323 14862
rect 8845 14922 8911 14925
rect 12065 14922 12131 14925
rect 8845 14920 12131 14922
rect 8845 14864 8850 14920
rect 8906 14864 12070 14920
rect 12126 14864 12131 14920
rect 8845 14862 12131 14864
rect 8845 14859 8911 14862
rect 12065 14859 12131 14862
rect 8201 14786 8267 14789
rect 8477 14786 8543 14789
rect 9213 14786 9279 14789
rect 8201 14784 9279 14786
rect 8201 14728 8206 14784
rect 8262 14728 8482 14784
rect 8538 14728 9218 14784
rect 9274 14728 9279 14784
rect 8201 14726 9279 14728
rect 8201 14723 8267 14726
rect 8477 14723 8543 14726
rect 9213 14723 9279 14726
rect 4354 14720 4750 14721
rect 4354 14656 4360 14720
rect 4424 14656 4440 14720
rect 4504 14656 4520 14720
rect 4584 14656 4600 14720
rect 4664 14656 4680 14720
rect 4744 14656 4750 14720
rect 4354 14655 4750 14656
rect 10354 14720 10750 14721
rect 10354 14656 10360 14720
rect 10424 14656 10440 14720
rect 10504 14656 10520 14720
rect 10584 14656 10600 14720
rect 10664 14656 10680 14720
rect 10744 14656 10750 14720
rect 10354 14655 10750 14656
rect 16354 14720 16750 14721
rect 16354 14656 16360 14720
rect 16424 14656 16440 14720
rect 16504 14656 16520 14720
rect 16584 14656 16600 14720
rect 16664 14656 16680 14720
rect 16744 14656 16750 14720
rect 16354 14655 16750 14656
rect 22354 14720 22750 14721
rect 22354 14656 22360 14720
rect 22424 14656 22440 14720
rect 22504 14656 22520 14720
rect 22584 14656 22600 14720
rect 22664 14656 22680 14720
rect 22744 14656 22750 14720
rect 22354 14655 22750 14656
rect 5993 14650 6059 14653
rect 9581 14650 9647 14653
rect 5993 14648 9647 14650
rect 5993 14592 5998 14648
rect 6054 14592 9586 14648
rect 9642 14592 9647 14648
rect 5993 14590 9647 14592
rect 5993 14587 6059 14590
rect 9581 14587 9647 14590
rect 10133 14648 10199 14653
rect 10133 14592 10138 14648
rect 10194 14592 10199 14648
rect 10133 14587 10199 14592
rect 11830 14588 11836 14652
rect 11900 14650 11906 14652
rect 12065 14650 12131 14653
rect 11900 14648 12131 14650
rect 11900 14592 12070 14648
rect 12126 14592 12131 14648
rect 11900 14590 12131 14592
rect 11900 14588 11906 14590
rect 12065 14587 12131 14590
rect 12709 14650 12775 14653
rect 12709 14648 16130 14650
rect 12709 14592 12714 14648
rect 12770 14592 16130 14648
rect 12709 14590 16130 14592
rect 12709 14587 12775 14590
rect 3877 14514 3943 14517
rect 5257 14514 5323 14517
rect 3877 14512 5323 14514
rect 3877 14456 3882 14512
rect 3938 14456 5262 14512
rect 5318 14456 5323 14512
rect 3877 14454 5323 14456
rect 3877 14451 3943 14454
rect 5257 14451 5323 14454
rect 8293 14514 8359 14517
rect 9029 14514 9095 14517
rect 8293 14512 9095 14514
rect 8293 14456 8298 14512
rect 8354 14456 9034 14512
rect 9090 14456 9095 14512
rect 8293 14454 9095 14456
rect 8293 14451 8359 14454
rect 9029 14451 9095 14454
rect 9765 14514 9831 14517
rect 10136 14514 10196 14587
rect 14089 14514 14155 14517
rect 9765 14512 14155 14514
rect 9765 14456 9770 14512
rect 9826 14456 14094 14512
rect 14150 14456 14155 14512
rect 9765 14454 14155 14456
rect 16070 14514 16130 14590
rect 19190 14514 19196 14516
rect 16070 14454 19196 14514
rect 9765 14451 9831 14454
rect 14089 14451 14155 14454
rect 19190 14452 19196 14454
rect 19260 14514 19266 14516
rect 19333 14514 19399 14517
rect 19260 14512 19399 14514
rect 19260 14456 19338 14512
rect 19394 14456 19399 14512
rect 19260 14454 19399 14456
rect 19260 14452 19266 14454
rect 19333 14451 19399 14454
rect 4613 14378 4679 14381
rect 5533 14378 5599 14381
rect 4613 14376 5599 14378
rect 4613 14320 4618 14376
rect 4674 14320 5538 14376
rect 5594 14320 5599 14376
rect 4613 14318 5599 14320
rect 4613 14315 4679 14318
rect 5533 14315 5599 14318
rect 10133 14378 10199 14381
rect 12157 14378 12223 14381
rect 10133 14376 12223 14378
rect 10133 14320 10138 14376
rect 10194 14320 12162 14376
rect 12218 14320 12223 14376
rect 10133 14318 12223 14320
rect 10133 14315 10199 14318
rect 12157 14315 12223 14318
rect 12617 14378 12683 14381
rect 15193 14378 15259 14381
rect 12617 14376 15259 14378
rect 12617 14320 12622 14376
rect 12678 14320 15198 14376
rect 15254 14320 15259 14376
rect 12617 14318 15259 14320
rect 12617 14315 12683 14318
rect 15193 14315 15259 14318
rect 10685 14242 10751 14245
rect 12934 14242 12940 14244
rect 10685 14240 12940 14242
rect 10685 14184 10690 14240
rect 10746 14184 12940 14240
rect 10685 14182 12940 14184
rect 10685 14179 10751 14182
rect 12934 14180 12940 14182
rect 13004 14180 13010 14244
rect 14549 14242 14615 14245
rect 18689 14242 18755 14245
rect 14549 14240 18755 14242
rect 14549 14184 14554 14240
rect 14610 14184 18694 14240
rect 18750 14184 18755 14240
rect 14549 14182 18755 14184
rect 14549 14179 14615 14182
rect 18689 14179 18755 14182
rect 1354 14176 1750 14177
rect 1354 14112 1360 14176
rect 1424 14112 1440 14176
rect 1504 14112 1520 14176
rect 1584 14112 1600 14176
rect 1664 14112 1680 14176
rect 1744 14112 1750 14176
rect 1354 14111 1750 14112
rect 7354 14176 7750 14177
rect 7354 14112 7360 14176
rect 7424 14112 7440 14176
rect 7504 14112 7520 14176
rect 7584 14112 7600 14176
rect 7664 14112 7680 14176
rect 7744 14112 7750 14176
rect 7354 14111 7750 14112
rect 13354 14176 13750 14177
rect 13354 14112 13360 14176
rect 13424 14112 13440 14176
rect 13504 14112 13520 14176
rect 13584 14112 13600 14176
rect 13664 14112 13680 14176
rect 13744 14112 13750 14176
rect 13354 14111 13750 14112
rect 19354 14176 19750 14177
rect 19354 14112 19360 14176
rect 19424 14112 19440 14176
rect 19504 14112 19520 14176
rect 19584 14112 19600 14176
rect 19664 14112 19680 14176
rect 19744 14112 19750 14176
rect 19354 14111 19750 14112
rect 10133 14106 10199 14109
rect 11053 14106 11119 14109
rect 10133 14104 11119 14106
rect 10133 14048 10138 14104
rect 10194 14048 11058 14104
rect 11114 14048 11119 14104
rect 10133 14046 11119 14048
rect 10133 14043 10199 14046
rect 11053 14043 11119 14046
rect 6085 13970 6151 13973
rect 7373 13970 7439 13973
rect 6085 13968 7439 13970
rect 6085 13912 6090 13968
rect 6146 13912 7378 13968
rect 7434 13912 7439 13968
rect 6085 13910 7439 13912
rect 6085 13907 6151 13910
rect 7373 13907 7439 13910
rect 8109 13970 8175 13973
rect 15837 13970 15903 13973
rect 8109 13968 15903 13970
rect 8109 13912 8114 13968
rect 8170 13912 15842 13968
rect 15898 13912 15903 13968
rect 8109 13910 15903 13912
rect 8109 13907 8175 13910
rect 15837 13907 15903 13910
rect 5533 13834 5599 13837
rect 5942 13834 5948 13836
rect 5533 13832 5948 13834
rect 5533 13776 5538 13832
rect 5594 13776 5948 13832
rect 5533 13774 5948 13776
rect 5533 13771 5599 13774
rect 5942 13772 5948 13774
rect 6012 13772 6018 13836
rect 10317 13834 10383 13837
rect 12249 13834 12315 13837
rect 13261 13834 13327 13837
rect 10182 13832 10978 13834
rect 10182 13776 10322 13832
rect 10378 13776 10978 13832
rect 10182 13774 10978 13776
rect 8017 13698 8083 13701
rect 9070 13698 9076 13700
rect 8017 13696 9076 13698
rect 8017 13640 8022 13696
rect 8078 13640 9076 13696
rect 8017 13638 9076 13640
rect 8017 13635 8083 13638
rect 9070 13636 9076 13638
rect 9140 13636 9146 13700
rect 9489 13698 9555 13701
rect 10182 13698 10242 13774
rect 10317 13771 10383 13774
rect 9489 13696 10242 13698
rect 9489 13640 9494 13696
rect 9550 13640 10242 13696
rect 9489 13638 10242 13640
rect 10918 13698 10978 13774
rect 12249 13832 13327 13834
rect 12249 13776 12254 13832
rect 12310 13776 13266 13832
rect 13322 13776 13327 13832
rect 12249 13774 13327 13776
rect 12249 13771 12315 13774
rect 13261 13771 13327 13774
rect 15745 13698 15811 13701
rect 10918 13696 15811 13698
rect 10918 13640 15750 13696
rect 15806 13640 15811 13696
rect 10918 13638 15811 13640
rect 9489 13635 9555 13638
rect 15745 13635 15811 13638
rect 4354 13632 4750 13633
rect 4354 13568 4360 13632
rect 4424 13568 4440 13632
rect 4504 13568 4520 13632
rect 4584 13568 4600 13632
rect 4664 13568 4680 13632
rect 4744 13568 4750 13632
rect 4354 13567 4750 13568
rect 10354 13632 10750 13633
rect 10354 13568 10360 13632
rect 10424 13568 10440 13632
rect 10504 13568 10520 13632
rect 10584 13568 10600 13632
rect 10664 13568 10680 13632
rect 10744 13568 10750 13632
rect 10354 13567 10750 13568
rect 16354 13632 16750 13633
rect 16354 13568 16360 13632
rect 16424 13568 16440 13632
rect 16504 13568 16520 13632
rect 16584 13568 16600 13632
rect 16664 13568 16680 13632
rect 16744 13568 16750 13632
rect 16354 13567 16750 13568
rect 22354 13632 22750 13633
rect 22354 13568 22360 13632
rect 22424 13568 22440 13632
rect 22504 13568 22520 13632
rect 22584 13568 22600 13632
rect 22664 13568 22680 13632
rect 22744 13568 22750 13632
rect 22354 13567 22750 13568
rect 7966 13500 7972 13564
rect 8036 13562 8042 13564
rect 8937 13562 9003 13565
rect 12709 13562 12775 13565
rect 8036 13560 9003 13562
rect 8036 13504 8942 13560
rect 8998 13504 9003 13560
rect 8036 13502 9003 13504
rect 8036 13500 8042 13502
rect 8937 13499 9003 13502
rect 12390 13560 12775 13562
rect 12390 13504 12714 13560
rect 12770 13504 12775 13560
rect 12390 13502 12775 13504
rect 4245 13426 4311 13429
rect 12390 13426 12450 13502
rect 12709 13499 12775 13502
rect 12801 13428 12867 13429
rect 4245 13424 12450 13426
rect 4245 13368 4250 13424
rect 4306 13368 12450 13424
rect 4245 13366 12450 13368
rect 4245 13363 4311 13366
rect 12750 13364 12756 13428
rect 12820 13426 12867 13428
rect 12820 13424 12912 13426
rect 12862 13368 12912 13424
rect 12820 13366 12912 13368
rect 12820 13364 12867 13366
rect 12801 13363 12867 13364
rect 6821 13290 6887 13293
rect 7649 13290 7715 13293
rect 6821 13288 7715 13290
rect 6821 13232 6826 13288
rect 6882 13232 7654 13288
rect 7710 13232 7715 13288
rect 6821 13230 7715 13232
rect 6821 13227 6887 13230
rect 7649 13227 7715 13230
rect 11646 13228 11652 13292
rect 11716 13290 11722 13292
rect 18454 13290 18460 13292
rect 11716 13230 18460 13290
rect 11716 13228 11722 13230
rect 18454 13228 18460 13230
rect 18524 13228 18530 13292
rect 12617 13154 12683 13157
rect 13118 13154 13124 13156
rect 12617 13152 13124 13154
rect 12617 13096 12622 13152
rect 12678 13096 13124 13152
rect 12617 13094 13124 13096
rect 12617 13091 12683 13094
rect 13118 13092 13124 13094
rect 13188 13092 13194 13156
rect 1354 13088 1750 13089
rect 1354 13024 1360 13088
rect 1424 13024 1440 13088
rect 1504 13024 1520 13088
rect 1584 13024 1600 13088
rect 1664 13024 1680 13088
rect 1744 13024 1750 13088
rect 1354 13023 1750 13024
rect 7354 13088 7750 13089
rect 7354 13024 7360 13088
rect 7424 13024 7440 13088
rect 7504 13024 7520 13088
rect 7584 13024 7600 13088
rect 7664 13024 7680 13088
rect 7744 13024 7750 13088
rect 7354 13023 7750 13024
rect 13354 13088 13750 13089
rect 13354 13024 13360 13088
rect 13424 13024 13440 13088
rect 13504 13024 13520 13088
rect 13584 13024 13600 13088
rect 13664 13024 13680 13088
rect 13744 13024 13750 13088
rect 13354 13023 13750 13024
rect 19354 13088 19750 13089
rect 19354 13024 19360 13088
rect 19424 13024 19440 13088
rect 19504 13024 19520 13088
rect 19584 13024 19600 13088
rect 19664 13024 19680 13088
rect 19744 13024 19750 13088
rect 19354 13023 19750 13024
rect 9765 13018 9831 13021
rect 9765 13016 13232 13018
rect 9765 12960 9770 13016
rect 9826 12960 13232 13016
rect 9765 12958 13232 12960
rect 9765 12955 9831 12958
rect 2313 12882 2379 12885
rect 9254 12882 9260 12884
rect 2313 12880 9260 12882
rect 2313 12824 2318 12880
rect 2374 12824 9260 12880
rect 2313 12822 9260 12824
rect 2313 12819 2379 12822
rect 9254 12820 9260 12822
rect 9324 12820 9330 12884
rect 9765 12882 9831 12885
rect 12341 12882 12407 12885
rect 12617 12882 12683 12885
rect 9765 12880 12683 12882
rect 9765 12824 9770 12880
rect 9826 12824 12346 12880
rect 12402 12824 12622 12880
rect 12678 12824 12683 12880
rect 9765 12822 12683 12824
rect 13172 12882 13232 12958
rect 13905 12882 13971 12885
rect 13172 12880 13971 12882
rect 13172 12824 13910 12880
rect 13966 12824 13971 12880
rect 13172 12822 13971 12824
rect 9765 12819 9831 12822
rect 12341 12819 12407 12822
rect 12617 12819 12683 12822
rect 13905 12819 13971 12822
rect 19333 12882 19399 12885
rect 19517 12882 19583 12885
rect 20161 12882 20227 12885
rect 20805 12884 20871 12885
rect 20805 12882 20852 12884
rect 19333 12880 20227 12882
rect 19333 12824 19338 12880
rect 19394 12824 19522 12880
rect 19578 12824 20166 12880
rect 20222 12824 20227 12880
rect 19333 12822 20227 12824
rect 20764 12880 20852 12882
rect 20916 12882 20922 12884
rect 21214 12882 21220 12884
rect 20764 12824 20810 12880
rect 20764 12822 20852 12824
rect 19333 12819 19399 12822
rect 19517 12819 19583 12822
rect 20161 12819 20227 12822
rect 20805 12820 20852 12822
rect 20916 12822 21220 12882
rect 20916 12820 20922 12822
rect 21214 12820 21220 12822
rect 21284 12820 21290 12884
rect 20805 12819 20871 12820
rect 8293 12746 8359 12749
rect 8569 12746 8635 12749
rect 8293 12744 10978 12746
rect 8293 12688 8298 12744
rect 8354 12688 8574 12744
rect 8630 12688 10978 12744
rect 8293 12686 10978 12688
rect 8293 12683 8359 12686
rect 8569 12683 8635 12686
rect 10918 12610 10978 12686
rect 12566 12610 12572 12612
rect 10918 12550 12572 12610
rect 12566 12548 12572 12550
rect 12636 12548 12642 12612
rect 4354 12544 4750 12545
rect 4354 12480 4360 12544
rect 4424 12480 4440 12544
rect 4504 12480 4520 12544
rect 4584 12480 4600 12544
rect 4664 12480 4680 12544
rect 4744 12480 4750 12544
rect 4354 12479 4750 12480
rect 10354 12544 10750 12545
rect 10354 12480 10360 12544
rect 10424 12480 10440 12544
rect 10504 12480 10520 12544
rect 10584 12480 10600 12544
rect 10664 12480 10680 12544
rect 10744 12480 10750 12544
rect 10354 12479 10750 12480
rect 16354 12544 16750 12545
rect 16354 12480 16360 12544
rect 16424 12480 16440 12544
rect 16504 12480 16520 12544
rect 16584 12480 16600 12544
rect 16664 12480 16680 12544
rect 16744 12480 16750 12544
rect 16354 12479 16750 12480
rect 22354 12544 22750 12545
rect 22354 12480 22360 12544
rect 22424 12480 22440 12544
rect 22504 12480 22520 12544
rect 22584 12480 22600 12544
rect 22664 12480 22680 12544
rect 22744 12480 22750 12544
rect 22354 12479 22750 12480
rect 12341 12474 12407 12477
rect 15469 12474 15535 12477
rect 12341 12472 15535 12474
rect 12341 12416 12346 12472
rect 12402 12416 15474 12472
rect 15530 12416 15535 12472
rect 12341 12414 15535 12416
rect 12341 12411 12407 12414
rect 15469 12411 15535 12414
rect 11329 12338 11395 12341
rect 11789 12338 11855 12341
rect 18045 12338 18111 12341
rect 11329 12336 18111 12338
rect 11329 12280 11334 12336
rect 11390 12280 11794 12336
rect 11850 12280 18050 12336
rect 18106 12280 18111 12336
rect 11329 12278 18111 12280
rect 11329 12275 11395 12278
rect 11789 12275 11855 12278
rect 18045 12275 18111 12278
rect 1485 12202 1551 12205
rect 1945 12202 2011 12205
rect 1485 12200 2011 12202
rect 1485 12144 1490 12200
rect 1546 12144 1950 12200
rect 2006 12144 2011 12200
rect 1485 12142 2011 12144
rect 1485 12139 1551 12142
rect 1945 12139 2011 12142
rect 5441 12202 5507 12205
rect 8385 12202 8451 12205
rect 9213 12202 9279 12205
rect 5441 12200 9279 12202
rect 5441 12144 5446 12200
rect 5502 12144 8390 12200
rect 8446 12144 9218 12200
rect 9274 12144 9279 12200
rect 5441 12142 9279 12144
rect 5441 12139 5507 12142
rect 8385 12139 8451 12142
rect 9213 12139 9279 12142
rect 12934 12140 12940 12204
rect 13004 12202 13010 12204
rect 16665 12202 16731 12205
rect 13004 12200 16731 12202
rect 13004 12144 16670 12200
rect 16726 12144 16731 12200
rect 13004 12142 16731 12144
rect 13004 12140 13010 12142
rect 16665 12139 16731 12142
rect 19517 12202 19583 12205
rect 20621 12204 20687 12205
rect 19517 12200 19948 12202
rect 19517 12144 19522 12200
rect 19578 12144 19948 12200
rect 19517 12142 19948 12144
rect 19517 12139 19583 12142
rect 10910 12004 10916 12068
rect 10980 12066 10986 12068
rect 11789 12066 11855 12069
rect 10980 12064 11855 12066
rect 10980 12008 11794 12064
rect 11850 12008 11855 12064
rect 10980 12006 11855 12008
rect 10980 12004 10986 12006
rect 11789 12003 11855 12006
rect 15377 12066 15443 12069
rect 17493 12066 17559 12069
rect 15377 12064 17559 12066
rect 15377 12008 15382 12064
rect 15438 12008 17498 12064
rect 17554 12008 17559 12064
rect 15377 12006 17559 12008
rect 15377 12003 15443 12006
rect 17493 12003 17559 12006
rect 1354 12000 1750 12001
rect 1354 11936 1360 12000
rect 1424 11936 1440 12000
rect 1504 11936 1520 12000
rect 1584 11936 1600 12000
rect 1664 11936 1680 12000
rect 1744 11936 1750 12000
rect 1354 11935 1750 11936
rect 7354 12000 7750 12001
rect 7354 11936 7360 12000
rect 7424 11936 7440 12000
rect 7504 11936 7520 12000
rect 7584 11936 7600 12000
rect 7664 11936 7680 12000
rect 7744 11936 7750 12000
rect 7354 11935 7750 11936
rect 13354 12000 13750 12001
rect 13354 11936 13360 12000
rect 13424 11936 13440 12000
rect 13504 11936 13520 12000
rect 13584 11936 13600 12000
rect 13664 11936 13680 12000
rect 13744 11936 13750 12000
rect 13354 11935 13750 11936
rect 19354 12000 19750 12001
rect 19354 11936 19360 12000
rect 19424 11936 19440 12000
rect 19504 11936 19520 12000
rect 19584 11936 19600 12000
rect 19664 11936 19680 12000
rect 19744 11936 19750 12000
rect 19354 11935 19750 11936
rect 10869 11930 10935 11933
rect 12617 11930 12683 11933
rect 10869 11928 12683 11930
rect 10869 11872 10874 11928
rect 10930 11872 12622 11928
rect 12678 11872 12683 11928
rect 10869 11870 12683 11872
rect 10869 11867 10935 11870
rect 12617 11867 12683 11870
rect 14181 11930 14247 11933
rect 18321 11930 18387 11933
rect 14181 11928 18387 11930
rect 14181 11872 14186 11928
rect 14242 11872 18326 11928
rect 18382 11872 18387 11928
rect 14181 11870 18387 11872
rect 14181 11867 14247 11870
rect 18321 11867 18387 11870
rect 4245 11794 4311 11797
rect 11278 11794 11284 11796
rect 4245 11792 11284 11794
rect 4245 11736 4250 11792
rect 4306 11736 11284 11792
rect 4245 11734 11284 11736
rect 4245 11731 4311 11734
rect 11278 11732 11284 11734
rect 11348 11732 11354 11796
rect 13169 11794 13235 11797
rect 19517 11794 19583 11797
rect 19888 11794 19948 12142
rect 20621 12200 20668 12204
rect 20732 12202 20738 12204
rect 20621 12144 20626 12200
rect 20621 12140 20668 12144
rect 20732 12142 20778 12202
rect 20732 12140 20738 12142
rect 20621 12139 20687 12140
rect 13169 11792 18154 11794
rect 13169 11736 13174 11792
rect 13230 11736 18154 11792
rect 13169 11734 18154 11736
rect 13169 11731 13235 11734
rect 18094 11661 18154 11734
rect 19517 11792 19948 11794
rect 19517 11736 19522 11792
rect 19578 11736 19948 11792
rect 19517 11734 19948 11736
rect 19517 11731 19583 11734
rect 10174 11596 10180 11660
rect 10244 11658 10250 11660
rect 11278 11658 11284 11660
rect 10244 11598 11284 11658
rect 10244 11596 10250 11598
rect 11278 11596 11284 11598
rect 11348 11596 11354 11660
rect 12617 11658 12683 11661
rect 13537 11658 13603 11661
rect 12617 11656 13603 11658
rect 12617 11600 12622 11656
rect 12678 11600 13542 11656
rect 13598 11600 13603 11656
rect 12617 11598 13603 11600
rect 12617 11595 12683 11598
rect 13537 11595 13603 11598
rect 14181 11656 14247 11661
rect 14181 11600 14186 11656
rect 14242 11600 14247 11656
rect 14181 11595 14247 11600
rect 14365 11658 14431 11661
rect 16573 11658 16639 11661
rect 14365 11656 16639 11658
rect 14365 11600 14370 11656
rect 14426 11600 16578 11656
rect 16634 11600 16639 11656
rect 14365 11598 16639 11600
rect 18094 11656 18203 11661
rect 18094 11600 18142 11656
rect 18198 11600 18203 11656
rect 18094 11598 18203 11600
rect 14365 11595 14431 11598
rect 16573 11595 16639 11598
rect 18137 11595 18203 11598
rect 12525 11524 12591 11525
rect 12525 11520 12572 11524
rect 12636 11522 12642 11524
rect 12525 11464 12530 11520
rect 12525 11460 12572 11464
rect 12636 11462 12682 11522
rect 12636 11460 12642 11462
rect 12525 11459 12591 11460
rect 4354 11456 4750 11457
rect 4354 11392 4360 11456
rect 4424 11392 4440 11456
rect 4504 11392 4520 11456
rect 4584 11392 4600 11456
rect 4664 11392 4680 11456
rect 4744 11392 4750 11456
rect 4354 11391 4750 11392
rect 10354 11456 10750 11457
rect 10354 11392 10360 11456
rect 10424 11392 10440 11456
rect 10504 11392 10520 11456
rect 10584 11392 10600 11456
rect 10664 11392 10680 11456
rect 10744 11392 10750 11456
rect 10354 11391 10750 11392
rect 11789 11386 11855 11389
rect 14184 11386 14244 11595
rect 18689 11522 18755 11525
rect 19057 11522 19123 11525
rect 18689 11520 19123 11522
rect 18689 11464 18694 11520
rect 18750 11464 19062 11520
rect 19118 11464 19123 11520
rect 18689 11462 19123 11464
rect 18689 11459 18755 11462
rect 19057 11459 19123 11462
rect 16354 11456 16750 11457
rect 16354 11392 16360 11456
rect 16424 11392 16440 11456
rect 16504 11392 16520 11456
rect 16584 11392 16600 11456
rect 16664 11392 16680 11456
rect 16744 11392 16750 11456
rect 16354 11391 16750 11392
rect 22354 11456 22750 11457
rect 22354 11392 22360 11456
rect 22424 11392 22440 11456
rect 22504 11392 22520 11456
rect 22584 11392 22600 11456
rect 22664 11392 22680 11456
rect 22744 11392 22750 11456
rect 22354 11391 22750 11392
rect 11789 11384 14244 11386
rect 11789 11328 11794 11384
rect 11850 11328 14244 11384
rect 11789 11326 14244 11328
rect 11789 11323 11855 11326
rect 8293 11250 8359 11253
rect 12709 11250 12775 11253
rect 13169 11250 13235 11253
rect 14273 11250 14339 11253
rect 8293 11248 12450 11250
rect 8293 11192 8298 11248
rect 8354 11192 12450 11248
rect 8293 11190 12450 11192
rect 8293 11187 8359 11190
rect 5022 11052 5028 11116
rect 5092 11114 5098 11116
rect 5257 11114 5323 11117
rect 5092 11112 5323 11114
rect 5092 11056 5262 11112
rect 5318 11056 5323 11112
rect 5092 11054 5323 11056
rect 5092 11052 5098 11054
rect 5257 11051 5323 11054
rect 7833 11114 7899 11117
rect 11513 11114 11579 11117
rect 12014 11114 12020 11116
rect 7833 11112 8034 11114
rect 7833 11056 7838 11112
rect 7894 11056 8034 11112
rect 7833 11054 8034 11056
rect 7833 11051 7899 11054
rect 7974 10980 8034 11054
rect 11513 11112 12020 11114
rect 11513 11056 11518 11112
rect 11574 11056 12020 11112
rect 11513 11054 12020 11056
rect 11513 11051 11579 11054
rect 12014 11052 12020 11054
rect 12084 11052 12090 11116
rect 12390 11114 12450 11190
rect 12709 11248 14339 11250
rect 12709 11192 12714 11248
rect 12770 11192 13174 11248
rect 13230 11192 14278 11248
rect 14334 11192 14339 11248
rect 12709 11190 14339 11192
rect 12709 11187 12775 11190
rect 13169 11187 13235 11190
rect 14273 11187 14339 11190
rect 15377 11250 15443 11253
rect 16297 11250 16363 11253
rect 15377 11248 16363 11250
rect 15377 11192 15382 11248
rect 15438 11192 16302 11248
rect 16358 11192 16363 11248
rect 15377 11190 16363 11192
rect 15377 11187 15443 11190
rect 16297 11187 16363 11190
rect 18873 11250 18939 11253
rect 20253 11250 20319 11253
rect 18873 11248 20319 11250
rect 18873 11192 18878 11248
rect 18934 11192 20258 11248
rect 20314 11192 20319 11248
rect 18873 11190 20319 11192
rect 18873 11187 18939 11190
rect 20253 11187 20319 11190
rect 12801 11114 12867 11117
rect 12390 11112 12867 11114
rect 12390 11056 12806 11112
rect 12862 11056 12867 11112
rect 12390 11054 12867 11056
rect 12801 11051 12867 11054
rect 13077 11114 13143 11117
rect 14181 11114 14247 11117
rect 13077 11112 14247 11114
rect 13077 11056 13082 11112
rect 13138 11056 14186 11112
rect 14242 11056 14247 11112
rect 13077 11054 14247 11056
rect 13077 11051 13143 11054
rect 14181 11051 14247 11054
rect 18321 11114 18387 11117
rect 19333 11114 19399 11117
rect 18321 11112 19399 11114
rect 18321 11056 18326 11112
rect 18382 11056 19338 11112
rect 19394 11056 19399 11112
rect 18321 11054 19399 11056
rect 18321 11051 18387 11054
rect 19333 11051 19399 11054
rect 7966 10916 7972 10980
rect 8036 10978 8042 10980
rect 11605 10978 11671 10981
rect 8036 10976 11671 10978
rect 8036 10920 11610 10976
rect 11666 10920 11671 10976
rect 8036 10918 11671 10920
rect 8036 10916 8042 10918
rect 11605 10915 11671 10918
rect 12065 10978 12131 10981
rect 12801 10978 12867 10981
rect 12065 10976 12867 10978
rect 12065 10920 12070 10976
rect 12126 10920 12806 10976
rect 12862 10920 12867 10976
rect 12065 10918 12867 10920
rect 12065 10915 12131 10918
rect 12801 10915 12867 10918
rect 16941 10978 17007 10981
rect 17125 10978 17191 10981
rect 16941 10976 17191 10978
rect 16941 10920 16946 10976
rect 17002 10920 17130 10976
rect 17186 10920 17191 10976
rect 16941 10918 17191 10920
rect 16941 10915 17007 10918
rect 17125 10915 17191 10918
rect 1354 10912 1750 10913
rect 1354 10848 1360 10912
rect 1424 10848 1440 10912
rect 1504 10848 1520 10912
rect 1584 10848 1600 10912
rect 1664 10848 1680 10912
rect 1744 10848 1750 10912
rect 1354 10847 1750 10848
rect 7354 10912 7750 10913
rect 7354 10848 7360 10912
rect 7424 10848 7440 10912
rect 7504 10848 7520 10912
rect 7584 10848 7600 10912
rect 7664 10848 7680 10912
rect 7744 10848 7750 10912
rect 7354 10847 7750 10848
rect 13354 10912 13750 10913
rect 13354 10848 13360 10912
rect 13424 10848 13440 10912
rect 13504 10848 13520 10912
rect 13584 10848 13600 10912
rect 13664 10848 13680 10912
rect 13744 10848 13750 10912
rect 13354 10847 13750 10848
rect 19354 10912 19750 10913
rect 19354 10848 19360 10912
rect 19424 10848 19440 10912
rect 19504 10848 19520 10912
rect 19584 10848 19600 10912
rect 19664 10848 19680 10912
rect 19744 10848 19750 10912
rect 19354 10847 19750 10848
rect 9121 10842 9187 10845
rect 13077 10842 13143 10845
rect 17769 10842 17835 10845
rect 9121 10840 13143 10842
rect 9121 10784 9126 10840
rect 9182 10784 13082 10840
rect 13138 10784 13143 10840
rect 9121 10782 13143 10784
rect 9121 10779 9187 10782
rect 13077 10779 13143 10782
rect 17726 10840 17835 10842
rect 17726 10784 17774 10840
rect 17830 10784 17835 10840
rect 17726 10779 17835 10784
rect 6545 10706 6611 10709
rect 6678 10706 6684 10708
rect 6545 10704 6684 10706
rect 6545 10648 6550 10704
rect 6606 10648 6684 10704
rect 6545 10646 6684 10648
rect 6545 10643 6611 10646
rect 6678 10644 6684 10646
rect 6748 10644 6754 10708
rect 8201 10706 8267 10709
rect 17585 10706 17651 10709
rect 17726 10706 17786 10779
rect 19241 10708 19307 10709
rect 19190 10706 19196 10708
rect 8201 10704 17786 10706
rect 8201 10648 8206 10704
rect 8262 10648 17590 10704
rect 17646 10648 17786 10704
rect 8201 10646 17786 10648
rect 19150 10646 19196 10706
rect 19260 10704 19307 10708
rect 19302 10648 19307 10704
rect 8201 10643 8267 10646
rect 17585 10643 17651 10646
rect 19190 10644 19196 10646
rect 19260 10644 19307 10648
rect 19241 10643 19307 10644
rect 8753 10570 8819 10573
rect 12249 10570 12315 10573
rect 12382 10570 12388 10572
rect 8753 10568 10932 10570
rect 8753 10512 8758 10568
rect 8814 10512 10932 10568
rect 8753 10510 10932 10512
rect 8753 10507 8819 10510
rect 4354 10368 4750 10369
rect 4354 10304 4360 10368
rect 4424 10304 4440 10368
rect 4504 10304 4520 10368
rect 4584 10304 4600 10368
rect 4664 10304 4680 10368
rect 4744 10304 4750 10368
rect 4354 10303 4750 10304
rect 10354 10368 10750 10369
rect 10354 10304 10360 10368
rect 10424 10304 10440 10368
rect 10504 10304 10520 10368
rect 10584 10304 10600 10368
rect 10664 10304 10680 10368
rect 10744 10304 10750 10368
rect 10354 10303 10750 10304
rect 9029 10298 9095 10301
rect 4846 10296 9095 10298
rect 4846 10240 9034 10296
rect 9090 10240 9095 10296
rect 4846 10238 9095 10240
rect 10872 10298 10932 10510
rect 12249 10568 12388 10570
rect 12249 10512 12254 10568
rect 12310 10512 12388 10568
rect 12249 10510 12388 10512
rect 12249 10507 12315 10510
rect 12382 10508 12388 10510
rect 12452 10508 12458 10572
rect 13118 10508 13124 10572
rect 13188 10570 13194 10572
rect 13445 10570 13511 10573
rect 13188 10568 13511 10570
rect 13188 10512 13450 10568
rect 13506 10512 13511 10568
rect 13188 10510 13511 10512
rect 13188 10508 13194 10510
rect 13445 10507 13511 10510
rect 14825 10570 14891 10573
rect 18229 10570 18295 10573
rect 19609 10570 19675 10573
rect 14825 10568 19675 10570
rect 14825 10512 14830 10568
rect 14886 10512 18234 10568
rect 18290 10512 19614 10568
rect 19670 10512 19675 10568
rect 14825 10510 19675 10512
rect 14825 10507 14891 10510
rect 18229 10507 18295 10510
rect 19609 10507 19675 10510
rect 12249 10434 12315 10437
rect 14641 10434 14707 10437
rect 12249 10432 14707 10434
rect 12249 10376 12254 10432
rect 12310 10376 14646 10432
rect 14702 10376 14707 10432
rect 12249 10374 14707 10376
rect 12249 10371 12315 10374
rect 14641 10371 14707 10374
rect 16354 10368 16750 10369
rect 16354 10304 16360 10368
rect 16424 10304 16440 10368
rect 16504 10304 16520 10368
rect 16584 10304 16600 10368
rect 16664 10304 16680 10368
rect 16744 10304 16750 10368
rect 16354 10303 16750 10304
rect 22354 10368 22750 10369
rect 22354 10304 22360 10368
rect 22424 10304 22440 10368
rect 22504 10304 22520 10368
rect 22584 10304 22600 10368
rect 22664 10304 22680 10368
rect 22744 10304 22750 10368
rect 22354 10303 22750 10304
rect 13629 10298 13695 10301
rect 10872 10296 13695 10298
rect 10872 10240 13634 10296
rect 13690 10240 13695 10296
rect 10872 10238 13695 10240
rect 4337 10162 4403 10165
rect 4846 10162 4906 10238
rect 9029 10235 9095 10238
rect 13629 10235 13695 10238
rect 17769 10298 17835 10301
rect 21725 10298 21791 10301
rect 17769 10296 21791 10298
rect 17769 10240 17774 10296
rect 17830 10240 21730 10296
rect 21786 10240 21791 10296
rect 17769 10238 21791 10240
rect 17769 10235 17835 10238
rect 21725 10235 21791 10238
rect 4337 10160 4906 10162
rect 4337 10104 4342 10160
rect 4398 10104 4906 10160
rect 4337 10102 4906 10104
rect 6729 10162 6795 10165
rect 16113 10162 16179 10165
rect 21449 10162 21515 10165
rect 6729 10160 16179 10162
rect 6729 10104 6734 10160
rect 6790 10104 16118 10160
rect 16174 10104 16179 10160
rect 6729 10102 16179 10104
rect 4337 10099 4403 10102
rect 6729 10099 6795 10102
rect 16113 10099 16179 10102
rect 16254 10160 21515 10162
rect 16254 10104 21454 10160
rect 21510 10104 21515 10160
rect 16254 10102 21515 10104
rect 6913 10026 6979 10029
rect 8201 10026 8267 10029
rect 6913 10024 8267 10026
rect 6913 9968 6918 10024
rect 6974 9968 8206 10024
rect 8262 9968 8267 10024
rect 6913 9966 8267 9968
rect 6913 9963 6979 9966
rect 8201 9963 8267 9966
rect 9213 10026 9279 10029
rect 14273 10026 14339 10029
rect 16254 10026 16314 10102
rect 21449 10099 21515 10102
rect 9213 10024 16314 10026
rect 9213 9968 9218 10024
rect 9274 9968 14278 10024
rect 14334 9968 16314 10024
rect 9213 9966 16314 9968
rect 16389 10026 16455 10029
rect 18597 10026 18663 10029
rect 16389 10024 18663 10026
rect 16389 9968 16394 10024
rect 16450 9968 18602 10024
rect 18658 9968 18663 10024
rect 16389 9966 18663 9968
rect 9213 9963 9279 9966
rect 14273 9963 14339 9966
rect 16389 9963 16455 9966
rect 18597 9963 18663 9966
rect 18822 9964 18828 10028
rect 18892 10026 18898 10028
rect 19926 10026 19932 10028
rect 18892 9966 19932 10026
rect 18892 9964 18898 9966
rect 19926 9964 19932 9966
rect 19996 9964 20002 10028
rect 10041 9890 10107 9893
rect 9998 9888 10107 9890
rect 9998 9832 10046 9888
rect 10102 9832 10107 9888
rect 9998 9827 10107 9832
rect 14825 9890 14891 9893
rect 18413 9890 18479 9893
rect 14825 9888 18479 9890
rect 14825 9832 14830 9888
rect 14886 9832 18418 9888
rect 18474 9832 18479 9888
rect 14825 9830 18479 9832
rect 14825 9827 14891 9830
rect 18413 9827 18479 9830
rect 1354 9824 1750 9825
rect 1354 9760 1360 9824
rect 1424 9760 1440 9824
rect 1504 9760 1520 9824
rect 1584 9760 1600 9824
rect 1664 9760 1680 9824
rect 1744 9760 1750 9824
rect 1354 9759 1750 9760
rect 7354 9824 7750 9825
rect 7354 9760 7360 9824
rect 7424 9760 7440 9824
rect 7504 9760 7520 9824
rect 7584 9760 7600 9824
rect 7664 9760 7680 9824
rect 7744 9760 7750 9824
rect 7354 9759 7750 9760
rect 9121 9754 9187 9757
rect 9622 9754 9628 9756
rect 9121 9752 9628 9754
rect 9121 9696 9126 9752
rect 9182 9696 9628 9752
rect 9121 9694 9628 9696
rect 9121 9691 9187 9694
rect 9622 9692 9628 9694
rect 9692 9692 9698 9756
rect 9857 9754 9923 9757
rect 9998 9754 10058 9827
rect 13354 9824 13750 9825
rect 13354 9760 13360 9824
rect 13424 9760 13440 9824
rect 13504 9760 13520 9824
rect 13584 9760 13600 9824
rect 13664 9760 13680 9824
rect 13744 9760 13750 9824
rect 13354 9759 13750 9760
rect 19354 9824 19750 9825
rect 19354 9760 19360 9824
rect 19424 9760 19440 9824
rect 19504 9760 19520 9824
rect 19584 9760 19600 9824
rect 19664 9760 19680 9824
rect 19744 9760 19750 9824
rect 19354 9759 19750 9760
rect 9857 9752 10058 9754
rect 9857 9696 9862 9752
rect 9918 9696 10058 9752
rect 9857 9694 10058 9696
rect 11053 9754 11119 9757
rect 12525 9754 12591 9757
rect 11053 9752 12591 9754
rect 11053 9696 11058 9752
rect 11114 9696 12530 9752
rect 12586 9696 12591 9752
rect 11053 9694 12591 9696
rect 9857 9691 9923 9694
rect 11053 9691 11119 9694
rect 12525 9691 12591 9694
rect 15285 9754 15351 9757
rect 15929 9754 15995 9757
rect 16757 9754 16823 9757
rect 18229 9756 18295 9757
rect 18229 9754 18276 9756
rect 15285 9752 15995 9754
rect 15285 9696 15290 9752
rect 15346 9696 15934 9752
rect 15990 9696 15995 9752
rect 15285 9694 15995 9696
rect 15285 9691 15351 9694
rect 15929 9691 15995 9694
rect 16438 9752 16823 9754
rect 16438 9696 16762 9752
rect 16818 9696 16823 9752
rect 16438 9694 16823 9696
rect 18184 9752 18276 9754
rect 18184 9696 18234 9752
rect 18184 9694 18276 9696
rect 16438 9621 16498 9694
rect 16757 9691 16823 9694
rect 18229 9692 18276 9694
rect 18340 9692 18346 9756
rect 18229 9691 18295 9692
rect 4061 9618 4127 9621
rect 9305 9618 9371 9621
rect 4061 9616 9371 9618
rect 4061 9560 4066 9616
rect 4122 9560 9310 9616
rect 9366 9560 9371 9616
rect 4061 9558 9371 9560
rect 4061 9555 4127 9558
rect 9305 9555 9371 9558
rect 13118 9556 13124 9620
rect 13188 9618 13194 9620
rect 16389 9618 16498 9621
rect 13188 9616 16498 9618
rect 13188 9560 16394 9616
rect 16450 9560 16498 9616
rect 13188 9558 16498 9560
rect 16757 9618 16823 9621
rect 21081 9618 21147 9621
rect 16757 9616 21147 9618
rect 16757 9560 16762 9616
rect 16818 9560 21086 9616
rect 21142 9560 21147 9616
rect 16757 9558 21147 9560
rect 13188 9556 13194 9558
rect 16389 9555 16455 9558
rect 16757 9555 16823 9558
rect 21081 9555 21147 9558
rect 1393 9482 1459 9485
rect 3325 9482 3391 9485
rect 1393 9480 3391 9482
rect 1393 9424 1398 9480
rect 1454 9424 3330 9480
rect 3386 9424 3391 9480
rect 1393 9422 3391 9424
rect 1393 9419 1459 9422
rect 3325 9419 3391 9422
rect 3601 9482 3667 9485
rect 9489 9482 9555 9485
rect 3601 9480 9555 9482
rect 3601 9424 3606 9480
rect 3662 9424 9494 9480
rect 9550 9424 9555 9480
rect 3601 9422 9555 9424
rect 3601 9419 3667 9422
rect 9489 9419 9555 9422
rect 10317 9482 10383 9485
rect 12525 9482 12591 9485
rect 16665 9482 16731 9485
rect 17861 9482 17927 9485
rect 19425 9482 19491 9485
rect 19885 9482 19951 9485
rect 10317 9480 12591 9482
rect 10317 9424 10322 9480
rect 10378 9424 12530 9480
rect 12586 9424 12591 9480
rect 10317 9422 12591 9424
rect 10317 9419 10383 9422
rect 12525 9419 12591 9422
rect 16070 9480 17786 9482
rect 16070 9424 16670 9480
rect 16726 9424 17786 9480
rect 16070 9422 17786 9424
rect 10869 9346 10935 9349
rect 15101 9346 15167 9349
rect 10869 9344 15167 9346
rect 10869 9288 10874 9344
rect 10930 9288 15106 9344
rect 15162 9288 15167 9344
rect 10869 9286 15167 9288
rect 10869 9283 10935 9286
rect 15101 9283 15167 9286
rect 4354 9280 4750 9281
rect 4354 9216 4360 9280
rect 4424 9216 4440 9280
rect 4504 9216 4520 9280
rect 4584 9216 4600 9280
rect 4664 9216 4680 9280
rect 4744 9216 4750 9280
rect 4354 9215 4750 9216
rect 10354 9280 10750 9281
rect 10354 9216 10360 9280
rect 10424 9216 10440 9280
rect 10504 9216 10520 9280
rect 10584 9216 10600 9280
rect 10664 9216 10680 9280
rect 10744 9216 10750 9280
rect 10354 9215 10750 9216
rect 1577 9210 1643 9213
rect 1945 9210 2011 9213
rect 3969 9210 4035 9213
rect 1577 9208 4035 9210
rect 1577 9152 1582 9208
rect 1638 9152 1950 9208
rect 2006 9152 3974 9208
rect 4030 9152 4035 9208
rect 1577 9150 4035 9152
rect 1577 9147 1643 9150
rect 1945 9147 2011 9150
rect 3969 9147 4035 9150
rect 7046 9148 7052 9212
rect 7116 9210 7122 9212
rect 7649 9210 7715 9213
rect 7116 9208 7715 9210
rect 7116 9152 7654 9208
rect 7710 9152 7715 9208
rect 7116 9150 7715 9152
rect 7116 9148 7122 9150
rect 7649 9147 7715 9150
rect 10910 9148 10916 9212
rect 10980 9210 10986 9212
rect 11145 9210 11211 9213
rect 10980 9208 11211 9210
rect 10980 9152 11150 9208
rect 11206 9152 11211 9208
rect 10980 9150 11211 9152
rect 10980 9148 10986 9150
rect 11145 9147 11211 9150
rect 11513 9210 11579 9213
rect 11697 9210 11763 9213
rect 12801 9210 12867 9213
rect 11513 9208 12867 9210
rect 11513 9152 11518 9208
rect 11574 9152 11702 9208
rect 11758 9152 12806 9208
rect 12862 9152 12867 9208
rect 11513 9150 12867 9152
rect 11513 9147 11579 9150
rect 11697 9147 11763 9150
rect 12801 9147 12867 9150
rect 13813 9210 13879 9213
rect 15285 9210 15351 9213
rect 13813 9208 15351 9210
rect 13813 9152 13818 9208
rect 13874 9152 15290 9208
rect 15346 9152 15351 9208
rect 13813 9150 15351 9152
rect 13813 9147 13879 9150
rect 15285 9147 15351 9150
rect 5349 9074 5415 9077
rect 6269 9074 6335 9077
rect 6545 9074 6611 9077
rect 14457 9074 14523 9077
rect 5349 9072 5642 9074
rect 5349 9016 5354 9072
rect 5410 9016 5642 9072
rect 5349 9014 5642 9016
rect 5349 9011 5415 9014
rect 5582 8941 5642 9014
rect 6269 9072 14523 9074
rect 6269 9016 6274 9072
rect 6330 9016 6550 9072
rect 6606 9016 14462 9072
rect 14518 9016 14523 9072
rect 6269 9014 14523 9016
rect 6269 9011 6335 9014
rect 6545 9011 6611 9014
rect 14457 9011 14523 9014
rect 14958 9012 14964 9076
rect 15028 9074 15034 9076
rect 15101 9074 15167 9077
rect 15028 9072 15167 9074
rect 15028 9016 15106 9072
rect 15162 9016 15167 9072
rect 15028 9014 15167 9016
rect 15028 9012 15034 9014
rect 15101 9011 15167 9014
rect 5582 8936 5691 8941
rect 5582 8880 5630 8936
rect 5686 8880 5691 8936
rect 5582 8878 5691 8880
rect 5625 8875 5691 8878
rect 7097 8938 7163 8941
rect 8109 8938 8175 8941
rect 16070 8938 16130 9422
rect 16665 9419 16731 9422
rect 17726 9346 17786 9422
rect 17861 9480 19350 9482
rect 17861 9424 17866 9480
rect 17922 9424 19350 9480
rect 17861 9422 19350 9424
rect 17861 9419 17927 9422
rect 18781 9346 18847 9349
rect 17726 9344 18847 9346
rect 17726 9288 18786 9344
rect 18842 9288 18847 9344
rect 17726 9286 18847 9288
rect 19290 9346 19350 9422
rect 19425 9480 19951 9482
rect 19425 9424 19430 9480
rect 19486 9424 19890 9480
rect 19946 9424 19951 9480
rect 19425 9422 19951 9424
rect 19425 9419 19491 9422
rect 19885 9419 19951 9422
rect 20069 9480 20135 9485
rect 20069 9424 20074 9480
rect 20130 9424 20135 9480
rect 20069 9419 20135 9424
rect 20072 9346 20132 9419
rect 20345 9346 20411 9349
rect 19290 9344 20411 9346
rect 19290 9288 20350 9344
rect 20406 9288 20411 9344
rect 19290 9286 20411 9288
rect 18781 9283 18847 9286
rect 20345 9283 20411 9286
rect 16354 9280 16750 9281
rect 16354 9216 16360 9280
rect 16424 9216 16440 9280
rect 16504 9216 16520 9280
rect 16584 9216 16600 9280
rect 16664 9216 16680 9280
rect 16744 9216 16750 9280
rect 16354 9215 16750 9216
rect 22354 9280 22750 9281
rect 22354 9216 22360 9280
rect 22424 9216 22440 9280
rect 22504 9216 22520 9280
rect 22584 9216 22600 9280
rect 22664 9216 22680 9280
rect 22744 9216 22750 9280
rect 22354 9215 22750 9216
rect 17309 9210 17375 9213
rect 17677 9210 17743 9213
rect 17309 9208 17743 9210
rect 17309 9152 17314 9208
rect 17370 9152 17682 9208
rect 17738 9152 17743 9208
rect 17309 9150 17743 9152
rect 17309 9147 17375 9150
rect 17677 9147 17743 9150
rect 18137 9210 18203 9213
rect 19333 9210 19399 9213
rect 20294 9210 20300 9212
rect 18137 9208 19258 9210
rect 18137 9152 18142 9208
rect 18198 9152 19258 9208
rect 18137 9150 19258 9152
rect 18137 9147 18203 9150
rect 17125 9074 17191 9077
rect 18137 9074 18203 9077
rect 19057 9074 19123 9077
rect 17125 9072 19123 9074
rect 17125 9016 17130 9072
rect 17186 9016 18142 9072
rect 18198 9016 19062 9072
rect 19118 9016 19123 9072
rect 17125 9014 19123 9016
rect 19198 9074 19258 9150
rect 19333 9208 20300 9210
rect 19333 9152 19338 9208
rect 19394 9152 20300 9208
rect 19333 9150 20300 9152
rect 19333 9147 19399 9150
rect 20294 9148 20300 9150
rect 20364 9148 20370 9212
rect 21449 9074 21515 9077
rect 19198 9072 21515 9074
rect 19198 9016 21454 9072
rect 21510 9016 21515 9072
rect 19198 9014 21515 9016
rect 17125 9011 17191 9014
rect 18137 9011 18203 9014
rect 19057 9011 19123 9014
rect 21449 9011 21515 9014
rect 18229 8940 18295 8941
rect 18229 8938 18276 8940
rect 7097 8936 16130 8938
rect 7097 8880 7102 8936
rect 7158 8880 8114 8936
rect 8170 8880 16130 8936
rect 7097 8878 16130 8880
rect 18184 8936 18276 8938
rect 18184 8880 18234 8936
rect 18184 8878 18276 8880
rect 7097 8875 7163 8878
rect 8109 8875 8175 8878
rect 18229 8876 18276 8878
rect 18340 8876 18346 8940
rect 19241 8938 19307 8941
rect 19701 8938 19767 8941
rect 19241 8936 19767 8938
rect 19241 8880 19246 8936
rect 19302 8880 19706 8936
rect 19762 8880 19767 8936
rect 19241 8878 19767 8880
rect 18229 8875 18295 8876
rect 19241 8875 19307 8878
rect 19701 8875 19767 8878
rect 7833 8802 7899 8805
rect 13118 8802 13124 8804
rect 7833 8800 13124 8802
rect 7833 8744 7838 8800
rect 7894 8744 13124 8800
rect 7833 8742 13124 8744
rect 7833 8739 7899 8742
rect 13118 8740 13124 8742
rect 13188 8740 13194 8804
rect 15101 8802 15167 8805
rect 18965 8802 19031 8805
rect 15101 8800 19031 8802
rect 15101 8744 15106 8800
rect 15162 8744 18970 8800
rect 19026 8744 19031 8800
rect 15101 8742 19031 8744
rect 15101 8739 15167 8742
rect 18965 8739 19031 8742
rect 1354 8736 1750 8737
rect 1354 8672 1360 8736
rect 1424 8672 1440 8736
rect 1504 8672 1520 8736
rect 1584 8672 1600 8736
rect 1664 8672 1680 8736
rect 1744 8672 1750 8736
rect 1354 8671 1750 8672
rect 7354 8736 7750 8737
rect 7354 8672 7360 8736
rect 7424 8672 7440 8736
rect 7504 8672 7520 8736
rect 7584 8672 7600 8736
rect 7664 8672 7680 8736
rect 7744 8672 7750 8736
rect 7354 8671 7750 8672
rect 13354 8736 13750 8737
rect 13354 8672 13360 8736
rect 13424 8672 13440 8736
rect 13504 8672 13520 8736
rect 13584 8672 13600 8736
rect 13664 8672 13680 8736
rect 13744 8672 13750 8736
rect 13354 8671 13750 8672
rect 19354 8736 19750 8737
rect 19354 8672 19360 8736
rect 19424 8672 19440 8736
rect 19504 8672 19520 8736
rect 19584 8672 19600 8736
rect 19664 8672 19680 8736
rect 19744 8672 19750 8736
rect 19354 8671 19750 8672
rect 2313 8666 2379 8669
rect 4797 8666 4863 8669
rect 5717 8668 5783 8669
rect 5717 8666 5764 8668
rect 2313 8664 4863 8666
rect 2313 8608 2318 8664
rect 2374 8608 4802 8664
rect 4858 8608 4863 8664
rect 2313 8606 4863 8608
rect 5672 8664 5764 8666
rect 5672 8608 5722 8664
rect 5672 8606 5764 8608
rect 2313 8603 2379 8606
rect 4797 8603 4863 8606
rect 5717 8604 5764 8606
rect 5828 8604 5834 8668
rect 9254 8604 9260 8668
rect 9324 8666 9330 8668
rect 9581 8666 9647 8669
rect 9324 8664 9647 8666
rect 9324 8608 9586 8664
rect 9642 8608 9647 8664
rect 9324 8606 9647 8608
rect 9324 8604 9330 8606
rect 5717 8603 5826 8604
rect 9581 8603 9647 8606
rect 15653 8666 15719 8669
rect 17585 8666 17651 8669
rect 15653 8664 17651 8666
rect 15653 8608 15658 8664
rect 15714 8608 17590 8664
rect 17646 8608 17651 8664
rect 15653 8606 17651 8608
rect 15653 8603 15719 8606
rect 17585 8603 17651 8606
rect 17861 8666 17927 8669
rect 18086 8666 18092 8668
rect 17861 8664 18092 8666
rect 17861 8608 17866 8664
rect 17922 8608 18092 8664
rect 17861 8606 18092 8608
rect 17861 8603 17927 8606
rect 18086 8604 18092 8606
rect 18156 8604 18162 8668
rect 18413 8666 18479 8669
rect 18689 8666 18755 8669
rect 18413 8664 18755 8666
rect 18413 8608 18418 8664
rect 18474 8608 18694 8664
rect 18750 8608 18755 8664
rect 18413 8606 18755 8608
rect 18413 8603 18479 8606
rect 18689 8603 18755 8606
rect 3141 8394 3207 8397
rect 3785 8394 3851 8397
rect 3141 8392 3851 8394
rect 3141 8336 3146 8392
rect 3202 8336 3790 8392
rect 3846 8336 3851 8392
rect 3141 8334 3851 8336
rect 3141 8331 3207 8334
rect 3785 8331 3851 8334
rect 4889 8394 4955 8397
rect 5390 8394 5396 8396
rect 4889 8392 5396 8394
rect 4889 8336 4894 8392
rect 4950 8336 5396 8392
rect 4889 8334 5396 8336
rect 4889 8331 4955 8334
rect 5390 8332 5396 8334
rect 5460 8332 5466 8396
rect 5766 8394 5826 8603
rect 8661 8530 8727 8533
rect 14917 8530 14983 8533
rect 8661 8528 14983 8530
rect 8661 8472 8666 8528
rect 8722 8472 14922 8528
rect 14978 8472 14983 8528
rect 8661 8470 14983 8472
rect 8661 8467 8727 8470
rect 14917 8467 14983 8470
rect 15101 8530 15167 8533
rect 21081 8530 21147 8533
rect 15101 8528 21147 8530
rect 15101 8472 15106 8528
rect 15162 8472 21086 8528
rect 21142 8472 21147 8528
rect 15101 8470 21147 8472
rect 15101 8467 15167 8470
rect 21081 8467 21147 8470
rect 9765 8394 9831 8397
rect 10317 8394 10383 8397
rect 5766 8334 9322 8394
rect 9262 8261 9322 8334
rect 9765 8392 10383 8394
rect 9765 8336 9770 8392
rect 9826 8336 10322 8392
rect 10378 8336 10383 8392
rect 9765 8334 10383 8336
rect 9765 8331 9831 8334
rect 10317 8331 10383 8334
rect 11605 8394 11671 8397
rect 15469 8394 15535 8397
rect 22829 8394 22895 8397
rect 11605 8392 22895 8394
rect 11605 8336 11610 8392
rect 11666 8336 15474 8392
rect 15530 8336 22834 8392
rect 22890 8336 22895 8392
rect 11605 8334 22895 8336
rect 11605 8331 11671 8334
rect 15469 8331 15535 8334
rect 22829 8331 22895 8334
rect 9262 8256 9371 8261
rect 9262 8200 9310 8256
rect 9366 8200 9371 8256
rect 9262 8198 9371 8200
rect 9305 8195 9371 8198
rect 12566 8196 12572 8260
rect 12636 8258 12642 8260
rect 15142 8258 15148 8260
rect 12636 8198 15148 8258
rect 12636 8196 12642 8198
rect 15142 8196 15148 8198
rect 15212 8196 15218 8260
rect 17953 8258 18019 8261
rect 19149 8258 19215 8261
rect 17953 8256 19215 8258
rect 17953 8200 17958 8256
rect 18014 8200 19154 8256
rect 19210 8200 19215 8256
rect 17953 8198 19215 8200
rect 17953 8195 18019 8198
rect 19149 8195 19215 8198
rect 4354 8192 4750 8193
rect 4354 8128 4360 8192
rect 4424 8128 4440 8192
rect 4504 8128 4520 8192
rect 4584 8128 4600 8192
rect 4664 8128 4680 8192
rect 4744 8128 4750 8192
rect 4354 8127 4750 8128
rect 10354 8192 10750 8193
rect 10354 8128 10360 8192
rect 10424 8128 10440 8192
rect 10504 8128 10520 8192
rect 10584 8128 10600 8192
rect 10664 8128 10680 8192
rect 10744 8128 10750 8192
rect 10354 8127 10750 8128
rect 16354 8192 16750 8193
rect 16354 8128 16360 8192
rect 16424 8128 16440 8192
rect 16504 8128 16520 8192
rect 16584 8128 16600 8192
rect 16664 8128 16680 8192
rect 16744 8128 16750 8192
rect 16354 8127 16750 8128
rect 22354 8192 22750 8193
rect 22354 8128 22360 8192
rect 22424 8128 22440 8192
rect 22504 8128 22520 8192
rect 22584 8128 22600 8192
rect 22664 8128 22680 8192
rect 22744 8128 22750 8192
rect 22354 8127 22750 8128
rect 12709 8122 12775 8125
rect 16021 8122 16087 8125
rect 12709 8120 16087 8122
rect 12709 8064 12714 8120
rect 12770 8064 16026 8120
rect 16082 8064 16087 8120
rect 12709 8062 16087 8064
rect 12709 8059 12775 8062
rect 16021 8059 16087 8062
rect 17493 8122 17559 8125
rect 17493 8120 18752 8122
rect 17493 8064 17498 8120
rect 17554 8064 18752 8120
rect 17493 8062 18752 8064
rect 17493 8059 17559 8062
rect 3141 7988 3207 7989
rect 3141 7986 3188 7988
rect 3096 7984 3188 7986
rect 3096 7928 3146 7984
rect 3096 7926 3188 7928
rect 3141 7924 3188 7926
rect 3252 7924 3258 7988
rect 6269 7986 6335 7989
rect 8385 7986 8451 7989
rect 6269 7984 8451 7986
rect 6269 7928 6274 7984
rect 6330 7928 8390 7984
rect 8446 7928 8451 7984
rect 6269 7926 8451 7928
rect 3141 7923 3207 7924
rect 6269 7923 6335 7926
rect 8385 7923 8451 7926
rect 8937 7986 9003 7989
rect 9254 7986 9260 7988
rect 8937 7984 9260 7986
rect 8937 7928 8942 7984
rect 8998 7928 9260 7984
rect 8937 7926 9260 7928
rect 8937 7923 9003 7926
rect 9254 7924 9260 7926
rect 9324 7986 9330 7988
rect 9581 7986 9647 7989
rect 9324 7984 9647 7986
rect 9324 7928 9586 7984
rect 9642 7928 9647 7984
rect 9324 7926 9647 7928
rect 9324 7924 9330 7926
rect 9581 7923 9647 7926
rect 10777 7986 10843 7989
rect 18413 7986 18479 7989
rect 10777 7984 18479 7986
rect 10777 7928 10782 7984
rect 10838 7928 18418 7984
rect 18474 7928 18479 7984
rect 10777 7926 18479 7928
rect 10777 7923 10843 7926
rect 18413 7923 18479 7926
rect 18692 7853 18752 8062
rect 7465 7850 7531 7853
rect 9121 7850 9187 7853
rect 17769 7850 17835 7853
rect 7465 7848 8218 7850
rect 7465 7792 7470 7848
rect 7526 7792 8218 7848
rect 7465 7790 8218 7792
rect 7465 7787 7531 7790
rect 1354 7648 1750 7649
rect 1354 7584 1360 7648
rect 1424 7584 1440 7648
rect 1504 7584 1520 7648
rect 1584 7584 1600 7648
rect 1664 7584 1680 7648
rect 1744 7584 1750 7648
rect 1354 7583 1750 7584
rect 7354 7648 7750 7649
rect 7354 7584 7360 7648
rect 7424 7584 7440 7648
rect 7504 7584 7520 7648
rect 7584 7584 7600 7648
rect 7664 7584 7680 7648
rect 7744 7584 7750 7648
rect 7354 7583 7750 7584
rect 6361 7442 6427 7445
rect 6729 7442 6795 7445
rect 6361 7440 6795 7442
rect 6361 7384 6366 7440
rect 6422 7384 6734 7440
rect 6790 7384 6795 7440
rect 6361 7382 6795 7384
rect 6361 7379 6427 7382
rect 6729 7379 6795 7382
rect 6545 7306 6611 7309
rect 8158 7306 8218 7790
rect 9121 7848 17835 7850
rect 9121 7792 9126 7848
rect 9182 7792 17774 7848
rect 17830 7792 17835 7848
rect 9121 7790 17835 7792
rect 9121 7787 9187 7790
rect 17769 7787 17835 7790
rect 18689 7848 18755 7853
rect 18689 7792 18694 7848
rect 18750 7792 18755 7848
rect 18689 7787 18755 7792
rect 14549 7714 14615 7717
rect 18965 7714 19031 7717
rect 14549 7712 19031 7714
rect 14549 7656 14554 7712
rect 14610 7656 18970 7712
rect 19026 7656 19031 7712
rect 14549 7654 19031 7656
rect 14549 7651 14615 7654
rect 18965 7651 19031 7654
rect 13354 7648 13750 7649
rect 13354 7584 13360 7648
rect 13424 7584 13440 7648
rect 13504 7584 13520 7648
rect 13584 7584 13600 7648
rect 13664 7584 13680 7648
rect 13744 7584 13750 7648
rect 13354 7583 13750 7584
rect 19354 7648 19750 7649
rect 19354 7584 19360 7648
rect 19424 7584 19440 7648
rect 19504 7584 19520 7648
rect 19584 7584 19600 7648
rect 19664 7584 19680 7648
rect 19744 7584 19750 7648
rect 19354 7583 19750 7584
rect 15561 7578 15627 7581
rect 18137 7578 18203 7581
rect 15561 7576 18203 7578
rect 15561 7520 15566 7576
rect 15622 7520 18142 7576
rect 18198 7520 18203 7576
rect 15561 7518 18203 7520
rect 15561 7515 15627 7518
rect 18137 7515 18203 7518
rect 8385 7442 8451 7445
rect 19241 7442 19307 7445
rect 8385 7440 19307 7442
rect 8385 7384 8390 7440
rect 8446 7384 19246 7440
rect 19302 7384 19307 7440
rect 8385 7382 19307 7384
rect 8385 7379 8451 7382
rect 19241 7379 19307 7382
rect 19609 7442 19675 7445
rect 20294 7442 20300 7444
rect 19609 7440 20300 7442
rect 19609 7384 19614 7440
rect 19670 7384 20300 7440
rect 19609 7382 20300 7384
rect 19609 7379 19675 7382
rect 20294 7380 20300 7382
rect 20364 7442 20370 7444
rect 21541 7442 21607 7445
rect 20364 7440 21607 7442
rect 20364 7384 21546 7440
rect 21602 7384 21607 7440
rect 20364 7382 21607 7384
rect 20364 7380 20370 7382
rect 21541 7379 21607 7382
rect 9673 7306 9739 7309
rect 6545 7304 6746 7306
rect 6545 7248 6550 7304
rect 6606 7248 6746 7304
rect 6545 7246 6746 7248
rect 8158 7304 9739 7306
rect 8158 7248 9678 7304
rect 9734 7248 9739 7304
rect 8158 7246 9739 7248
rect 6545 7243 6611 7246
rect 6686 7170 6746 7246
rect 9673 7243 9739 7246
rect 13629 7306 13695 7309
rect 13905 7306 13971 7309
rect 17493 7306 17559 7309
rect 13629 7304 17559 7306
rect 13629 7248 13634 7304
rect 13690 7248 13910 7304
rect 13966 7248 17498 7304
rect 17554 7248 17559 7304
rect 13629 7246 17559 7248
rect 13629 7243 13695 7246
rect 13905 7243 13971 7246
rect 17493 7243 17559 7246
rect 6821 7170 6887 7173
rect 6686 7168 6887 7170
rect 6686 7112 6826 7168
rect 6882 7112 6887 7168
rect 6686 7110 6887 7112
rect 6821 7107 6887 7110
rect 12014 7108 12020 7172
rect 12084 7170 12090 7172
rect 15561 7170 15627 7173
rect 12084 7168 15627 7170
rect 12084 7112 15566 7168
rect 15622 7112 15627 7168
rect 12084 7110 15627 7112
rect 12084 7108 12090 7110
rect 15561 7107 15627 7110
rect 4354 7104 4750 7105
rect 4354 7040 4360 7104
rect 4424 7040 4440 7104
rect 4504 7040 4520 7104
rect 4584 7040 4600 7104
rect 4664 7040 4680 7104
rect 4744 7040 4750 7104
rect 4354 7039 4750 7040
rect 10354 7104 10750 7105
rect 10354 7040 10360 7104
rect 10424 7040 10440 7104
rect 10504 7040 10520 7104
rect 10584 7040 10600 7104
rect 10664 7040 10680 7104
rect 10744 7040 10750 7104
rect 10354 7039 10750 7040
rect 16354 7104 16750 7105
rect 16354 7040 16360 7104
rect 16424 7040 16440 7104
rect 16504 7040 16520 7104
rect 16584 7040 16600 7104
rect 16664 7040 16680 7104
rect 16744 7040 16750 7104
rect 16354 7039 16750 7040
rect 22354 7104 22750 7105
rect 22354 7040 22360 7104
rect 22424 7040 22440 7104
rect 22504 7040 22520 7104
rect 22584 7040 22600 7104
rect 22664 7040 22680 7104
rect 22744 7040 22750 7104
rect 22354 7039 22750 7040
rect 5533 7034 5599 7037
rect 5942 7034 5948 7036
rect 5533 7032 5948 7034
rect 5533 6976 5538 7032
rect 5594 6976 5948 7032
rect 5533 6974 5948 6976
rect 5533 6971 5599 6974
rect 5942 6972 5948 6974
rect 6012 6972 6018 7036
rect 6453 7034 6519 7037
rect 6678 7034 6684 7036
rect 6453 7032 6684 7034
rect 6453 6976 6458 7032
rect 6514 6976 6684 7032
rect 6453 6974 6684 6976
rect 6453 6971 6519 6974
rect 6678 6972 6684 6974
rect 6748 6972 6754 7036
rect 11697 7034 11763 7037
rect 15377 7034 15443 7037
rect 10918 7032 11763 7034
rect 10918 6976 11702 7032
rect 11758 6976 11763 7032
rect 10918 6974 11763 6976
rect 10409 6898 10475 6901
rect 10918 6898 10978 6974
rect 11697 6971 11763 6974
rect 12758 7032 15443 7034
rect 12758 6976 15382 7032
rect 15438 6976 15443 7032
rect 12758 6974 15443 6976
rect 10409 6896 10978 6898
rect 10409 6840 10414 6896
rect 10470 6840 10978 6896
rect 10409 6838 10978 6840
rect 10409 6835 10475 6838
rect 11094 6836 11100 6900
rect 11164 6898 11170 6900
rect 12758 6898 12818 6974
rect 15377 6971 15443 6974
rect 11164 6838 12818 6898
rect 19793 6898 19859 6901
rect 20253 6898 20319 6901
rect 19793 6896 20319 6898
rect 19793 6840 19798 6896
rect 19854 6840 20258 6896
rect 20314 6840 20319 6896
rect 19793 6838 20319 6840
rect 11164 6836 11170 6838
rect 19793 6835 19859 6838
rect 20253 6835 20319 6838
rect 21909 6898 21975 6901
rect 22093 6898 22159 6901
rect 21909 6896 22159 6898
rect 21909 6840 21914 6896
rect 21970 6840 22098 6896
rect 22154 6840 22159 6896
rect 21909 6838 22159 6840
rect 21909 6835 21975 6838
rect 22093 6835 22159 6838
rect 6453 6762 6519 6765
rect 13905 6762 13971 6765
rect 6453 6760 13971 6762
rect 6453 6704 6458 6760
rect 6514 6704 13910 6760
rect 13966 6704 13971 6760
rect 6453 6702 13971 6704
rect 6453 6699 6519 6702
rect 13905 6699 13971 6702
rect 19701 6762 19767 6765
rect 19701 6760 21972 6762
rect 19701 6704 19706 6760
rect 19762 6704 21972 6760
rect 19701 6702 21972 6704
rect 19701 6699 19767 6702
rect 21912 6629 21972 6702
rect 8477 6626 8543 6629
rect 9029 6626 9095 6629
rect 8477 6624 9095 6626
rect 8477 6568 8482 6624
rect 8538 6568 9034 6624
rect 9090 6568 9095 6624
rect 8477 6566 9095 6568
rect 8477 6563 8543 6566
rect 9029 6563 9095 6566
rect 10501 6626 10567 6629
rect 11697 6626 11763 6629
rect 10501 6624 11763 6626
rect 10501 6568 10506 6624
rect 10562 6568 11702 6624
rect 11758 6568 11763 6624
rect 10501 6566 11763 6568
rect 10501 6563 10567 6566
rect 11697 6563 11763 6566
rect 21909 6624 21975 6629
rect 21909 6568 21914 6624
rect 21970 6568 21975 6624
rect 21909 6563 21975 6568
rect 1354 6560 1750 6561
rect 1354 6496 1360 6560
rect 1424 6496 1440 6560
rect 1504 6496 1520 6560
rect 1584 6496 1600 6560
rect 1664 6496 1680 6560
rect 1744 6496 1750 6560
rect 1354 6495 1750 6496
rect 7354 6560 7750 6561
rect 7354 6496 7360 6560
rect 7424 6496 7440 6560
rect 7504 6496 7520 6560
rect 7584 6496 7600 6560
rect 7664 6496 7680 6560
rect 7744 6496 7750 6560
rect 7354 6495 7750 6496
rect 13354 6560 13750 6561
rect 13354 6496 13360 6560
rect 13424 6496 13440 6560
rect 13504 6496 13520 6560
rect 13584 6496 13600 6560
rect 13664 6496 13680 6560
rect 13744 6496 13750 6560
rect 13354 6495 13750 6496
rect 19354 6560 19750 6561
rect 19354 6496 19360 6560
rect 19424 6496 19440 6560
rect 19504 6496 19520 6560
rect 19584 6496 19600 6560
rect 19664 6496 19680 6560
rect 19744 6496 19750 6560
rect 19354 6495 19750 6496
rect 7046 6428 7052 6492
rect 7116 6490 7122 6492
rect 7189 6490 7255 6493
rect 7116 6488 7255 6490
rect 7116 6432 7194 6488
rect 7250 6432 7255 6488
rect 7116 6430 7255 6432
rect 7116 6428 7122 6430
rect 7189 6427 7255 6430
rect 5942 6292 5948 6356
rect 6012 6354 6018 6356
rect 9213 6354 9279 6357
rect 6012 6352 9279 6354
rect 6012 6296 9218 6352
rect 9274 6296 9279 6352
rect 6012 6294 9279 6296
rect 6012 6292 6018 6294
rect 9213 6291 9279 6294
rect 9581 6354 9647 6357
rect 10869 6354 10935 6357
rect 9581 6352 10935 6354
rect 9581 6296 9586 6352
rect 9642 6296 10874 6352
rect 10930 6296 10935 6352
rect 9581 6294 10935 6296
rect 9581 6291 9647 6294
rect 10869 6291 10935 6294
rect 19425 6354 19491 6357
rect 19926 6354 19932 6356
rect 19425 6352 19932 6354
rect 19425 6296 19430 6352
rect 19486 6296 19932 6352
rect 19425 6294 19932 6296
rect 19425 6291 19491 6294
rect 19926 6292 19932 6294
rect 19996 6292 20002 6356
rect 8109 6218 8175 6221
rect 16297 6218 16363 6221
rect 21357 6218 21423 6221
rect 8109 6216 21423 6218
rect 8109 6160 8114 6216
rect 8170 6160 16302 6216
rect 16358 6160 21362 6216
rect 21418 6160 21423 6216
rect 8109 6158 21423 6160
rect 8109 6155 8175 6158
rect 16297 6155 16363 6158
rect 21357 6155 21423 6158
rect 7741 6082 7807 6085
rect 10041 6082 10107 6085
rect 7741 6080 10107 6082
rect 7741 6024 7746 6080
rect 7802 6024 10046 6080
rect 10102 6024 10107 6080
rect 7741 6022 10107 6024
rect 7741 6019 7807 6022
rect 10041 6019 10107 6022
rect 12985 6082 13051 6085
rect 15193 6082 15259 6085
rect 15377 6082 15443 6085
rect 12985 6080 15443 6082
rect 12985 6024 12990 6080
rect 13046 6024 15198 6080
rect 15254 6024 15382 6080
rect 15438 6024 15443 6080
rect 12985 6022 15443 6024
rect 12985 6019 13051 6022
rect 15193 6019 15259 6022
rect 15377 6019 15443 6022
rect 4354 6016 4750 6017
rect 4354 5952 4360 6016
rect 4424 5952 4440 6016
rect 4504 5952 4520 6016
rect 4584 5952 4600 6016
rect 4664 5952 4680 6016
rect 4744 5952 4750 6016
rect 4354 5951 4750 5952
rect 10354 6016 10750 6017
rect 10354 5952 10360 6016
rect 10424 5952 10440 6016
rect 10504 5952 10520 6016
rect 10584 5952 10600 6016
rect 10664 5952 10680 6016
rect 10744 5952 10750 6016
rect 10354 5951 10750 5952
rect 16354 6016 16750 6017
rect 16354 5952 16360 6016
rect 16424 5952 16440 6016
rect 16504 5952 16520 6016
rect 16584 5952 16600 6016
rect 16664 5952 16680 6016
rect 16744 5952 16750 6016
rect 16354 5951 16750 5952
rect 22354 6016 22750 6017
rect 22354 5952 22360 6016
rect 22424 5952 22440 6016
rect 22504 5952 22520 6016
rect 22584 5952 22600 6016
rect 22664 5952 22680 6016
rect 22744 5952 22750 6016
rect 22354 5951 22750 5952
rect 9949 5946 10015 5949
rect 10174 5946 10180 5948
rect 9949 5944 10180 5946
rect 9949 5888 9954 5944
rect 10010 5888 10180 5944
rect 9949 5886 10180 5888
rect 9949 5883 10015 5886
rect 10174 5884 10180 5886
rect 10244 5884 10250 5948
rect 15694 5748 15700 5812
rect 15764 5810 15770 5812
rect 19517 5810 19583 5813
rect 15764 5808 19583 5810
rect 15764 5752 19522 5808
rect 19578 5752 19583 5808
rect 15764 5750 19583 5752
rect 15764 5748 15770 5750
rect 19517 5747 19583 5750
rect 3601 5674 3667 5677
rect 8109 5674 8175 5677
rect 3601 5672 8175 5674
rect 3601 5616 3606 5672
rect 3662 5616 8114 5672
rect 8170 5616 8175 5672
rect 3601 5614 8175 5616
rect 3601 5611 3667 5614
rect 8109 5611 8175 5614
rect 20069 5674 20135 5677
rect 20846 5674 20852 5676
rect 20069 5672 20852 5674
rect 20069 5616 20074 5672
rect 20130 5616 20852 5672
rect 20069 5614 20852 5616
rect 20069 5611 20135 5614
rect 20846 5612 20852 5614
rect 20916 5612 20922 5676
rect 7966 5476 7972 5540
rect 8036 5538 8042 5540
rect 8109 5538 8175 5541
rect 8036 5536 8175 5538
rect 8036 5480 8114 5536
rect 8170 5480 8175 5536
rect 8036 5478 8175 5480
rect 8036 5476 8042 5478
rect 8109 5475 8175 5478
rect 10041 5538 10107 5541
rect 10910 5538 10916 5540
rect 10041 5536 10916 5538
rect 10041 5480 10046 5536
rect 10102 5480 10916 5536
rect 10041 5478 10916 5480
rect 10041 5475 10107 5478
rect 10910 5476 10916 5478
rect 10980 5476 10986 5540
rect 1354 5472 1750 5473
rect 1354 5408 1360 5472
rect 1424 5408 1440 5472
rect 1504 5408 1520 5472
rect 1584 5408 1600 5472
rect 1664 5408 1680 5472
rect 1744 5408 1750 5472
rect 1354 5407 1750 5408
rect 7354 5472 7750 5473
rect 7354 5408 7360 5472
rect 7424 5408 7440 5472
rect 7504 5408 7520 5472
rect 7584 5408 7600 5472
rect 7664 5408 7680 5472
rect 7744 5408 7750 5472
rect 7354 5407 7750 5408
rect 13354 5472 13750 5473
rect 13354 5408 13360 5472
rect 13424 5408 13440 5472
rect 13504 5408 13520 5472
rect 13584 5408 13600 5472
rect 13664 5408 13680 5472
rect 13744 5408 13750 5472
rect 13354 5407 13750 5408
rect 19354 5472 19750 5473
rect 19354 5408 19360 5472
rect 19424 5408 19440 5472
rect 19504 5408 19520 5472
rect 19584 5408 19600 5472
rect 19664 5408 19680 5472
rect 19744 5408 19750 5472
rect 19354 5407 19750 5408
rect 10133 5402 10199 5405
rect 10133 5400 12450 5402
rect 10133 5344 10138 5400
rect 10194 5344 12450 5400
rect 10133 5342 12450 5344
rect 10133 5339 10199 5342
rect 9622 5204 9628 5268
rect 9692 5266 9698 5268
rect 11329 5266 11395 5269
rect 9692 5264 11395 5266
rect 9692 5208 11334 5264
rect 11390 5208 11395 5264
rect 9692 5206 11395 5208
rect 12390 5266 12450 5342
rect 12893 5266 12959 5269
rect 12390 5264 12959 5266
rect 12390 5208 12898 5264
rect 12954 5208 12959 5264
rect 12390 5206 12959 5208
rect 9692 5204 9698 5206
rect 11329 5203 11395 5206
rect 12893 5203 12959 5206
rect 15142 5204 15148 5268
rect 15212 5266 15218 5268
rect 17401 5266 17467 5269
rect 15212 5264 17467 5266
rect 15212 5208 17406 5264
rect 17462 5208 17467 5264
rect 15212 5206 17467 5208
rect 15212 5204 15218 5206
rect 17401 5203 17467 5206
rect 19006 5204 19012 5268
rect 19076 5266 19082 5268
rect 19701 5266 19767 5269
rect 19076 5264 19767 5266
rect 19076 5208 19706 5264
rect 19762 5208 19767 5264
rect 19076 5206 19767 5208
rect 19076 5204 19082 5206
rect 19701 5203 19767 5206
rect 4337 5130 4403 5133
rect 4110 5128 4403 5130
rect 4110 5072 4342 5128
rect 4398 5072 4403 5128
rect 4110 5070 4403 5072
rect 3693 4724 3759 4725
rect 3693 4722 3740 4724
rect 3648 4720 3740 4722
rect 3648 4664 3698 4720
rect 3648 4662 3740 4664
rect 3693 4660 3740 4662
rect 3804 4660 3810 4724
rect 4110 4722 4170 5070
rect 4337 5067 4403 5070
rect 12341 5130 12407 5133
rect 19149 5130 19215 5133
rect 12341 5128 19215 5130
rect 12341 5072 12346 5128
rect 12402 5072 19154 5128
rect 19210 5072 19215 5128
rect 12341 5070 19215 5072
rect 12341 5067 12407 5070
rect 19149 5067 19215 5070
rect 12249 4994 12315 4997
rect 12617 4994 12683 4997
rect 12249 4992 12683 4994
rect 12249 4936 12254 4992
rect 12310 4936 12622 4992
rect 12678 4936 12683 4992
rect 12249 4934 12683 4936
rect 12249 4931 12315 4934
rect 12617 4931 12683 4934
rect 4354 4928 4750 4929
rect 4354 4864 4360 4928
rect 4424 4864 4440 4928
rect 4504 4864 4520 4928
rect 4584 4864 4600 4928
rect 4664 4864 4680 4928
rect 4744 4864 4750 4928
rect 4354 4863 4750 4864
rect 10354 4928 10750 4929
rect 10354 4864 10360 4928
rect 10424 4864 10440 4928
rect 10504 4864 10520 4928
rect 10584 4864 10600 4928
rect 10664 4864 10680 4928
rect 10744 4864 10750 4928
rect 10354 4863 10750 4864
rect 16354 4928 16750 4929
rect 16354 4864 16360 4928
rect 16424 4864 16440 4928
rect 16504 4864 16520 4928
rect 16584 4864 16600 4928
rect 16664 4864 16680 4928
rect 16744 4864 16750 4928
rect 16354 4863 16750 4864
rect 22354 4928 22750 4929
rect 22354 4864 22360 4928
rect 22424 4864 22440 4928
rect 22504 4864 22520 4928
rect 22584 4864 22600 4928
rect 22664 4864 22680 4928
rect 22744 4864 22750 4928
rect 22354 4863 22750 4864
rect 12249 4858 12315 4861
rect 14917 4858 14983 4861
rect 12249 4856 14983 4858
rect 12249 4800 12254 4856
rect 12310 4800 14922 4856
rect 14978 4800 14983 4856
rect 12249 4798 14983 4800
rect 12249 4795 12315 4798
rect 14917 4795 14983 4798
rect 4337 4722 4403 4725
rect 4110 4720 4403 4722
rect 4110 4664 4342 4720
rect 4398 4664 4403 4720
rect 4110 4662 4403 4664
rect 3693 4659 3759 4660
rect 4337 4659 4403 4662
rect 11329 4722 11395 4725
rect 12893 4722 12959 4725
rect 11329 4720 12959 4722
rect 11329 4664 11334 4720
rect 11390 4664 12898 4720
rect 12954 4664 12959 4720
rect 11329 4662 12959 4664
rect 11329 4659 11395 4662
rect 12893 4659 12959 4662
rect 12893 4586 12959 4589
rect 18045 4586 18111 4589
rect 12893 4584 18111 4586
rect 12893 4528 12898 4584
rect 12954 4528 18050 4584
rect 18106 4528 18111 4584
rect 12893 4526 18111 4528
rect 12893 4523 12959 4526
rect 18045 4523 18111 4526
rect 1354 4384 1750 4385
rect 1354 4320 1360 4384
rect 1424 4320 1440 4384
rect 1504 4320 1520 4384
rect 1584 4320 1600 4384
rect 1664 4320 1680 4384
rect 1744 4320 1750 4384
rect 1354 4319 1750 4320
rect 7354 4384 7750 4385
rect 7354 4320 7360 4384
rect 7424 4320 7440 4384
rect 7504 4320 7520 4384
rect 7584 4320 7600 4384
rect 7664 4320 7680 4384
rect 7744 4320 7750 4384
rect 7354 4319 7750 4320
rect 13354 4384 13750 4385
rect 13354 4320 13360 4384
rect 13424 4320 13440 4384
rect 13504 4320 13520 4384
rect 13584 4320 13600 4384
rect 13664 4320 13680 4384
rect 13744 4320 13750 4384
rect 13354 4319 13750 4320
rect 19354 4384 19750 4385
rect 19354 4320 19360 4384
rect 19424 4320 19440 4384
rect 19504 4320 19520 4384
rect 19584 4320 19600 4384
rect 19664 4320 19680 4384
rect 19744 4320 19750 4384
rect 19354 4319 19750 4320
rect 14181 4314 14247 4317
rect 19057 4314 19123 4317
rect 14181 4312 19123 4314
rect 14181 4256 14186 4312
rect 14242 4256 19062 4312
rect 19118 4256 19123 4312
rect 14181 4254 19123 4256
rect 14181 4251 14247 4254
rect 19057 4251 19123 4254
rect 8017 4178 8083 4181
rect 9990 4178 9996 4180
rect 8017 4176 9996 4178
rect 8017 4120 8022 4176
rect 8078 4120 9996 4176
rect 8017 4118 9996 4120
rect 8017 4115 8083 4118
rect 9990 4116 9996 4118
rect 10060 4116 10066 4180
rect 15745 4178 15811 4181
rect 16297 4178 16363 4181
rect 15745 4176 16363 4178
rect 15745 4120 15750 4176
rect 15806 4120 16302 4176
rect 16358 4120 16363 4176
rect 15745 4118 16363 4120
rect 15745 4115 15811 4118
rect 16297 4115 16363 4118
rect 21081 4178 21147 4181
rect 21582 4178 21588 4180
rect 21081 4176 21588 4178
rect 21081 4120 21086 4176
rect 21142 4120 21588 4176
rect 21081 4118 21588 4120
rect 21081 4115 21147 4118
rect 21582 4116 21588 4118
rect 21652 4116 21658 4180
rect 3918 3980 3924 4044
rect 3988 4042 3994 4044
rect 4981 4042 5047 4045
rect 3988 4040 5047 4042
rect 3988 3984 4986 4040
rect 5042 3984 5047 4040
rect 3988 3982 5047 3984
rect 3988 3980 3994 3982
rect 4981 3979 5047 3982
rect 10041 4042 10107 4045
rect 10685 4042 10751 4045
rect 19977 4042 20043 4045
rect 10041 4040 20043 4042
rect 10041 3984 10046 4040
rect 10102 3984 10690 4040
rect 10746 3984 19982 4040
rect 20038 3984 20043 4040
rect 10041 3982 20043 3984
rect 10041 3979 10107 3982
rect 10685 3979 10751 3982
rect 19977 3979 20043 3982
rect 20253 4042 20319 4045
rect 21030 4042 21036 4044
rect 20253 4040 21036 4042
rect 20253 3984 20258 4040
rect 20314 3984 21036 4040
rect 20253 3982 21036 3984
rect 20253 3979 20319 3982
rect 21030 3980 21036 3982
rect 21100 3980 21106 4044
rect 4354 3840 4750 3841
rect 4354 3776 4360 3840
rect 4424 3776 4440 3840
rect 4504 3776 4520 3840
rect 4584 3776 4600 3840
rect 4664 3776 4680 3840
rect 4744 3776 4750 3840
rect 4354 3775 4750 3776
rect 10354 3840 10750 3841
rect 10354 3776 10360 3840
rect 10424 3776 10440 3840
rect 10504 3776 10520 3840
rect 10584 3776 10600 3840
rect 10664 3776 10680 3840
rect 10744 3776 10750 3840
rect 10354 3775 10750 3776
rect 16354 3840 16750 3841
rect 16354 3776 16360 3840
rect 16424 3776 16440 3840
rect 16504 3776 16520 3840
rect 16584 3776 16600 3840
rect 16664 3776 16680 3840
rect 16744 3776 16750 3840
rect 16354 3775 16750 3776
rect 22354 3840 22750 3841
rect 22354 3776 22360 3840
rect 22424 3776 22440 3840
rect 22504 3776 22520 3840
rect 22584 3776 22600 3840
rect 22664 3776 22680 3840
rect 22744 3776 22750 3840
rect 22354 3775 22750 3776
rect 9029 3634 9095 3637
rect 10501 3634 10567 3637
rect 9029 3632 10567 3634
rect 9029 3576 9034 3632
rect 9090 3576 10506 3632
rect 10562 3576 10567 3632
rect 9029 3574 10567 3576
rect 9029 3571 9095 3574
rect 10501 3571 10567 3574
rect 14089 3634 14155 3637
rect 19517 3634 19583 3637
rect 14089 3632 19583 3634
rect 14089 3576 14094 3632
rect 14150 3576 19522 3632
rect 19578 3576 19583 3632
rect 14089 3574 19583 3576
rect 14089 3571 14155 3574
rect 19517 3571 19583 3574
rect 19885 3634 19951 3637
rect 21081 3636 21147 3637
rect 20110 3634 20116 3636
rect 19885 3632 20116 3634
rect 19885 3576 19890 3632
rect 19946 3576 20116 3632
rect 19885 3574 20116 3576
rect 19885 3571 19951 3574
rect 20110 3572 20116 3574
rect 20180 3572 20186 3636
rect 21030 3572 21036 3636
rect 21100 3634 21147 3636
rect 21100 3632 21192 3634
rect 21142 3576 21192 3632
rect 21100 3574 21192 3576
rect 21100 3572 21147 3574
rect 21081 3571 21147 3572
rect 10225 3498 10291 3501
rect 11278 3498 11284 3500
rect 10225 3496 11284 3498
rect 10225 3440 10230 3496
rect 10286 3440 11284 3496
rect 10225 3438 11284 3440
rect 10225 3435 10291 3438
rect 11278 3436 11284 3438
rect 11348 3498 11354 3500
rect 18873 3498 18939 3501
rect 11348 3496 18939 3498
rect 11348 3440 18878 3496
rect 18934 3440 18939 3496
rect 11348 3438 18939 3440
rect 11348 3436 11354 3438
rect 18873 3435 18939 3438
rect 19333 3498 19399 3501
rect 21173 3498 21239 3501
rect 19333 3496 21239 3498
rect 19333 3440 19338 3496
rect 19394 3440 21178 3496
rect 21234 3440 21239 3496
rect 19333 3438 21239 3440
rect 19333 3435 19399 3438
rect 21173 3435 21239 3438
rect 10593 3362 10659 3365
rect 11513 3362 11579 3365
rect 10593 3360 11579 3362
rect 10593 3304 10598 3360
rect 10654 3304 11518 3360
rect 11574 3304 11579 3360
rect 10593 3302 11579 3304
rect 10593 3299 10659 3302
rect 11513 3299 11579 3302
rect 1354 3296 1750 3297
rect 1354 3232 1360 3296
rect 1424 3232 1440 3296
rect 1504 3232 1520 3296
rect 1584 3232 1600 3296
rect 1664 3232 1680 3296
rect 1744 3232 1750 3296
rect 1354 3231 1750 3232
rect 7354 3296 7750 3297
rect 7354 3232 7360 3296
rect 7424 3232 7440 3296
rect 7504 3232 7520 3296
rect 7584 3232 7600 3296
rect 7664 3232 7680 3296
rect 7744 3232 7750 3296
rect 7354 3231 7750 3232
rect 13354 3296 13750 3297
rect 13354 3232 13360 3296
rect 13424 3232 13440 3296
rect 13504 3232 13520 3296
rect 13584 3232 13600 3296
rect 13664 3232 13680 3296
rect 13744 3232 13750 3296
rect 13354 3231 13750 3232
rect 19354 3296 19750 3297
rect 19354 3232 19360 3296
rect 19424 3232 19440 3296
rect 19504 3232 19520 3296
rect 19584 3232 19600 3296
rect 19664 3232 19680 3296
rect 19744 3232 19750 3296
rect 19354 3231 19750 3232
rect 4981 3092 5047 3093
rect 4981 3090 5028 3092
rect 4936 3088 5028 3090
rect 4936 3032 4986 3088
rect 4936 3030 5028 3032
rect 4981 3028 5028 3030
rect 5092 3028 5098 3092
rect 7741 3090 7807 3093
rect 11094 3090 11100 3092
rect 7741 3088 11100 3090
rect 7741 3032 7746 3088
rect 7802 3032 11100 3088
rect 7741 3030 11100 3032
rect 4981 3027 5047 3028
rect 7741 3027 7807 3030
rect 11094 3028 11100 3030
rect 11164 3028 11170 3092
rect 11329 3090 11395 3093
rect 20345 3090 20411 3093
rect 11329 3088 20411 3090
rect 11329 3032 11334 3088
rect 11390 3032 20350 3088
rect 20406 3032 20411 3088
rect 11329 3030 20411 3032
rect 11329 3027 11395 3030
rect 20345 3027 20411 3030
rect 9581 2954 9647 2957
rect 14089 2954 14155 2957
rect 9581 2952 14155 2954
rect 9581 2896 9586 2952
rect 9642 2896 14094 2952
rect 14150 2896 14155 2952
rect 9581 2894 14155 2896
rect 9581 2891 9647 2894
rect 14089 2891 14155 2894
rect 10961 2820 11027 2821
rect 10910 2756 10916 2820
rect 10980 2818 11027 2820
rect 11605 2818 11671 2821
rect 12617 2818 12683 2821
rect 13721 2818 13787 2821
rect 10980 2816 11072 2818
rect 11022 2760 11072 2816
rect 10980 2758 11072 2760
rect 11605 2816 13787 2818
rect 11605 2760 11610 2816
rect 11666 2760 12622 2816
rect 12678 2760 13726 2816
rect 13782 2760 13787 2816
rect 11605 2758 13787 2760
rect 10980 2756 11027 2758
rect 10961 2755 11027 2756
rect 11605 2755 11671 2758
rect 12617 2755 12683 2758
rect 13721 2755 13787 2758
rect 4354 2752 4750 2753
rect 4354 2688 4360 2752
rect 4424 2688 4440 2752
rect 4504 2688 4520 2752
rect 4584 2688 4600 2752
rect 4664 2688 4680 2752
rect 4744 2688 4750 2752
rect 4354 2687 4750 2688
rect 10354 2752 10750 2753
rect 10354 2688 10360 2752
rect 10424 2688 10440 2752
rect 10504 2688 10520 2752
rect 10584 2688 10600 2752
rect 10664 2688 10680 2752
rect 10744 2688 10750 2752
rect 10354 2687 10750 2688
rect 16354 2752 16750 2753
rect 16354 2688 16360 2752
rect 16424 2688 16440 2752
rect 16504 2688 16520 2752
rect 16584 2688 16600 2752
rect 16664 2688 16680 2752
rect 16744 2688 16750 2752
rect 16354 2687 16750 2688
rect 22354 2752 22750 2753
rect 22354 2688 22360 2752
rect 22424 2688 22440 2752
rect 22504 2688 22520 2752
rect 22584 2688 22600 2752
rect 22664 2688 22680 2752
rect 22744 2688 22750 2752
rect 22354 2687 22750 2688
rect 11329 2682 11395 2685
rect 11881 2682 11947 2685
rect 18505 2682 18571 2685
rect 21817 2682 21883 2685
rect 11329 2680 15256 2682
rect 11329 2624 11334 2680
rect 11390 2624 11886 2680
rect 11942 2624 15256 2680
rect 11329 2622 15256 2624
rect 11329 2619 11395 2622
rect 11881 2619 11947 2622
rect 15196 2549 15256 2622
rect 18505 2680 21883 2682
rect 18505 2624 18510 2680
rect 18566 2624 21822 2680
rect 21878 2624 21883 2680
rect 18505 2622 21883 2624
rect 18505 2619 18571 2622
rect 21817 2619 21883 2622
rect 12433 2546 12499 2549
rect 15193 2546 15259 2549
rect 16297 2546 16363 2549
rect 12433 2544 15072 2546
rect 12433 2488 12438 2544
rect 12494 2488 15072 2544
rect 12433 2486 15072 2488
rect 12433 2483 12499 2486
rect 8293 2410 8359 2413
rect 10225 2412 10291 2413
rect 9438 2410 9444 2412
rect 8293 2408 9444 2410
rect 8293 2352 8298 2408
rect 8354 2352 9444 2408
rect 8293 2350 9444 2352
rect 8293 2347 8359 2350
rect 9438 2348 9444 2350
rect 9508 2348 9514 2412
rect 10174 2348 10180 2412
rect 10244 2410 10291 2412
rect 10961 2410 11027 2413
rect 10244 2408 11027 2410
rect 10286 2352 10966 2408
rect 11022 2352 11027 2408
rect 10244 2350 11027 2352
rect 10244 2348 10291 2350
rect 10225 2347 10291 2348
rect 10961 2347 11027 2350
rect 11237 2410 11303 2413
rect 14181 2410 14247 2413
rect 11237 2408 14247 2410
rect 11237 2352 11242 2408
rect 11298 2352 14186 2408
rect 14242 2352 14247 2408
rect 11237 2350 14247 2352
rect 15012 2410 15072 2486
rect 15193 2544 20776 2546
rect 15193 2488 15198 2544
rect 15254 2488 16302 2544
rect 16358 2488 20776 2544
rect 15193 2486 20776 2488
rect 15193 2483 15259 2486
rect 16297 2483 16363 2486
rect 17677 2410 17743 2413
rect 15012 2408 17743 2410
rect 15012 2352 17682 2408
rect 17738 2352 17743 2408
rect 15012 2350 17743 2352
rect 11237 2347 11303 2350
rect 14181 2347 14247 2350
rect 17677 2347 17743 2350
rect 17861 2410 17927 2413
rect 20069 2410 20135 2413
rect 17861 2408 20135 2410
rect 17861 2352 17866 2408
rect 17922 2352 20074 2408
rect 20130 2352 20135 2408
rect 17861 2350 20135 2352
rect 20716 2410 20776 2486
rect 22185 2410 22251 2413
rect 20716 2408 22251 2410
rect 20716 2352 22190 2408
rect 22246 2352 22251 2408
rect 20716 2350 22251 2352
rect 17861 2347 17927 2350
rect 20069 2347 20135 2350
rect 22185 2347 22251 2350
rect 9673 2274 9739 2277
rect 11881 2274 11947 2277
rect 12433 2274 12499 2277
rect 9673 2272 12499 2274
rect 9673 2216 9678 2272
rect 9734 2216 11886 2272
rect 11942 2216 12438 2272
rect 12494 2216 12499 2272
rect 9673 2214 12499 2216
rect 9673 2211 9739 2214
rect 11881 2211 11947 2214
rect 12433 2211 12499 2214
rect 14273 2274 14339 2277
rect 18045 2274 18111 2277
rect 14273 2272 18111 2274
rect 14273 2216 14278 2272
rect 14334 2216 18050 2272
rect 18106 2216 18111 2272
rect 14273 2214 18111 2216
rect 14273 2211 14339 2214
rect 18045 2211 18111 2214
rect 19885 2274 19951 2277
rect 22461 2274 22527 2277
rect 19885 2272 22527 2274
rect 19885 2216 19890 2272
rect 19946 2216 22466 2272
rect 22522 2216 22527 2272
rect 19885 2214 22527 2216
rect 19885 2211 19951 2214
rect 22461 2211 22527 2214
rect 1354 2208 1750 2209
rect 1354 2144 1360 2208
rect 1424 2144 1440 2208
rect 1504 2144 1520 2208
rect 1584 2144 1600 2208
rect 1664 2144 1680 2208
rect 1744 2144 1750 2208
rect 1354 2143 1750 2144
rect 7354 2208 7750 2209
rect 7354 2144 7360 2208
rect 7424 2144 7440 2208
rect 7504 2144 7520 2208
rect 7584 2144 7600 2208
rect 7664 2144 7680 2208
rect 7744 2144 7750 2208
rect 7354 2143 7750 2144
rect 13354 2208 13750 2209
rect 13354 2144 13360 2208
rect 13424 2144 13440 2208
rect 13504 2144 13520 2208
rect 13584 2144 13600 2208
rect 13664 2144 13680 2208
rect 13744 2144 13750 2208
rect 13354 2143 13750 2144
rect 19354 2208 19750 2209
rect 19354 2144 19360 2208
rect 19424 2144 19440 2208
rect 19504 2144 19520 2208
rect 19584 2144 19600 2208
rect 19664 2144 19680 2208
rect 19744 2144 19750 2208
rect 19354 2143 19750 2144
rect 9070 2076 9076 2140
rect 9140 2138 9146 2140
rect 9949 2138 10015 2141
rect 12157 2138 12223 2141
rect 13077 2138 13143 2141
rect 9140 2136 13143 2138
rect 9140 2080 9954 2136
rect 10010 2080 12162 2136
rect 12218 2080 13082 2136
rect 13138 2080 13143 2136
rect 9140 2078 13143 2080
rect 9140 2076 9146 2078
rect 9949 2075 10015 2078
rect 12157 2075 12223 2078
rect 13077 2075 13143 2078
rect 13813 2138 13879 2141
rect 13813 2136 18154 2138
rect 13813 2080 13818 2136
rect 13874 2080 18154 2136
rect 13813 2078 18154 2080
rect 13813 2075 13879 2078
rect 6494 1940 6500 2004
rect 6564 2002 6570 2004
rect 6637 2002 6703 2005
rect 6564 2000 6703 2002
rect 6564 1944 6642 2000
rect 6698 1944 6703 2000
rect 6564 1942 6703 1944
rect 6564 1940 6570 1942
rect 6637 1939 6703 1942
rect 9857 2002 9923 2005
rect 17769 2002 17835 2005
rect 9857 2000 17835 2002
rect 9857 1944 9862 2000
rect 9918 1944 17774 2000
rect 17830 1944 17835 2000
rect 9857 1942 17835 1944
rect 9857 1939 9923 1942
rect 17769 1939 17835 1942
rect 10041 1866 10107 1869
rect 12433 1866 12499 1869
rect 12617 1866 12683 1869
rect 10041 1864 12499 1866
rect 10041 1808 10046 1864
rect 10102 1808 12438 1864
rect 12494 1808 12499 1864
rect 10041 1806 12499 1808
rect 10041 1803 10107 1806
rect 12433 1803 12499 1806
rect 12574 1864 12683 1866
rect 12574 1808 12622 1864
rect 12678 1808 12683 1864
rect 12574 1803 12683 1808
rect 12801 1866 12867 1869
rect 14549 1866 14615 1869
rect 12801 1864 14615 1866
rect 12801 1808 12806 1864
rect 12862 1808 14554 1864
rect 14610 1808 14615 1864
rect 12801 1806 14615 1808
rect 18094 1866 18154 2078
rect 18454 1940 18460 2004
rect 18524 2002 18530 2004
rect 18689 2002 18755 2005
rect 18524 2000 18755 2002
rect 18524 1944 18694 2000
rect 18750 1944 18755 2000
rect 18524 1942 18755 1944
rect 18524 1940 18530 1942
rect 18689 1939 18755 1942
rect 20437 1866 20503 1869
rect 22553 1866 22619 1869
rect 18094 1864 22619 1866
rect 18094 1808 20442 1864
rect 20498 1808 22558 1864
rect 22614 1808 22619 1864
rect 18094 1806 22619 1808
rect 12801 1803 12867 1806
rect 14549 1803 14615 1806
rect 20437 1803 20503 1806
rect 22553 1803 22619 1806
rect 12574 1730 12634 1803
rect 15009 1730 15075 1733
rect 12574 1728 15075 1730
rect 12574 1672 15014 1728
rect 15070 1672 15075 1728
rect 12574 1670 15075 1672
rect 15009 1667 15075 1670
rect 19333 1730 19399 1733
rect 19926 1730 19932 1732
rect 19333 1728 19932 1730
rect 19333 1672 19338 1728
rect 19394 1672 19932 1728
rect 19333 1670 19932 1672
rect 19333 1667 19399 1670
rect 19926 1668 19932 1670
rect 19996 1730 20002 1732
rect 20345 1730 20411 1733
rect 19996 1728 20411 1730
rect 19996 1672 20350 1728
rect 20406 1672 20411 1728
rect 19996 1670 20411 1672
rect 19996 1668 20002 1670
rect 20345 1667 20411 1670
rect 4354 1664 4750 1665
rect 4354 1600 4360 1664
rect 4424 1600 4440 1664
rect 4504 1600 4520 1664
rect 4584 1600 4600 1664
rect 4664 1600 4680 1664
rect 4744 1600 4750 1664
rect 4354 1599 4750 1600
rect 10354 1664 10750 1665
rect 10354 1600 10360 1664
rect 10424 1600 10440 1664
rect 10504 1600 10520 1664
rect 10584 1600 10600 1664
rect 10664 1600 10680 1664
rect 10744 1600 10750 1664
rect 10354 1599 10750 1600
rect 16354 1664 16750 1665
rect 16354 1600 16360 1664
rect 16424 1600 16440 1664
rect 16504 1600 16520 1664
rect 16584 1600 16600 1664
rect 16664 1600 16680 1664
rect 16744 1600 16750 1664
rect 16354 1599 16750 1600
rect 22354 1664 22750 1665
rect 22354 1600 22360 1664
rect 22424 1600 22440 1664
rect 22504 1600 22520 1664
rect 22584 1600 22600 1664
rect 22664 1600 22680 1664
rect 22744 1600 22750 1664
rect 22354 1599 22750 1600
rect 5441 1596 5507 1597
rect 5390 1532 5396 1596
rect 5460 1594 5507 1596
rect 12065 1594 12131 1597
rect 15193 1594 15259 1597
rect 15929 1594 15995 1597
rect 5460 1592 5552 1594
rect 5502 1536 5552 1592
rect 5460 1534 5552 1536
rect 12065 1592 15995 1594
rect 12065 1536 12070 1592
rect 12126 1536 15198 1592
rect 15254 1536 15934 1592
rect 15990 1536 15995 1592
rect 12065 1534 15995 1536
rect 5460 1532 5507 1534
rect 5441 1531 5507 1532
rect 12065 1531 12131 1534
rect 15193 1531 15259 1534
rect 15929 1531 15995 1534
rect 6729 1460 6795 1461
rect 6678 1396 6684 1460
rect 6748 1458 6795 1460
rect 8937 1458 9003 1461
rect 10961 1458 11027 1461
rect 13353 1458 13419 1461
rect 19701 1458 19767 1461
rect 20069 1458 20135 1461
rect 6748 1456 6840 1458
rect 6790 1400 6840 1456
rect 6748 1398 6840 1400
rect 8937 1456 10794 1458
rect 8937 1400 8942 1456
rect 8998 1400 10794 1456
rect 8937 1398 10794 1400
rect 6748 1396 6795 1398
rect 6729 1395 6795 1396
rect 8937 1395 9003 1398
rect 9857 1324 9923 1325
rect 9806 1260 9812 1324
rect 9876 1322 9923 1324
rect 10734 1322 10794 1398
rect 10961 1456 13186 1458
rect 10961 1400 10966 1456
rect 11022 1400 13186 1456
rect 10961 1398 13186 1400
rect 10961 1395 11027 1398
rect 11094 1322 11100 1324
rect 9876 1320 9968 1322
rect 9918 1264 9968 1320
rect 9876 1262 9968 1264
rect 10734 1262 11100 1322
rect 9876 1260 9923 1262
rect 11094 1260 11100 1262
rect 11164 1260 11170 1324
rect 13126 1322 13186 1398
rect 13353 1456 20135 1458
rect 13353 1400 13358 1456
rect 13414 1400 19706 1456
rect 19762 1400 20074 1456
rect 20130 1400 20135 1456
rect 13353 1398 20135 1400
rect 13353 1395 13419 1398
rect 19701 1395 19767 1398
rect 20069 1395 20135 1398
rect 19793 1322 19859 1325
rect 20161 1322 20227 1325
rect 20621 1322 20687 1325
rect 13126 1320 20040 1322
rect 13126 1264 19798 1320
rect 19854 1264 20040 1320
rect 13126 1262 20040 1264
rect 9857 1259 9923 1260
rect 19793 1259 19859 1262
rect 14549 1186 14615 1189
rect 16849 1186 16915 1189
rect 14549 1184 16915 1186
rect 14549 1128 14554 1184
rect 14610 1128 16854 1184
rect 16910 1128 16915 1184
rect 14549 1126 16915 1128
rect 19980 1186 20040 1262
rect 20161 1320 20687 1322
rect 20161 1264 20166 1320
rect 20222 1264 20626 1320
rect 20682 1264 20687 1320
rect 20161 1262 20687 1264
rect 20161 1259 20227 1262
rect 20621 1259 20687 1262
rect 20437 1186 20503 1189
rect 19980 1184 20503 1186
rect 19980 1128 20442 1184
rect 20498 1128 20503 1184
rect 19980 1126 20503 1128
rect 14549 1123 14615 1126
rect 16849 1123 16915 1126
rect 20437 1123 20503 1126
rect 1354 1120 1750 1121
rect 1354 1056 1360 1120
rect 1424 1056 1440 1120
rect 1504 1056 1520 1120
rect 1584 1056 1600 1120
rect 1664 1056 1680 1120
rect 1744 1056 1750 1120
rect 1354 1055 1750 1056
rect 7354 1120 7750 1121
rect 7354 1056 7360 1120
rect 7424 1056 7440 1120
rect 7504 1056 7520 1120
rect 7584 1056 7600 1120
rect 7664 1056 7680 1120
rect 7744 1056 7750 1120
rect 7354 1055 7750 1056
rect 13354 1120 13750 1121
rect 13354 1056 13360 1120
rect 13424 1056 13440 1120
rect 13504 1056 13520 1120
rect 13584 1056 13600 1120
rect 13664 1056 13680 1120
rect 13744 1056 13750 1120
rect 13354 1055 13750 1056
rect 19354 1120 19750 1121
rect 19354 1056 19360 1120
rect 19424 1056 19440 1120
rect 19504 1056 19520 1120
rect 19584 1056 19600 1120
rect 19664 1056 19680 1120
rect 19744 1056 19750 1120
rect 19354 1055 19750 1056
rect 14181 1050 14247 1053
rect 14406 1050 14412 1052
rect 14181 1048 14412 1050
rect 14181 992 14186 1048
rect 14242 992 14412 1048
rect 14181 990 14412 992
rect 14181 987 14247 990
rect 14406 988 14412 990
rect 14476 1050 14482 1052
rect 17861 1050 17927 1053
rect 14476 1048 17927 1050
rect 14476 992 17866 1048
rect 17922 992 17927 1048
rect 14476 990 17927 992
rect 14476 988 14482 990
rect 17861 987 17927 990
rect 19885 1050 19951 1053
rect 20713 1050 20779 1053
rect 19885 1048 20779 1050
rect 19885 992 19890 1048
rect 19946 992 20718 1048
rect 20774 992 20779 1048
rect 19885 990 20779 992
rect 19885 987 19951 990
rect 20713 987 20779 990
rect 7097 914 7163 917
rect 21633 914 21699 917
rect 7097 912 21699 914
rect 7097 856 7102 912
rect 7158 856 21638 912
rect 21694 856 21699 912
rect 7097 854 21699 856
rect 7097 851 7163 854
rect 21633 851 21699 854
rect 4521 778 4587 781
rect 5257 778 5323 781
rect 18597 778 18663 781
rect 4521 776 18663 778
rect 4521 720 4526 776
rect 4582 720 5262 776
rect 5318 720 18602 776
rect 18658 720 18663 776
rect 4521 718 18663 720
rect 4521 715 4587 718
rect 5257 715 5323 718
rect 18597 715 18663 718
rect 4354 576 4750 577
rect 4354 512 4360 576
rect 4424 512 4440 576
rect 4504 512 4520 576
rect 4584 512 4600 576
rect 4664 512 4680 576
rect 4744 512 4750 576
rect 4354 511 4750 512
rect 10354 576 10750 577
rect 10354 512 10360 576
rect 10424 512 10440 576
rect 10504 512 10520 576
rect 10584 512 10600 576
rect 10664 512 10680 576
rect 10744 512 10750 576
rect 10354 511 10750 512
rect 16354 576 16750 577
rect 16354 512 16360 576
rect 16424 512 16440 576
rect 16504 512 16520 576
rect 16584 512 16600 576
rect 16664 512 16680 576
rect 16744 512 16750 576
rect 16354 511 16750 512
rect 22354 576 22750 577
rect 22354 512 22360 576
rect 22424 512 22440 576
rect 22504 512 22520 576
rect 22584 512 22600 576
rect 22664 512 22680 576
rect 22744 512 22750 576
rect 22354 511 22750 512
rect 20621 506 20687 509
rect 21817 506 21883 509
rect 20621 504 21883 506
rect 20621 448 20626 504
rect 20682 448 21822 504
rect 21878 448 21883 504
rect 20621 446 21883 448
rect 20621 443 20687 446
rect 21817 443 21883 446
rect 11094 308 11100 372
rect 11164 370 11170 372
rect 19926 370 19932 372
rect 11164 310 19932 370
rect 11164 308 11170 310
rect 19926 308 19932 310
rect 19996 308 20002 372
rect 10041 234 10107 237
rect 17861 234 17927 237
rect 10041 232 17927 234
rect 10041 176 10046 232
rect 10102 176 17866 232
rect 17922 176 17927 232
rect 10041 174 17927 176
rect 10041 171 10107 174
rect 17861 171 17927 174
rect 12065 98 12131 101
rect 17585 98 17651 101
rect 12065 96 17651 98
rect 12065 40 12070 96
rect 12126 40 17590 96
rect 17646 40 17651 96
rect 12065 38 17651 40
rect 12065 35 12131 38
rect 17585 35 17651 38
<< via3 >>
rect 4360 23420 4424 23424
rect 4360 23364 4364 23420
rect 4364 23364 4420 23420
rect 4420 23364 4424 23420
rect 4360 23360 4424 23364
rect 4440 23420 4504 23424
rect 4440 23364 4444 23420
rect 4444 23364 4500 23420
rect 4500 23364 4504 23420
rect 4440 23360 4504 23364
rect 4520 23420 4584 23424
rect 4520 23364 4524 23420
rect 4524 23364 4580 23420
rect 4580 23364 4584 23420
rect 4520 23360 4584 23364
rect 4600 23420 4664 23424
rect 4600 23364 4604 23420
rect 4604 23364 4660 23420
rect 4660 23364 4664 23420
rect 4600 23360 4664 23364
rect 4680 23420 4744 23424
rect 4680 23364 4684 23420
rect 4684 23364 4740 23420
rect 4740 23364 4744 23420
rect 4680 23360 4744 23364
rect 10360 23420 10424 23424
rect 10360 23364 10364 23420
rect 10364 23364 10420 23420
rect 10420 23364 10424 23420
rect 10360 23360 10424 23364
rect 10440 23420 10504 23424
rect 10440 23364 10444 23420
rect 10444 23364 10500 23420
rect 10500 23364 10504 23420
rect 10440 23360 10504 23364
rect 10520 23420 10584 23424
rect 10520 23364 10524 23420
rect 10524 23364 10580 23420
rect 10580 23364 10584 23420
rect 10520 23360 10584 23364
rect 10600 23420 10664 23424
rect 10600 23364 10604 23420
rect 10604 23364 10660 23420
rect 10660 23364 10664 23420
rect 10600 23360 10664 23364
rect 10680 23420 10744 23424
rect 10680 23364 10684 23420
rect 10684 23364 10740 23420
rect 10740 23364 10744 23420
rect 10680 23360 10744 23364
rect 16360 23420 16424 23424
rect 16360 23364 16364 23420
rect 16364 23364 16420 23420
rect 16420 23364 16424 23420
rect 16360 23360 16424 23364
rect 16440 23420 16504 23424
rect 16440 23364 16444 23420
rect 16444 23364 16500 23420
rect 16500 23364 16504 23420
rect 16440 23360 16504 23364
rect 16520 23420 16584 23424
rect 16520 23364 16524 23420
rect 16524 23364 16580 23420
rect 16580 23364 16584 23420
rect 16520 23360 16584 23364
rect 16600 23420 16664 23424
rect 16600 23364 16604 23420
rect 16604 23364 16660 23420
rect 16660 23364 16664 23420
rect 16600 23360 16664 23364
rect 16680 23420 16744 23424
rect 16680 23364 16684 23420
rect 16684 23364 16740 23420
rect 16740 23364 16744 23420
rect 16680 23360 16744 23364
rect 22360 23420 22424 23424
rect 22360 23364 22364 23420
rect 22364 23364 22420 23420
rect 22420 23364 22424 23420
rect 22360 23360 22424 23364
rect 22440 23420 22504 23424
rect 22440 23364 22444 23420
rect 22444 23364 22500 23420
rect 22500 23364 22504 23420
rect 22440 23360 22504 23364
rect 22520 23420 22584 23424
rect 22520 23364 22524 23420
rect 22524 23364 22580 23420
rect 22580 23364 22584 23420
rect 22520 23360 22584 23364
rect 22600 23420 22664 23424
rect 22600 23364 22604 23420
rect 22604 23364 22660 23420
rect 22660 23364 22664 23420
rect 22600 23360 22664 23364
rect 22680 23420 22744 23424
rect 22680 23364 22684 23420
rect 22684 23364 22740 23420
rect 22740 23364 22744 23420
rect 22680 23360 22744 23364
rect 21588 22944 21652 22948
rect 21588 22888 21638 22944
rect 21638 22888 21652 22944
rect 21588 22884 21652 22888
rect 1360 22876 1424 22880
rect 1360 22820 1364 22876
rect 1364 22820 1420 22876
rect 1420 22820 1424 22876
rect 1360 22816 1424 22820
rect 1440 22876 1504 22880
rect 1440 22820 1444 22876
rect 1444 22820 1500 22876
rect 1500 22820 1504 22876
rect 1440 22816 1504 22820
rect 1520 22876 1584 22880
rect 1520 22820 1524 22876
rect 1524 22820 1580 22876
rect 1580 22820 1584 22876
rect 1520 22816 1584 22820
rect 1600 22876 1664 22880
rect 1600 22820 1604 22876
rect 1604 22820 1660 22876
rect 1660 22820 1664 22876
rect 1600 22816 1664 22820
rect 1680 22876 1744 22880
rect 1680 22820 1684 22876
rect 1684 22820 1740 22876
rect 1740 22820 1744 22876
rect 1680 22816 1744 22820
rect 7360 22876 7424 22880
rect 7360 22820 7364 22876
rect 7364 22820 7420 22876
rect 7420 22820 7424 22876
rect 7360 22816 7424 22820
rect 7440 22876 7504 22880
rect 7440 22820 7444 22876
rect 7444 22820 7500 22876
rect 7500 22820 7504 22876
rect 7440 22816 7504 22820
rect 7520 22876 7584 22880
rect 7520 22820 7524 22876
rect 7524 22820 7580 22876
rect 7580 22820 7584 22876
rect 7520 22816 7584 22820
rect 7600 22876 7664 22880
rect 7600 22820 7604 22876
rect 7604 22820 7660 22876
rect 7660 22820 7664 22876
rect 7600 22816 7664 22820
rect 7680 22876 7744 22880
rect 7680 22820 7684 22876
rect 7684 22820 7740 22876
rect 7740 22820 7744 22876
rect 7680 22816 7744 22820
rect 13360 22876 13424 22880
rect 13360 22820 13364 22876
rect 13364 22820 13420 22876
rect 13420 22820 13424 22876
rect 13360 22816 13424 22820
rect 13440 22876 13504 22880
rect 13440 22820 13444 22876
rect 13444 22820 13500 22876
rect 13500 22820 13504 22876
rect 13440 22816 13504 22820
rect 13520 22876 13584 22880
rect 13520 22820 13524 22876
rect 13524 22820 13580 22876
rect 13580 22820 13584 22876
rect 13520 22816 13584 22820
rect 13600 22876 13664 22880
rect 13600 22820 13604 22876
rect 13604 22820 13660 22876
rect 13660 22820 13664 22876
rect 13600 22816 13664 22820
rect 13680 22876 13744 22880
rect 13680 22820 13684 22876
rect 13684 22820 13740 22876
rect 13740 22820 13744 22876
rect 13680 22816 13744 22820
rect 19360 22876 19424 22880
rect 19360 22820 19364 22876
rect 19364 22820 19420 22876
rect 19420 22820 19424 22876
rect 19360 22816 19424 22820
rect 19440 22876 19504 22880
rect 19440 22820 19444 22876
rect 19444 22820 19500 22876
rect 19500 22820 19504 22876
rect 19440 22816 19504 22820
rect 19520 22876 19584 22880
rect 19520 22820 19524 22876
rect 19524 22820 19580 22876
rect 19580 22820 19584 22876
rect 19520 22816 19584 22820
rect 19600 22876 19664 22880
rect 19600 22820 19604 22876
rect 19604 22820 19660 22876
rect 19660 22820 19664 22876
rect 19600 22816 19664 22820
rect 19680 22876 19744 22880
rect 19680 22820 19684 22876
rect 19684 22820 19740 22876
rect 19740 22820 19744 22876
rect 19680 22816 19744 22820
rect 11652 22612 11716 22676
rect 9996 22536 10060 22540
rect 9996 22480 10046 22536
rect 10046 22480 10060 22536
rect 9996 22476 10060 22480
rect 3188 22340 3252 22404
rect 6500 22340 6564 22404
rect 4360 22332 4424 22336
rect 4360 22276 4364 22332
rect 4364 22276 4420 22332
rect 4420 22276 4424 22332
rect 4360 22272 4424 22276
rect 4440 22332 4504 22336
rect 4440 22276 4444 22332
rect 4444 22276 4500 22332
rect 4500 22276 4504 22332
rect 4440 22272 4504 22276
rect 4520 22332 4584 22336
rect 4520 22276 4524 22332
rect 4524 22276 4580 22332
rect 4580 22276 4584 22332
rect 4520 22272 4584 22276
rect 4600 22332 4664 22336
rect 4600 22276 4604 22332
rect 4604 22276 4660 22332
rect 4660 22276 4664 22332
rect 4600 22272 4664 22276
rect 4680 22332 4744 22336
rect 4680 22276 4684 22332
rect 4684 22276 4740 22332
rect 4740 22276 4744 22332
rect 4680 22272 4744 22276
rect 10360 22332 10424 22336
rect 10360 22276 10364 22332
rect 10364 22276 10420 22332
rect 10420 22276 10424 22332
rect 10360 22272 10424 22276
rect 10440 22332 10504 22336
rect 10440 22276 10444 22332
rect 10444 22276 10500 22332
rect 10500 22276 10504 22332
rect 10440 22272 10504 22276
rect 10520 22332 10584 22336
rect 10520 22276 10524 22332
rect 10524 22276 10580 22332
rect 10580 22276 10584 22332
rect 10520 22272 10584 22276
rect 10600 22332 10664 22336
rect 10600 22276 10604 22332
rect 10604 22276 10660 22332
rect 10660 22276 10664 22332
rect 10600 22272 10664 22276
rect 10680 22332 10744 22336
rect 10680 22276 10684 22332
rect 10684 22276 10740 22332
rect 10740 22276 10744 22332
rect 10680 22272 10744 22276
rect 16360 22332 16424 22336
rect 16360 22276 16364 22332
rect 16364 22276 16420 22332
rect 16420 22276 16424 22332
rect 16360 22272 16424 22276
rect 16440 22332 16504 22336
rect 16440 22276 16444 22332
rect 16444 22276 16500 22332
rect 16500 22276 16504 22332
rect 16440 22272 16504 22276
rect 16520 22332 16584 22336
rect 16520 22276 16524 22332
rect 16524 22276 16580 22332
rect 16580 22276 16584 22332
rect 16520 22272 16584 22276
rect 16600 22332 16664 22336
rect 16600 22276 16604 22332
rect 16604 22276 16660 22332
rect 16660 22276 16664 22332
rect 16600 22272 16664 22276
rect 16680 22332 16744 22336
rect 16680 22276 16684 22332
rect 16684 22276 16740 22332
rect 16740 22276 16744 22332
rect 16680 22272 16744 22276
rect 22360 22332 22424 22336
rect 22360 22276 22364 22332
rect 22364 22276 22420 22332
rect 22420 22276 22424 22332
rect 22360 22272 22424 22276
rect 22440 22332 22504 22336
rect 22440 22276 22444 22332
rect 22444 22276 22500 22332
rect 22500 22276 22504 22332
rect 22440 22272 22504 22276
rect 22520 22332 22584 22336
rect 22520 22276 22524 22332
rect 22524 22276 22580 22332
rect 22580 22276 22584 22332
rect 22520 22272 22584 22276
rect 22600 22332 22664 22336
rect 22600 22276 22604 22332
rect 22604 22276 22660 22332
rect 22660 22276 22664 22332
rect 22600 22272 22664 22276
rect 22680 22332 22744 22336
rect 22680 22276 22684 22332
rect 22684 22276 22740 22332
rect 22740 22276 22744 22332
rect 22680 22272 22744 22276
rect 21220 22204 21284 22268
rect 3924 22068 3988 22132
rect 9812 21796 9876 21860
rect 14412 21796 14476 21860
rect 1360 21788 1424 21792
rect 1360 21732 1364 21788
rect 1364 21732 1420 21788
rect 1420 21732 1424 21788
rect 1360 21728 1424 21732
rect 1440 21788 1504 21792
rect 1440 21732 1444 21788
rect 1444 21732 1500 21788
rect 1500 21732 1504 21788
rect 1440 21728 1504 21732
rect 1520 21788 1584 21792
rect 1520 21732 1524 21788
rect 1524 21732 1580 21788
rect 1580 21732 1584 21788
rect 1520 21728 1584 21732
rect 1600 21788 1664 21792
rect 1600 21732 1604 21788
rect 1604 21732 1660 21788
rect 1660 21732 1664 21788
rect 1600 21728 1664 21732
rect 1680 21788 1744 21792
rect 1680 21732 1684 21788
rect 1684 21732 1740 21788
rect 1740 21732 1744 21788
rect 1680 21728 1744 21732
rect 7360 21788 7424 21792
rect 7360 21732 7364 21788
rect 7364 21732 7420 21788
rect 7420 21732 7424 21788
rect 7360 21728 7424 21732
rect 7440 21788 7504 21792
rect 7440 21732 7444 21788
rect 7444 21732 7500 21788
rect 7500 21732 7504 21788
rect 7440 21728 7504 21732
rect 7520 21788 7584 21792
rect 7520 21732 7524 21788
rect 7524 21732 7580 21788
rect 7580 21732 7584 21788
rect 7520 21728 7584 21732
rect 7600 21788 7664 21792
rect 7600 21732 7604 21788
rect 7604 21732 7660 21788
rect 7660 21732 7664 21788
rect 7600 21728 7664 21732
rect 7680 21788 7744 21792
rect 7680 21732 7684 21788
rect 7684 21732 7740 21788
rect 7740 21732 7744 21788
rect 7680 21728 7744 21732
rect 13360 21788 13424 21792
rect 13360 21732 13364 21788
rect 13364 21732 13420 21788
rect 13420 21732 13424 21788
rect 13360 21728 13424 21732
rect 13440 21788 13504 21792
rect 13440 21732 13444 21788
rect 13444 21732 13500 21788
rect 13500 21732 13504 21788
rect 13440 21728 13504 21732
rect 13520 21788 13584 21792
rect 13520 21732 13524 21788
rect 13524 21732 13580 21788
rect 13580 21732 13584 21788
rect 13520 21728 13584 21732
rect 13600 21788 13664 21792
rect 13600 21732 13604 21788
rect 13604 21732 13660 21788
rect 13660 21732 13664 21788
rect 13600 21728 13664 21732
rect 13680 21788 13744 21792
rect 13680 21732 13684 21788
rect 13684 21732 13740 21788
rect 13740 21732 13744 21788
rect 13680 21728 13744 21732
rect 19360 21788 19424 21792
rect 19360 21732 19364 21788
rect 19364 21732 19420 21788
rect 19420 21732 19424 21788
rect 19360 21728 19424 21732
rect 19440 21788 19504 21792
rect 19440 21732 19444 21788
rect 19444 21732 19500 21788
rect 19500 21732 19504 21788
rect 19440 21728 19504 21732
rect 19520 21788 19584 21792
rect 19520 21732 19524 21788
rect 19524 21732 19580 21788
rect 19580 21732 19584 21788
rect 19520 21728 19584 21732
rect 19600 21788 19664 21792
rect 19600 21732 19604 21788
rect 19604 21732 19660 21788
rect 19660 21732 19664 21788
rect 19600 21728 19664 21732
rect 19680 21788 19744 21792
rect 19680 21732 19684 21788
rect 19684 21732 19740 21788
rect 19740 21732 19744 21788
rect 19680 21728 19744 21732
rect 4360 21244 4424 21248
rect 4360 21188 4364 21244
rect 4364 21188 4420 21244
rect 4420 21188 4424 21244
rect 4360 21184 4424 21188
rect 4440 21244 4504 21248
rect 4440 21188 4444 21244
rect 4444 21188 4500 21244
rect 4500 21188 4504 21244
rect 4440 21184 4504 21188
rect 4520 21244 4584 21248
rect 4520 21188 4524 21244
rect 4524 21188 4580 21244
rect 4580 21188 4584 21244
rect 4520 21184 4584 21188
rect 4600 21244 4664 21248
rect 4600 21188 4604 21244
rect 4604 21188 4660 21244
rect 4660 21188 4664 21244
rect 4600 21184 4664 21188
rect 4680 21244 4744 21248
rect 4680 21188 4684 21244
rect 4684 21188 4740 21244
rect 4740 21188 4744 21244
rect 4680 21184 4744 21188
rect 10360 21244 10424 21248
rect 10360 21188 10364 21244
rect 10364 21188 10420 21244
rect 10420 21188 10424 21244
rect 10360 21184 10424 21188
rect 10440 21244 10504 21248
rect 10440 21188 10444 21244
rect 10444 21188 10500 21244
rect 10500 21188 10504 21244
rect 10440 21184 10504 21188
rect 10520 21244 10584 21248
rect 10520 21188 10524 21244
rect 10524 21188 10580 21244
rect 10580 21188 10584 21244
rect 10520 21184 10584 21188
rect 10600 21244 10664 21248
rect 10600 21188 10604 21244
rect 10604 21188 10660 21244
rect 10660 21188 10664 21244
rect 10600 21184 10664 21188
rect 10680 21244 10744 21248
rect 10680 21188 10684 21244
rect 10684 21188 10740 21244
rect 10740 21188 10744 21244
rect 10680 21184 10744 21188
rect 16360 21244 16424 21248
rect 16360 21188 16364 21244
rect 16364 21188 16420 21244
rect 16420 21188 16424 21244
rect 16360 21184 16424 21188
rect 16440 21244 16504 21248
rect 16440 21188 16444 21244
rect 16444 21188 16500 21244
rect 16500 21188 16504 21244
rect 16440 21184 16504 21188
rect 16520 21244 16584 21248
rect 16520 21188 16524 21244
rect 16524 21188 16580 21244
rect 16580 21188 16584 21244
rect 16520 21184 16584 21188
rect 16600 21244 16664 21248
rect 16600 21188 16604 21244
rect 16604 21188 16660 21244
rect 16660 21188 16664 21244
rect 16600 21184 16664 21188
rect 16680 21244 16744 21248
rect 16680 21188 16684 21244
rect 16684 21188 16740 21244
rect 16740 21188 16744 21244
rect 16680 21184 16744 21188
rect 22360 21244 22424 21248
rect 22360 21188 22364 21244
rect 22364 21188 22420 21244
rect 22420 21188 22424 21244
rect 22360 21184 22424 21188
rect 22440 21244 22504 21248
rect 22440 21188 22444 21244
rect 22444 21188 22500 21244
rect 22500 21188 22504 21244
rect 22440 21184 22504 21188
rect 22520 21244 22584 21248
rect 22520 21188 22524 21244
rect 22524 21188 22580 21244
rect 22580 21188 22584 21244
rect 22520 21184 22584 21188
rect 22600 21244 22664 21248
rect 22600 21188 22604 21244
rect 22604 21188 22660 21244
rect 22660 21188 22664 21244
rect 22600 21184 22664 21188
rect 22680 21244 22744 21248
rect 22680 21188 22684 21244
rect 22684 21188 22740 21244
rect 22740 21188 22744 21244
rect 22680 21184 22744 21188
rect 6684 20708 6748 20772
rect 12756 20768 12820 20772
rect 12756 20712 12806 20768
rect 12806 20712 12820 20768
rect 12756 20708 12820 20712
rect 1360 20700 1424 20704
rect 1360 20644 1364 20700
rect 1364 20644 1420 20700
rect 1420 20644 1424 20700
rect 1360 20640 1424 20644
rect 1440 20700 1504 20704
rect 1440 20644 1444 20700
rect 1444 20644 1500 20700
rect 1500 20644 1504 20700
rect 1440 20640 1504 20644
rect 1520 20700 1584 20704
rect 1520 20644 1524 20700
rect 1524 20644 1580 20700
rect 1580 20644 1584 20700
rect 1520 20640 1584 20644
rect 1600 20700 1664 20704
rect 1600 20644 1604 20700
rect 1604 20644 1660 20700
rect 1660 20644 1664 20700
rect 1600 20640 1664 20644
rect 1680 20700 1744 20704
rect 1680 20644 1684 20700
rect 1684 20644 1740 20700
rect 1740 20644 1744 20700
rect 1680 20640 1744 20644
rect 7360 20700 7424 20704
rect 7360 20644 7364 20700
rect 7364 20644 7420 20700
rect 7420 20644 7424 20700
rect 7360 20640 7424 20644
rect 7440 20700 7504 20704
rect 7440 20644 7444 20700
rect 7444 20644 7500 20700
rect 7500 20644 7504 20700
rect 7440 20640 7504 20644
rect 7520 20700 7584 20704
rect 7520 20644 7524 20700
rect 7524 20644 7580 20700
rect 7580 20644 7584 20700
rect 7520 20640 7584 20644
rect 7600 20700 7664 20704
rect 7600 20644 7604 20700
rect 7604 20644 7660 20700
rect 7660 20644 7664 20700
rect 7600 20640 7664 20644
rect 7680 20700 7744 20704
rect 7680 20644 7684 20700
rect 7684 20644 7740 20700
rect 7740 20644 7744 20700
rect 7680 20640 7744 20644
rect 13360 20700 13424 20704
rect 13360 20644 13364 20700
rect 13364 20644 13420 20700
rect 13420 20644 13424 20700
rect 13360 20640 13424 20644
rect 13440 20700 13504 20704
rect 13440 20644 13444 20700
rect 13444 20644 13500 20700
rect 13500 20644 13504 20700
rect 13440 20640 13504 20644
rect 13520 20700 13584 20704
rect 13520 20644 13524 20700
rect 13524 20644 13580 20700
rect 13580 20644 13584 20700
rect 13520 20640 13584 20644
rect 13600 20700 13664 20704
rect 13600 20644 13604 20700
rect 13604 20644 13660 20700
rect 13660 20644 13664 20700
rect 13600 20640 13664 20644
rect 13680 20700 13744 20704
rect 13680 20644 13684 20700
rect 13684 20644 13740 20700
rect 13740 20644 13744 20700
rect 13680 20640 13744 20644
rect 21036 20844 21100 20908
rect 19360 20700 19424 20704
rect 19360 20644 19364 20700
rect 19364 20644 19420 20700
rect 19420 20644 19424 20700
rect 19360 20640 19424 20644
rect 19440 20700 19504 20704
rect 19440 20644 19444 20700
rect 19444 20644 19500 20700
rect 19500 20644 19504 20700
rect 19440 20640 19504 20644
rect 19520 20700 19584 20704
rect 19520 20644 19524 20700
rect 19524 20644 19580 20700
rect 19580 20644 19584 20700
rect 19520 20640 19584 20644
rect 19600 20700 19664 20704
rect 19600 20644 19604 20700
rect 19604 20644 19660 20700
rect 19660 20644 19664 20700
rect 19600 20640 19664 20644
rect 19680 20700 19744 20704
rect 19680 20644 19684 20700
rect 19684 20644 19740 20700
rect 19740 20644 19744 20700
rect 19680 20640 19744 20644
rect 4360 20156 4424 20160
rect 4360 20100 4364 20156
rect 4364 20100 4420 20156
rect 4420 20100 4424 20156
rect 4360 20096 4424 20100
rect 4440 20156 4504 20160
rect 4440 20100 4444 20156
rect 4444 20100 4500 20156
rect 4500 20100 4504 20156
rect 4440 20096 4504 20100
rect 4520 20156 4584 20160
rect 4520 20100 4524 20156
rect 4524 20100 4580 20156
rect 4580 20100 4584 20156
rect 4520 20096 4584 20100
rect 4600 20156 4664 20160
rect 4600 20100 4604 20156
rect 4604 20100 4660 20156
rect 4660 20100 4664 20156
rect 4600 20096 4664 20100
rect 4680 20156 4744 20160
rect 4680 20100 4684 20156
rect 4684 20100 4740 20156
rect 4740 20100 4744 20156
rect 4680 20096 4744 20100
rect 10360 20156 10424 20160
rect 10360 20100 10364 20156
rect 10364 20100 10420 20156
rect 10420 20100 10424 20156
rect 10360 20096 10424 20100
rect 10440 20156 10504 20160
rect 10440 20100 10444 20156
rect 10444 20100 10500 20156
rect 10500 20100 10504 20156
rect 10440 20096 10504 20100
rect 10520 20156 10584 20160
rect 10520 20100 10524 20156
rect 10524 20100 10580 20156
rect 10580 20100 10584 20156
rect 10520 20096 10584 20100
rect 10600 20156 10664 20160
rect 10600 20100 10604 20156
rect 10604 20100 10660 20156
rect 10660 20100 10664 20156
rect 10600 20096 10664 20100
rect 10680 20156 10744 20160
rect 10680 20100 10684 20156
rect 10684 20100 10740 20156
rect 10740 20100 10744 20156
rect 10680 20096 10744 20100
rect 16360 20156 16424 20160
rect 16360 20100 16364 20156
rect 16364 20100 16420 20156
rect 16420 20100 16424 20156
rect 16360 20096 16424 20100
rect 16440 20156 16504 20160
rect 16440 20100 16444 20156
rect 16444 20100 16500 20156
rect 16500 20100 16504 20156
rect 16440 20096 16504 20100
rect 16520 20156 16584 20160
rect 16520 20100 16524 20156
rect 16524 20100 16580 20156
rect 16580 20100 16584 20156
rect 16520 20096 16584 20100
rect 16600 20156 16664 20160
rect 16600 20100 16604 20156
rect 16604 20100 16660 20156
rect 16660 20100 16664 20156
rect 16600 20096 16664 20100
rect 16680 20156 16744 20160
rect 16680 20100 16684 20156
rect 16684 20100 16740 20156
rect 16740 20100 16744 20156
rect 16680 20096 16744 20100
rect 22360 20156 22424 20160
rect 22360 20100 22364 20156
rect 22364 20100 22420 20156
rect 22420 20100 22424 20156
rect 22360 20096 22424 20100
rect 22440 20156 22504 20160
rect 22440 20100 22444 20156
rect 22444 20100 22500 20156
rect 22500 20100 22504 20156
rect 22440 20096 22504 20100
rect 22520 20156 22584 20160
rect 22520 20100 22524 20156
rect 22524 20100 22580 20156
rect 22580 20100 22584 20156
rect 22520 20096 22584 20100
rect 22600 20156 22664 20160
rect 22600 20100 22604 20156
rect 22604 20100 22660 20156
rect 22660 20100 22664 20156
rect 22600 20096 22664 20100
rect 22680 20156 22744 20160
rect 22680 20100 22684 20156
rect 22684 20100 22740 20156
rect 22740 20100 22744 20156
rect 22680 20096 22744 20100
rect 1360 19612 1424 19616
rect 1360 19556 1364 19612
rect 1364 19556 1420 19612
rect 1420 19556 1424 19612
rect 1360 19552 1424 19556
rect 1440 19612 1504 19616
rect 1440 19556 1444 19612
rect 1444 19556 1500 19612
rect 1500 19556 1504 19612
rect 1440 19552 1504 19556
rect 1520 19612 1584 19616
rect 1520 19556 1524 19612
rect 1524 19556 1580 19612
rect 1580 19556 1584 19612
rect 1520 19552 1584 19556
rect 1600 19612 1664 19616
rect 1600 19556 1604 19612
rect 1604 19556 1660 19612
rect 1660 19556 1664 19612
rect 1600 19552 1664 19556
rect 1680 19612 1744 19616
rect 1680 19556 1684 19612
rect 1684 19556 1740 19612
rect 1740 19556 1744 19612
rect 1680 19552 1744 19556
rect 7360 19612 7424 19616
rect 7360 19556 7364 19612
rect 7364 19556 7420 19612
rect 7420 19556 7424 19612
rect 7360 19552 7424 19556
rect 7440 19612 7504 19616
rect 7440 19556 7444 19612
rect 7444 19556 7500 19612
rect 7500 19556 7504 19612
rect 7440 19552 7504 19556
rect 7520 19612 7584 19616
rect 7520 19556 7524 19612
rect 7524 19556 7580 19612
rect 7580 19556 7584 19612
rect 7520 19552 7584 19556
rect 7600 19612 7664 19616
rect 7600 19556 7604 19612
rect 7604 19556 7660 19612
rect 7660 19556 7664 19612
rect 7600 19552 7664 19556
rect 7680 19612 7744 19616
rect 7680 19556 7684 19612
rect 7684 19556 7740 19612
rect 7740 19556 7744 19612
rect 7680 19552 7744 19556
rect 18828 19620 18892 19684
rect 13360 19612 13424 19616
rect 13360 19556 13364 19612
rect 13364 19556 13420 19612
rect 13420 19556 13424 19612
rect 13360 19552 13424 19556
rect 13440 19612 13504 19616
rect 13440 19556 13444 19612
rect 13444 19556 13500 19612
rect 13500 19556 13504 19612
rect 13440 19552 13504 19556
rect 13520 19612 13584 19616
rect 13520 19556 13524 19612
rect 13524 19556 13580 19612
rect 13580 19556 13584 19612
rect 13520 19552 13584 19556
rect 13600 19612 13664 19616
rect 13600 19556 13604 19612
rect 13604 19556 13660 19612
rect 13660 19556 13664 19612
rect 13600 19552 13664 19556
rect 13680 19612 13744 19616
rect 13680 19556 13684 19612
rect 13684 19556 13740 19612
rect 13740 19556 13744 19612
rect 13680 19552 13744 19556
rect 19360 19612 19424 19616
rect 19360 19556 19364 19612
rect 19364 19556 19420 19612
rect 19420 19556 19424 19612
rect 19360 19552 19424 19556
rect 19440 19612 19504 19616
rect 19440 19556 19444 19612
rect 19444 19556 19500 19612
rect 19500 19556 19504 19612
rect 19440 19552 19504 19556
rect 19520 19612 19584 19616
rect 19520 19556 19524 19612
rect 19524 19556 19580 19612
rect 19580 19556 19584 19612
rect 19520 19552 19584 19556
rect 19600 19612 19664 19616
rect 19600 19556 19604 19612
rect 19604 19556 19660 19612
rect 19660 19556 19664 19612
rect 19600 19552 19664 19556
rect 19680 19612 19744 19616
rect 19680 19556 19684 19612
rect 19684 19556 19740 19612
rect 19740 19556 19744 19612
rect 19680 19552 19744 19556
rect 19012 19408 19076 19412
rect 19012 19352 19026 19408
rect 19026 19352 19076 19408
rect 19012 19348 19076 19352
rect 15700 19212 15764 19276
rect 21220 19212 21284 19276
rect 10180 19076 10244 19140
rect 4360 19068 4424 19072
rect 4360 19012 4364 19068
rect 4364 19012 4420 19068
rect 4420 19012 4424 19068
rect 4360 19008 4424 19012
rect 4440 19068 4504 19072
rect 4440 19012 4444 19068
rect 4444 19012 4500 19068
rect 4500 19012 4504 19068
rect 4440 19008 4504 19012
rect 4520 19068 4584 19072
rect 4520 19012 4524 19068
rect 4524 19012 4580 19068
rect 4580 19012 4584 19068
rect 4520 19008 4584 19012
rect 4600 19068 4664 19072
rect 4600 19012 4604 19068
rect 4604 19012 4660 19068
rect 4660 19012 4664 19068
rect 4600 19008 4664 19012
rect 4680 19068 4744 19072
rect 4680 19012 4684 19068
rect 4684 19012 4740 19068
rect 4740 19012 4744 19068
rect 4680 19008 4744 19012
rect 10360 19068 10424 19072
rect 10360 19012 10364 19068
rect 10364 19012 10420 19068
rect 10420 19012 10424 19068
rect 10360 19008 10424 19012
rect 10440 19068 10504 19072
rect 10440 19012 10444 19068
rect 10444 19012 10500 19068
rect 10500 19012 10504 19068
rect 10440 19008 10504 19012
rect 10520 19068 10584 19072
rect 10520 19012 10524 19068
rect 10524 19012 10580 19068
rect 10580 19012 10584 19068
rect 10520 19008 10584 19012
rect 10600 19068 10664 19072
rect 10600 19012 10604 19068
rect 10604 19012 10660 19068
rect 10660 19012 10664 19068
rect 10600 19008 10664 19012
rect 10680 19068 10744 19072
rect 10680 19012 10684 19068
rect 10684 19012 10740 19068
rect 10740 19012 10744 19068
rect 10680 19008 10744 19012
rect 16360 19068 16424 19072
rect 16360 19012 16364 19068
rect 16364 19012 16420 19068
rect 16420 19012 16424 19068
rect 16360 19008 16424 19012
rect 16440 19068 16504 19072
rect 16440 19012 16444 19068
rect 16444 19012 16500 19068
rect 16500 19012 16504 19068
rect 16440 19008 16504 19012
rect 16520 19068 16584 19072
rect 16520 19012 16524 19068
rect 16524 19012 16580 19068
rect 16580 19012 16584 19068
rect 16520 19008 16584 19012
rect 16600 19068 16664 19072
rect 16600 19012 16604 19068
rect 16604 19012 16660 19068
rect 16660 19012 16664 19068
rect 16600 19008 16664 19012
rect 16680 19068 16744 19072
rect 16680 19012 16684 19068
rect 16684 19012 16740 19068
rect 16740 19012 16744 19068
rect 16680 19008 16744 19012
rect 22360 19068 22424 19072
rect 22360 19012 22364 19068
rect 22364 19012 22420 19068
rect 22420 19012 22424 19068
rect 22360 19008 22424 19012
rect 22440 19068 22504 19072
rect 22440 19012 22444 19068
rect 22444 19012 22500 19068
rect 22500 19012 22504 19068
rect 22440 19008 22504 19012
rect 22520 19068 22584 19072
rect 22520 19012 22524 19068
rect 22524 19012 22580 19068
rect 22580 19012 22584 19068
rect 22520 19008 22584 19012
rect 22600 19068 22664 19072
rect 22600 19012 22604 19068
rect 22604 19012 22660 19068
rect 22660 19012 22664 19068
rect 22600 19008 22664 19012
rect 22680 19068 22744 19072
rect 22680 19012 22684 19068
rect 22684 19012 22740 19068
rect 22740 19012 22744 19068
rect 22680 19008 22744 19012
rect 19932 18592 19996 18596
rect 19932 18536 19946 18592
rect 19946 18536 19996 18592
rect 19932 18532 19996 18536
rect 1360 18524 1424 18528
rect 1360 18468 1364 18524
rect 1364 18468 1420 18524
rect 1420 18468 1424 18524
rect 1360 18464 1424 18468
rect 1440 18524 1504 18528
rect 1440 18468 1444 18524
rect 1444 18468 1500 18524
rect 1500 18468 1504 18524
rect 1440 18464 1504 18468
rect 1520 18524 1584 18528
rect 1520 18468 1524 18524
rect 1524 18468 1580 18524
rect 1580 18468 1584 18524
rect 1520 18464 1584 18468
rect 1600 18524 1664 18528
rect 1600 18468 1604 18524
rect 1604 18468 1660 18524
rect 1660 18468 1664 18524
rect 1600 18464 1664 18468
rect 1680 18524 1744 18528
rect 1680 18468 1684 18524
rect 1684 18468 1740 18524
rect 1740 18468 1744 18524
rect 1680 18464 1744 18468
rect 7360 18524 7424 18528
rect 7360 18468 7364 18524
rect 7364 18468 7420 18524
rect 7420 18468 7424 18524
rect 7360 18464 7424 18468
rect 7440 18524 7504 18528
rect 7440 18468 7444 18524
rect 7444 18468 7500 18524
rect 7500 18468 7504 18524
rect 7440 18464 7504 18468
rect 7520 18524 7584 18528
rect 7520 18468 7524 18524
rect 7524 18468 7580 18524
rect 7580 18468 7584 18524
rect 7520 18464 7584 18468
rect 7600 18524 7664 18528
rect 7600 18468 7604 18524
rect 7604 18468 7660 18524
rect 7660 18468 7664 18524
rect 7600 18464 7664 18468
rect 7680 18524 7744 18528
rect 7680 18468 7684 18524
rect 7684 18468 7740 18524
rect 7740 18468 7744 18524
rect 7680 18464 7744 18468
rect 13360 18524 13424 18528
rect 13360 18468 13364 18524
rect 13364 18468 13420 18524
rect 13420 18468 13424 18524
rect 13360 18464 13424 18468
rect 13440 18524 13504 18528
rect 13440 18468 13444 18524
rect 13444 18468 13500 18524
rect 13500 18468 13504 18524
rect 13440 18464 13504 18468
rect 13520 18524 13584 18528
rect 13520 18468 13524 18524
rect 13524 18468 13580 18524
rect 13580 18468 13584 18524
rect 13520 18464 13584 18468
rect 13600 18524 13664 18528
rect 13600 18468 13604 18524
rect 13604 18468 13660 18524
rect 13660 18468 13664 18524
rect 13600 18464 13664 18468
rect 13680 18524 13744 18528
rect 13680 18468 13684 18524
rect 13684 18468 13740 18524
rect 13740 18468 13744 18524
rect 13680 18464 13744 18468
rect 19360 18524 19424 18528
rect 19360 18468 19364 18524
rect 19364 18468 19420 18524
rect 19420 18468 19424 18524
rect 19360 18464 19424 18468
rect 19440 18524 19504 18528
rect 19440 18468 19444 18524
rect 19444 18468 19500 18524
rect 19500 18468 19504 18524
rect 19440 18464 19504 18468
rect 19520 18524 19584 18528
rect 19520 18468 19524 18524
rect 19524 18468 19580 18524
rect 19580 18468 19584 18524
rect 19520 18464 19584 18468
rect 19600 18524 19664 18528
rect 19600 18468 19604 18524
rect 19604 18468 19660 18524
rect 19660 18468 19664 18524
rect 19600 18464 19664 18468
rect 19680 18524 19744 18528
rect 19680 18468 19684 18524
rect 19684 18468 19740 18524
rect 19740 18468 19744 18524
rect 19680 18464 19744 18468
rect 9444 18124 9508 18188
rect 14964 17988 15028 18052
rect 20668 17988 20732 18052
rect 21588 18048 21652 18052
rect 21588 17992 21602 18048
rect 21602 17992 21652 18048
rect 21588 17988 21652 17992
rect 4360 17980 4424 17984
rect 4360 17924 4364 17980
rect 4364 17924 4420 17980
rect 4420 17924 4424 17980
rect 4360 17920 4424 17924
rect 4440 17980 4504 17984
rect 4440 17924 4444 17980
rect 4444 17924 4500 17980
rect 4500 17924 4504 17980
rect 4440 17920 4504 17924
rect 4520 17980 4584 17984
rect 4520 17924 4524 17980
rect 4524 17924 4580 17980
rect 4580 17924 4584 17980
rect 4520 17920 4584 17924
rect 4600 17980 4664 17984
rect 4600 17924 4604 17980
rect 4604 17924 4660 17980
rect 4660 17924 4664 17980
rect 4600 17920 4664 17924
rect 4680 17980 4744 17984
rect 4680 17924 4684 17980
rect 4684 17924 4740 17980
rect 4740 17924 4744 17980
rect 4680 17920 4744 17924
rect 10360 17980 10424 17984
rect 10360 17924 10364 17980
rect 10364 17924 10420 17980
rect 10420 17924 10424 17980
rect 10360 17920 10424 17924
rect 10440 17980 10504 17984
rect 10440 17924 10444 17980
rect 10444 17924 10500 17980
rect 10500 17924 10504 17980
rect 10440 17920 10504 17924
rect 10520 17980 10584 17984
rect 10520 17924 10524 17980
rect 10524 17924 10580 17980
rect 10580 17924 10584 17980
rect 10520 17920 10584 17924
rect 10600 17980 10664 17984
rect 10600 17924 10604 17980
rect 10604 17924 10660 17980
rect 10660 17924 10664 17980
rect 10600 17920 10664 17924
rect 10680 17980 10744 17984
rect 10680 17924 10684 17980
rect 10684 17924 10740 17980
rect 10740 17924 10744 17980
rect 10680 17920 10744 17924
rect 16360 17980 16424 17984
rect 16360 17924 16364 17980
rect 16364 17924 16420 17980
rect 16420 17924 16424 17980
rect 16360 17920 16424 17924
rect 16440 17980 16504 17984
rect 16440 17924 16444 17980
rect 16444 17924 16500 17980
rect 16500 17924 16504 17980
rect 16440 17920 16504 17924
rect 16520 17980 16584 17984
rect 16520 17924 16524 17980
rect 16524 17924 16580 17980
rect 16580 17924 16584 17980
rect 16520 17920 16584 17924
rect 16600 17980 16664 17984
rect 16600 17924 16604 17980
rect 16604 17924 16660 17980
rect 16660 17924 16664 17980
rect 16600 17920 16664 17924
rect 16680 17980 16744 17984
rect 16680 17924 16684 17980
rect 16684 17924 16740 17980
rect 16740 17924 16744 17980
rect 16680 17920 16744 17924
rect 22360 17980 22424 17984
rect 22360 17924 22364 17980
rect 22364 17924 22420 17980
rect 22420 17924 22424 17980
rect 22360 17920 22424 17924
rect 22440 17980 22504 17984
rect 22440 17924 22444 17980
rect 22444 17924 22500 17980
rect 22500 17924 22504 17980
rect 22440 17920 22504 17924
rect 22520 17980 22584 17984
rect 22520 17924 22524 17980
rect 22524 17924 22580 17980
rect 22580 17924 22584 17980
rect 22520 17920 22584 17924
rect 22600 17980 22664 17984
rect 22600 17924 22604 17980
rect 22604 17924 22660 17980
rect 22660 17924 22664 17980
rect 22600 17920 22664 17924
rect 22680 17980 22744 17984
rect 22680 17924 22684 17980
rect 22684 17924 22740 17980
rect 22740 17924 22744 17980
rect 22680 17920 22744 17924
rect 7972 17852 8036 17916
rect 11836 17580 11900 17644
rect 21036 17580 21100 17644
rect 1360 17436 1424 17440
rect 1360 17380 1364 17436
rect 1364 17380 1420 17436
rect 1420 17380 1424 17436
rect 1360 17376 1424 17380
rect 1440 17436 1504 17440
rect 1440 17380 1444 17436
rect 1444 17380 1500 17436
rect 1500 17380 1504 17436
rect 1440 17376 1504 17380
rect 1520 17436 1584 17440
rect 1520 17380 1524 17436
rect 1524 17380 1580 17436
rect 1580 17380 1584 17436
rect 1520 17376 1584 17380
rect 1600 17436 1664 17440
rect 1600 17380 1604 17436
rect 1604 17380 1660 17436
rect 1660 17380 1664 17436
rect 1600 17376 1664 17380
rect 1680 17436 1744 17440
rect 1680 17380 1684 17436
rect 1684 17380 1740 17436
rect 1740 17380 1744 17436
rect 1680 17376 1744 17380
rect 7360 17436 7424 17440
rect 7360 17380 7364 17436
rect 7364 17380 7420 17436
rect 7420 17380 7424 17436
rect 7360 17376 7424 17380
rect 7440 17436 7504 17440
rect 7440 17380 7444 17436
rect 7444 17380 7500 17436
rect 7500 17380 7504 17436
rect 7440 17376 7504 17380
rect 7520 17436 7584 17440
rect 7520 17380 7524 17436
rect 7524 17380 7580 17436
rect 7580 17380 7584 17436
rect 7520 17376 7584 17380
rect 7600 17436 7664 17440
rect 7600 17380 7604 17436
rect 7604 17380 7660 17436
rect 7660 17380 7664 17436
rect 7600 17376 7664 17380
rect 7680 17436 7744 17440
rect 7680 17380 7684 17436
rect 7684 17380 7740 17436
rect 7740 17380 7744 17436
rect 7680 17376 7744 17380
rect 13360 17436 13424 17440
rect 13360 17380 13364 17436
rect 13364 17380 13420 17436
rect 13420 17380 13424 17436
rect 13360 17376 13424 17380
rect 13440 17436 13504 17440
rect 13440 17380 13444 17436
rect 13444 17380 13500 17436
rect 13500 17380 13504 17436
rect 13440 17376 13504 17380
rect 13520 17436 13584 17440
rect 13520 17380 13524 17436
rect 13524 17380 13580 17436
rect 13580 17380 13584 17436
rect 13520 17376 13584 17380
rect 13600 17436 13664 17440
rect 13600 17380 13604 17436
rect 13604 17380 13660 17436
rect 13660 17380 13664 17436
rect 13600 17376 13664 17380
rect 13680 17436 13744 17440
rect 13680 17380 13684 17436
rect 13684 17380 13740 17436
rect 13740 17380 13744 17436
rect 13680 17376 13744 17380
rect 19360 17436 19424 17440
rect 19360 17380 19364 17436
rect 19364 17380 19420 17436
rect 19420 17380 19424 17436
rect 19360 17376 19424 17380
rect 19440 17436 19504 17440
rect 19440 17380 19444 17436
rect 19444 17380 19500 17436
rect 19500 17380 19504 17436
rect 19440 17376 19504 17380
rect 19520 17436 19584 17440
rect 19520 17380 19524 17436
rect 19524 17380 19580 17436
rect 19580 17380 19584 17436
rect 19520 17376 19584 17380
rect 19600 17436 19664 17440
rect 19600 17380 19604 17436
rect 19604 17380 19660 17436
rect 19660 17380 19664 17436
rect 19600 17376 19664 17380
rect 19680 17436 19744 17440
rect 19680 17380 19684 17436
rect 19684 17380 19740 17436
rect 19740 17380 19744 17436
rect 19680 17376 19744 17380
rect 9444 17172 9508 17236
rect 5764 17096 5828 17100
rect 5764 17040 5814 17096
rect 5814 17040 5828 17096
rect 5764 17036 5828 17040
rect 4360 16892 4424 16896
rect 4360 16836 4364 16892
rect 4364 16836 4420 16892
rect 4420 16836 4424 16892
rect 4360 16832 4424 16836
rect 4440 16892 4504 16896
rect 4440 16836 4444 16892
rect 4444 16836 4500 16892
rect 4500 16836 4504 16892
rect 4440 16832 4504 16836
rect 4520 16892 4584 16896
rect 4520 16836 4524 16892
rect 4524 16836 4580 16892
rect 4580 16836 4584 16892
rect 4520 16832 4584 16836
rect 4600 16892 4664 16896
rect 4600 16836 4604 16892
rect 4604 16836 4660 16892
rect 4660 16836 4664 16892
rect 4600 16832 4664 16836
rect 4680 16892 4744 16896
rect 4680 16836 4684 16892
rect 4684 16836 4740 16892
rect 4740 16836 4744 16892
rect 4680 16832 4744 16836
rect 10360 16892 10424 16896
rect 10360 16836 10364 16892
rect 10364 16836 10420 16892
rect 10420 16836 10424 16892
rect 10360 16832 10424 16836
rect 10440 16892 10504 16896
rect 10440 16836 10444 16892
rect 10444 16836 10500 16892
rect 10500 16836 10504 16892
rect 10440 16832 10504 16836
rect 10520 16892 10584 16896
rect 10520 16836 10524 16892
rect 10524 16836 10580 16892
rect 10580 16836 10584 16892
rect 10520 16832 10584 16836
rect 10600 16892 10664 16896
rect 10600 16836 10604 16892
rect 10604 16836 10660 16892
rect 10660 16836 10664 16892
rect 10600 16832 10664 16836
rect 10680 16892 10744 16896
rect 10680 16836 10684 16892
rect 10684 16836 10740 16892
rect 10740 16836 10744 16892
rect 10680 16832 10744 16836
rect 16360 16892 16424 16896
rect 16360 16836 16364 16892
rect 16364 16836 16420 16892
rect 16420 16836 16424 16892
rect 16360 16832 16424 16836
rect 16440 16892 16504 16896
rect 16440 16836 16444 16892
rect 16444 16836 16500 16892
rect 16500 16836 16504 16892
rect 16440 16832 16504 16836
rect 16520 16892 16584 16896
rect 16520 16836 16524 16892
rect 16524 16836 16580 16892
rect 16580 16836 16584 16892
rect 16520 16832 16584 16836
rect 16600 16892 16664 16896
rect 16600 16836 16604 16892
rect 16604 16836 16660 16892
rect 16660 16836 16664 16892
rect 16600 16832 16664 16836
rect 16680 16892 16744 16896
rect 16680 16836 16684 16892
rect 16684 16836 16740 16892
rect 16740 16836 16744 16892
rect 16680 16832 16744 16836
rect 22360 16892 22424 16896
rect 22360 16836 22364 16892
rect 22364 16836 22420 16892
rect 22420 16836 22424 16892
rect 22360 16832 22424 16836
rect 22440 16892 22504 16896
rect 22440 16836 22444 16892
rect 22444 16836 22500 16892
rect 22500 16836 22504 16892
rect 22440 16832 22504 16836
rect 22520 16892 22584 16896
rect 22520 16836 22524 16892
rect 22524 16836 22580 16892
rect 22580 16836 22584 16892
rect 22520 16832 22584 16836
rect 22600 16892 22664 16896
rect 22600 16836 22604 16892
rect 22604 16836 22660 16892
rect 22660 16836 22664 16892
rect 22600 16832 22664 16836
rect 22680 16892 22744 16896
rect 22680 16836 22684 16892
rect 22684 16836 22740 16892
rect 22740 16836 22744 16892
rect 22680 16832 22744 16836
rect 1360 16348 1424 16352
rect 1360 16292 1364 16348
rect 1364 16292 1420 16348
rect 1420 16292 1424 16348
rect 1360 16288 1424 16292
rect 1440 16348 1504 16352
rect 1440 16292 1444 16348
rect 1444 16292 1500 16348
rect 1500 16292 1504 16348
rect 1440 16288 1504 16292
rect 1520 16348 1584 16352
rect 1520 16292 1524 16348
rect 1524 16292 1580 16348
rect 1580 16292 1584 16348
rect 1520 16288 1584 16292
rect 1600 16348 1664 16352
rect 1600 16292 1604 16348
rect 1604 16292 1660 16348
rect 1660 16292 1664 16348
rect 1600 16288 1664 16292
rect 1680 16348 1744 16352
rect 1680 16292 1684 16348
rect 1684 16292 1740 16348
rect 1740 16292 1744 16348
rect 1680 16288 1744 16292
rect 7360 16348 7424 16352
rect 7360 16292 7364 16348
rect 7364 16292 7420 16348
rect 7420 16292 7424 16348
rect 7360 16288 7424 16292
rect 7440 16348 7504 16352
rect 7440 16292 7444 16348
rect 7444 16292 7500 16348
rect 7500 16292 7504 16348
rect 7440 16288 7504 16292
rect 7520 16348 7584 16352
rect 7520 16292 7524 16348
rect 7524 16292 7580 16348
rect 7580 16292 7584 16348
rect 7520 16288 7584 16292
rect 7600 16348 7664 16352
rect 7600 16292 7604 16348
rect 7604 16292 7660 16348
rect 7660 16292 7664 16348
rect 7600 16288 7664 16292
rect 7680 16348 7744 16352
rect 7680 16292 7684 16348
rect 7684 16292 7740 16348
rect 7740 16292 7744 16348
rect 7680 16288 7744 16292
rect 13360 16348 13424 16352
rect 13360 16292 13364 16348
rect 13364 16292 13420 16348
rect 13420 16292 13424 16348
rect 13360 16288 13424 16292
rect 13440 16348 13504 16352
rect 13440 16292 13444 16348
rect 13444 16292 13500 16348
rect 13500 16292 13504 16348
rect 13440 16288 13504 16292
rect 13520 16348 13584 16352
rect 13520 16292 13524 16348
rect 13524 16292 13580 16348
rect 13580 16292 13584 16348
rect 13520 16288 13584 16292
rect 13600 16348 13664 16352
rect 13600 16292 13604 16348
rect 13604 16292 13660 16348
rect 13660 16292 13664 16348
rect 13600 16288 13664 16292
rect 13680 16348 13744 16352
rect 13680 16292 13684 16348
rect 13684 16292 13740 16348
rect 13740 16292 13744 16348
rect 13680 16288 13744 16292
rect 19360 16348 19424 16352
rect 19360 16292 19364 16348
rect 19364 16292 19420 16348
rect 19420 16292 19424 16348
rect 19360 16288 19424 16292
rect 19440 16348 19504 16352
rect 19440 16292 19444 16348
rect 19444 16292 19500 16348
rect 19500 16292 19504 16348
rect 19440 16288 19504 16292
rect 19520 16348 19584 16352
rect 19520 16292 19524 16348
rect 19524 16292 19580 16348
rect 19580 16292 19584 16348
rect 19520 16288 19584 16292
rect 19600 16348 19664 16352
rect 19600 16292 19604 16348
rect 19604 16292 19660 16348
rect 19660 16292 19664 16348
rect 19600 16288 19664 16292
rect 19680 16348 19744 16352
rect 19680 16292 19684 16348
rect 19684 16292 19740 16348
rect 19740 16292 19744 16348
rect 19680 16288 19744 16292
rect 4360 15804 4424 15808
rect 4360 15748 4364 15804
rect 4364 15748 4420 15804
rect 4420 15748 4424 15804
rect 4360 15744 4424 15748
rect 4440 15804 4504 15808
rect 4440 15748 4444 15804
rect 4444 15748 4500 15804
rect 4500 15748 4504 15804
rect 4440 15744 4504 15748
rect 4520 15804 4584 15808
rect 4520 15748 4524 15804
rect 4524 15748 4580 15804
rect 4580 15748 4584 15804
rect 4520 15744 4584 15748
rect 4600 15804 4664 15808
rect 4600 15748 4604 15804
rect 4604 15748 4660 15804
rect 4660 15748 4664 15804
rect 4600 15744 4664 15748
rect 4680 15804 4744 15808
rect 4680 15748 4684 15804
rect 4684 15748 4740 15804
rect 4740 15748 4744 15804
rect 4680 15744 4744 15748
rect 10360 15804 10424 15808
rect 10360 15748 10364 15804
rect 10364 15748 10420 15804
rect 10420 15748 10424 15804
rect 10360 15744 10424 15748
rect 10440 15804 10504 15808
rect 10440 15748 10444 15804
rect 10444 15748 10500 15804
rect 10500 15748 10504 15804
rect 10440 15744 10504 15748
rect 10520 15804 10584 15808
rect 10520 15748 10524 15804
rect 10524 15748 10580 15804
rect 10580 15748 10584 15804
rect 10520 15744 10584 15748
rect 10600 15804 10664 15808
rect 10600 15748 10604 15804
rect 10604 15748 10660 15804
rect 10660 15748 10664 15804
rect 10600 15744 10664 15748
rect 10680 15804 10744 15808
rect 10680 15748 10684 15804
rect 10684 15748 10740 15804
rect 10740 15748 10744 15804
rect 10680 15744 10744 15748
rect 16360 15804 16424 15808
rect 16360 15748 16364 15804
rect 16364 15748 16420 15804
rect 16420 15748 16424 15804
rect 16360 15744 16424 15748
rect 16440 15804 16504 15808
rect 16440 15748 16444 15804
rect 16444 15748 16500 15804
rect 16500 15748 16504 15804
rect 16440 15744 16504 15748
rect 16520 15804 16584 15808
rect 16520 15748 16524 15804
rect 16524 15748 16580 15804
rect 16580 15748 16584 15804
rect 16520 15744 16584 15748
rect 16600 15804 16664 15808
rect 16600 15748 16604 15804
rect 16604 15748 16660 15804
rect 16660 15748 16664 15804
rect 16600 15744 16664 15748
rect 16680 15804 16744 15808
rect 16680 15748 16684 15804
rect 16684 15748 16740 15804
rect 16740 15748 16744 15804
rect 16680 15744 16744 15748
rect 22360 15804 22424 15808
rect 22360 15748 22364 15804
rect 22364 15748 22420 15804
rect 22420 15748 22424 15804
rect 22360 15744 22424 15748
rect 22440 15804 22504 15808
rect 22440 15748 22444 15804
rect 22444 15748 22500 15804
rect 22500 15748 22504 15804
rect 22440 15744 22504 15748
rect 22520 15804 22584 15808
rect 22520 15748 22524 15804
rect 22524 15748 22580 15804
rect 22580 15748 22584 15804
rect 22520 15744 22584 15748
rect 22600 15804 22664 15808
rect 22600 15748 22604 15804
rect 22604 15748 22660 15804
rect 22660 15748 22664 15804
rect 22600 15744 22664 15748
rect 22680 15804 22744 15808
rect 22680 15748 22684 15804
rect 22684 15748 22740 15804
rect 22740 15748 22744 15804
rect 22680 15744 22744 15748
rect 3740 15404 3804 15468
rect 1360 15260 1424 15264
rect 1360 15204 1364 15260
rect 1364 15204 1420 15260
rect 1420 15204 1424 15260
rect 1360 15200 1424 15204
rect 1440 15260 1504 15264
rect 1440 15204 1444 15260
rect 1444 15204 1500 15260
rect 1500 15204 1504 15260
rect 1440 15200 1504 15204
rect 1520 15260 1584 15264
rect 1520 15204 1524 15260
rect 1524 15204 1580 15260
rect 1580 15204 1584 15260
rect 1520 15200 1584 15204
rect 1600 15260 1664 15264
rect 1600 15204 1604 15260
rect 1604 15204 1660 15260
rect 1660 15204 1664 15260
rect 1600 15200 1664 15204
rect 1680 15260 1744 15264
rect 1680 15204 1684 15260
rect 1684 15204 1740 15260
rect 1740 15204 1744 15260
rect 1680 15200 1744 15204
rect 18092 15540 18156 15604
rect 11284 15268 11348 15332
rect 7360 15260 7424 15264
rect 7360 15204 7364 15260
rect 7364 15204 7420 15260
rect 7420 15204 7424 15260
rect 7360 15200 7424 15204
rect 7440 15260 7504 15264
rect 7440 15204 7444 15260
rect 7444 15204 7500 15260
rect 7500 15204 7504 15260
rect 7440 15200 7504 15204
rect 7520 15260 7584 15264
rect 7520 15204 7524 15260
rect 7524 15204 7580 15260
rect 7580 15204 7584 15260
rect 7520 15200 7584 15204
rect 7600 15260 7664 15264
rect 7600 15204 7604 15260
rect 7604 15204 7660 15260
rect 7660 15204 7664 15260
rect 7600 15200 7664 15204
rect 7680 15260 7744 15264
rect 7680 15204 7684 15260
rect 7684 15204 7740 15260
rect 7740 15204 7744 15260
rect 7680 15200 7744 15204
rect 13360 15260 13424 15264
rect 13360 15204 13364 15260
rect 13364 15204 13420 15260
rect 13420 15204 13424 15260
rect 13360 15200 13424 15204
rect 13440 15260 13504 15264
rect 13440 15204 13444 15260
rect 13444 15204 13500 15260
rect 13500 15204 13504 15260
rect 13440 15200 13504 15204
rect 13520 15260 13584 15264
rect 13520 15204 13524 15260
rect 13524 15204 13580 15260
rect 13580 15204 13584 15260
rect 13520 15200 13584 15204
rect 13600 15260 13664 15264
rect 13600 15204 13604 15260
rect 13604 15204 13660 15260
rect 13660 15204 13664 15260
rect 13600 15200 13664 15204
rect 13680 15260 13744 15264
rect 13680 15204 13684 15260
rect 13684 15204 13740 15260
rect 13740 15204 13744 15260
rect 13680 15200 13744 15204
rect 19360 15260 19424 15264
rect 19360 15204 19364 15260
rect 19364 15204 19420 15260
rect 19420 15204 19424 15260
rect 19360 15200 19424 15204
rect 19440 15260 19504 15264
rect 19440 15204 19444 15260
rect 19444 15204 19500 15260
rect 19500 15204 19504 15260
rect 19440 15200 19504 15204
rect 19520 15260 19584 15264
rect 19520 15204 19524 15260
rect 19524 15204 19580 15260
rect 19580 15204 19584 15260
rect 19520 15200 19584 15204
rect 19600 15260 19664 15264
rect 19600 15204 19604 15260
rect 19604 15204 19660 15260
rect 19660 15204 19664 15260
rect 19600 15200 19664 15204
rect 19680 15260 19744 15264
rect 19680 15204 19684 15260
rect 19684 15204 19740 15260
rect 19740 15204 19744 15260
rect 19680 15200 19744 15204
rect 10916 14996 10980 15060
rect 4360 14716 4424 14720
rect 4360 14660 4364 14716
rect 4364 14660 4420 14716
rect 4420 14660 4424 14716
rect 4360 14656 4424 14660
rect 4440 14716 4504 14720
rect 4440 14660 4444 14716
rect 4444 14660 4500 14716
rect 4500 14660 4504 14716
rect 4440 14656 4504 14660
rect 4520 14716 4584 14720
rect 4520 14660 4524 14716
rect 4524 14660 4580 14716
rect 4580 14660 4584 14716
rect 4520 14656 4584 14660
rect 4600 14716 4664 14720
rect 4600 14660 4604 14716
rect 4604 14660 4660 14716
rect 4660 14660 4664 14716
rect 4600 14656 4664 14660
rect 4680 14716 4744 14720
rect 4680 14660 4684 14716
rect 4684 14660 4740 14716
rect 4740 14660 4744 14716
rect 4680 14656 4744 14660
rect 10360 14716 10424 14720
rect 10360 14660 10364 14716
rect 10364 14660 10420 14716
rect 10420 14660 10424 14716
rect 10360 14656 10424 14660
rect 10440 14716 10504 14720
rect 10440 14660 10444 14716
rect 10444 14660 10500 14716
rect 10500 14660 10504 14716
rect 10440 14656 10504 14660
rect 10520 14716 10584 14720
rect 10520 14660 10524 14716
rect 10524 14660 10580 14716
rect 10580 14660 10584 14716
rect 10520 14656 10584 14660
rect 10600 14716 10664 14720
rect 10600 14660 10604 14716
rect 10604 14660 10660 14716
rect 10660 14660 10664 14716
rect 10600 14656 10664 14660
rect 10680 14716 10744 14720
rect 10680 14660 10684 14716
rect 10684 14660 10740 14716
rect 10740 14660 10744 14716
rect 10680 14656 10744 14660
rect 16360 14716 16424 14720
rect 16360 14660 16364 14716
rect 16364 14660 16420 14716
rect 16420 14660 16424 14716
rect 16360 14656 16424 14660
rect 16440 14716 16504 14720
rect 16440 14660 16444 14716
rect 16444 14660 16500 14716
rect 16500 14660 16504 14716
rect 16440 14656 16504 14660
rect 16520 14716 16584 14720
rect 16520 14660 16524 14716
rect 16524 14660 16580 14716
rect 16580 14660 16584 14716
rect 16520 14656 16584 14660
rect 16600 14716 16664 14720
rect 16600 14660 16604 14716
rect 16604 14660 16660 14716
rect 16660 14660 16664 14716
rect 16600 14656 16664 14660
rect 16680 14716 16744 14720
rect 16680 14660 16684 14716
rect 16684 14660 16740 14716
rect 16740 14660 16744 14716
rect 16680 14656 16744 14660
rect 22360 14716 22424 14720
rect 22360 14660 22364 14716
rect 22364 14660 22420 14716
rect 22420 14660 22424 14716
rect 22360 14656 22424 14660
rect 22440 14716 22504 14720
rect 22440 14660 22444 14716
rect 22444 14660 22500 14716
rect 22500 14660 22504 14716
rect 22440 14656 22504 14660
rect 22520 14716 22584 14720
rect 22520 14660 22524 14716
rect 22524 14660 22580 14716
rect 22580 14660 22584 14716
rect 22520 14656 22584 14660
rect 22600 14716 22664 14720
rect 22600 14660 22604 14716
rect 22604 14660 22660 14716
rect 22660 14660 22664 14716
rect 22600 14656 22664 14660
rect 22680 14716 22744 14720
rect 22680 14660 22684 14716
rect 22684 14660 22740 14716
rect 22740 14660 22744 14716
rect 22680 14656 22744 14660
rect 11836 14588 11900 14652
rect 19196 14452 19260 14516
rect 12940 14180 13004 14244
rect 1360 14172 1424 14176
rect 1360 14116 1364 14172
rect 1364 14116 1420 14172
rect 1420 14116 1424 14172
rect 1360 14112 1424 14116
rect 1440 14172 1504 14176
rect 1440 14116 1444 14172
rect 1444 14116 1500 14172
rect 1500 14116 1504 14172
rect 1440 14112 1504 14116
rect 1520 14172 1584 14176
rect 1520 14116 1524 14172
rect 1524 14116 1580 14172
rect 1580 14116 1584 14172
rect 1520 14112 1584 14116
rect 1600 14172 1664 14176
rect 1600 14116 1604 14172
rect 1604 14116 1660 14172
rect 1660 14116 1664 14172
rect 1600 14112 1664 14116
rect 1680 14172 1744 14176
rect 1680 14116 1684 14172
rect 1684 14116 1740 14172
rect 1740 14116 1744 14172
rect 1680 14112 1744 14116
rect 7360 14172 7424 14176
rect 7360 14116 7364 14172
rect 7364 14116 7420 14172
rect 7420 14116 7424 14172
rect 7360 14112 7424 14116
rect 7440 14172 7504 14176
rect 7440 14116 7444 14172
rect 7444 14116 7500 14172
rect 7500 14116 7504 14172
rect 7440 14112 7504 14116
rect 7520 14172 7584 14176
rect 7520 14116 7524 14172
rect 7524 14116 7580 14172
rect 7580 14116 7584 14172
rect 7520 14112 7584 14116
rect 7600 14172 7664 14176
rect 7600 14116 7604 14172
rect 7604 14116 7660 14172
rect 7660 14116 7664 14172
rect 7600 14112 7664 14116
rect 7680 14172 7744 14176
rect 7680 14116 7684 14172
rect 7684 14116 7740 14172
rect 7740 14116 7744 14172
rect 7680 14112 7744 14116
rect 13360 14172 13424 14176
rect 13360 14116 13364 14172
rect 13364 14116 13420 14172
rect 13420 14116 13424 14172
rect 13360 14112 13424 14116
rect 13440 14172 13504 14176
rect 13440 14116 13444 14172
rect 13444 14116 13500 14172
rect 13500 14116 13504 14172
rect 13440 14112 13504 14116
rect 13520 14172 13584 14176
rect 13520 14116 13524 14172
rect 13524 14116 13580 14172
rect 13580 14116 13584 14172
rect 13520 14112 13584 14116
rect 13600 14172 13664 14176
rect 13600 14116 13604 14172
rect 13604 14116 13660 14172
rect 13660 14116 13664 14172
rect 13600 14112 13664 14116
rect 13680 14172 13744 14176
rect 13680 14116 13684 14172
rect 13684 14116 13740 14172
rect 13740 14116 13744 14172
rect 13680 14112 13744 14116
rect 19360 14172 19424 14176
rect 19360 14116 19364 14172
rect 19364 14116 19420 14172
rect 19420 14116 19424 14172
rect 19360 14112 19424 14116
rect 19440 14172 19504 14176
rect 19440 14116 19444 14172
rect 19444 14116 19500 14172
rect 19500 14116 19504 14172
rect 19440 14112 19504 14116
rect 19520 14172 19584 14176
rect 19520 14116 19524 14172
rect 19524 14116 19580 14172
rect 19580 14116 19584 14172
rect 19520 14112 19584 14116
rect 19600 14172 19664 14176
rect 19600 14116 19604 14172
rect 19604 14116 19660 14172
rect 19660 14116 19664 14172
rect 19600 14112 19664 14116
rect 19680 14172 19744 14176
rect 19680 14116 19684 14172
rect 19684 14116 19740 14172
rect 19740 14116 19744 14172
rect 19680 14112 19744 14116
rect 5948 13772 6012 13836
rect 9076 13636 9140 13700
rect 4360 13628 4424 13632
rect 4360 13572 4364 13628
rect 4364 13572 4420 13628
rect 4420 13572 4424 13628
rect 4360 13568 4424 13572
rect 4440 13628 4504 13632
rect 4440 13572 4444 13628
rect 4444 13572 4500 13628
rect 4500 13572 4504 13628
rect 4440 13568 4504 13572
rect 4520 13628 4584 13632
rect 4520 13572 4524 13628
rect 4524 13572 4580 13628
rect 4580 13572 4584 13628
rect 4520 13568 4584 13572
rect 4600 13628 4664 13632
rect 4600 13572 4604 13628
rect 4604 13572 4660 13628
rect 4660 13572 4664 13628
rect 4600 13568 4664 13572
rect 4680 13628 4744 13632
rect 4680 13572 4684 13628
rect 4684 13572 4740 13628
rect 4740 13572 4744 13628
rect 4680 13568 4744 13572
rect 10360 13628 10424 13632
rect 10360 13572 10364 13628
rect 10364 13572 10420 13628
rect 10420 13572 10424 13628
rect 10360 13568 10424 13572
rect 10440 13628 10504 13632
rect 10440 13572 10444 13628
rect 10444 13572 10500 13628
rect 10500 13572 10504 13628
rect 10440 13568 10504 13572
rect 10520 13628 10584 13632
rect 10520 13572 10524 13628
rect 10524 13572 10580 13628
rect 10580 13572 10584 13628
rect 10520 13568 10584 13572
rect 10600 13628 10664 13632
rect 10600 13572 10604 13628
rect 10604 13572 10660 13628
rect 10660 13572 10664 13628
rect 10600 13568 10664 13572
rect 10680 13628 10744 13632
rect 10680 13572 10684 13628
rect 10684 13572 10740 13628
rect 10740 13572 10744 13628
rect 10680 13568 10744 13572
rect 16360 13628 16424 13632
rect 16360 13572 16364 13628
rect 16364 13572 16420 13628
rect 16420 13572 16424 13628
rect 16360 13568 16424 13572
rect 16440 13628 16504 13632
rect 16440 13572 16444 13628
rect 16444 13572 16500 13628
rect 16500 13572 16504 13628
rect 16440 13568 16504 13572
rect 16520 13628 16584 13632
rect 16520 13572 16524 13628
rect 16524 13572 16580 13628
rect 16580 13572 16584 13628
rect 16520 13568 16584 13572
rect 16600 13628 16664 13632
rect 16600 13572 16604 13628
rect 16604 13572 16660 13628
rect 16660 13572 16664 13628
rect 16600 13568 16664 13572
rect 16680 13628 16744 13632
rect 16680 13572 16684 13628
rect 16684 13572 16740 13628
rect 16740 13572 16744 13628
rect 16680 13568 16744 13572
rect 22360 13628 22424 13632
rect 22360 13572 22364 13628
rect 22364 13572 22420 13628
rect 22420 13572 22424 13628
rect 22360 13568 22424 13572
rect 22440 13628 22504 13632
rect 22440 13572 22444 13628
rect 22444 13572 22500 13628
rect 22500 13572 22504 13628
rect 22440 13568 22504 13572
rect 22520 13628 22584 13632
rect 22520 13572 22524 13628
rect 22524 13572 22580 13628
rect 22580 13572 22584 13628
rect 22520 13568 22584 13572
rect 22600 13628 22664 13632
rect 22600 13572 22604 13628
rect 22604 13572 22660 13628
rect 22660 13572 22664 13628
rect 22600 13568 22664 13572
rect 22680 13628 22744 13632
rect 22680 13572 22684 13628
rect 22684 13572 22740 13628
rect 22740 13572 22744 13628
rect 22680 13568 22744 13572
rect 7972 13500 8036 13564
rect 12756 13424 12820 13428
rect 12756 13368 12806 13424
rect 12806 13368 12820 13424
rect 12756 13364 12820 13368
rect 11652 13228 11716 13292
rect 18460 13228 18524 13292
rect 13124 13092 13188 13156
rect 1360 13084 1424 13088
rect 1360 13028 1364 13084
rect 1364 13028 1420 13084
rect 1420 13028 1424 13084
rect 1360 13024 1424 13028
rect 1440 13084 1504 13088
rect 1440 13028 1444 13084
rect 1444 13028 1500 13084
rect 1500 13028 1504 13084
rect 1440 13024 1504 13028
rect 1520 13084 1584 13088
rect 1520 13028 1524 13084
rect 1524 13028 1580 13084
rect 1580 13028 1584 13084
rect 1520 13024 1584 13028
rect 1600 13084 1664 13088
rect 1600 13028 1604 13084
rect 1604 13028 1660 13084
rect 1660 13028 1664 13084
rect 1600 13024 1664 13028
rect 1680 13084 1744 13088
rect 1680 13028 1684 13084
rect 1684 13028 1740 13084
rect 1740 13028 1744 13084
rect 1680 13024 1744 13028
rect 7360 13084 7424 13088
rect 7360 13028 7364 13084
rect 7364 13028 7420 13084
rect 7420 13028 7424 13084
rect 7360 13024 7424 13028
rect 7440 13084 7504 13088
rect 7440 13028 7444 13084
rect 7444 13028 7500 13084
rect 7500 13028 7504 13084
rect 7440 13024 7504 13028
rect 7520 13084 7584 13088
rect 7520 13028 7524 13084
rect 7524 13028 7580 13084
rect 7580 13028 7584 13084
rect 7520 13024 7584 13028
rect 7600 13084 7664 13088
rect 7600 13028 7604 13084
rect 7604 13028 7660 13084
rect 7660 13028 7664 13084
rect 7600 13024 7664 13028
rect 7680 13084 7744 13088
rect 7680 13028 7684 13084
rect 7684 13028 7740 13084
rect 7740 13028 7744 13084
rect 7680 13024 7744 13028
rect 13360 13084 13424 13088
rect 13360 13028 13364 13084
rect 13364 13028 13420 13084
rect 13420 13028 13424 13084
rect 13360 13024 13424 13028
rect 13440 13084 13504 13088
rect 13440 13028 13444 13084
rect 13444 13028 13500 13084
rect 13500 13028 13504 13084
rect 13440 13024 13504 13028
rect 13520 13084 13584 13088
rect 13520 13028 13524 13084
rect 13524 13028 13580 13084
rect 13580 13028 13584 13084
rect 13520 13024 13584 13028
rect 13600 13084 13664 13088
rect 13600 13028 13604 13084
rect 13604 13028 13660 13084
rect 13660 13028 13664 13084
rect 13600 13024 13664 13028
rect 13680 13084 13744 13088
rect 13680 13028 13684 13084
rect 13684 13028 13740 13084
rect 13740 13028 13744 13084
rect 13680 13024 13744 13028
rect 19360 13084 19424 13088
rect 19360 13028 19364 13084
rect 19364 13028 19420 13084
rect 19420 13028 19424 13084
rect 19360 13024 19424 13028
rect 19440 13084 19504 13088
rect 19440 13028 19444 13084
rect 19444 13028 19500 13084
rect 19500 13028 19504 13084
rect 19440 13024 19504 13028
rect 19520 13084 19584 13088
rect 19520 13028 19524 13084
rect 19524 13028 19580 13084
rect 19580 13028 19584 13084
rect 19520 13024 19584 13028
rect 19600 13084 19664 13088
rect 19600 13028 19604 13084
rect 19604 13028 19660 13084
rect 19660 13028 19664 13084
rect 19600 13024 19664 13028
rect 19680 13084 19744 13088
rect 19680 13028 19684 13084
rect 19684 13028 19740 13084
rect 19740 13028 19744 13084
rect 19680 13024 19744 13028
rect 9260 12820 9324 12884
rect 20852 12880 20916 12884
rect 20852 12824 20866 12880
rect 20866 12824 20916 12880
rect 20852 12820 20916 12824
rect 21220 12820 21284 12884
rect 12572 12548 12636 12612
rect 4360 12540 4424 12544
rect 4360 12484 4364 12540
rect 4364 12484 4420 12540
rect 4420 12484 4424 12540
rect 4360 12480 4424 12484
rect 4440 12540 4504 12544
rect 4440 12484 4444 12540
rect 4444 12484 4500 12540
rect 4500 12484 4504 12540
rect 4440 12480 4504 12484
rect 4520 12540 4584 12544
rect 4520 12484 4524 12540
rect 4524 12484 4580 12540
rect 4580 12484 4584 12540
rect 4520 12480 4584 12484
rect 4600 12540 4664 12544
rect 4600 12484 4604 12540
rect 4604 12484 4660 12540
rect 4660 12484 4664 12540
rect 4600 12480 4664 12484
rect 4680 12540 4744 12544
rect 4680 12484 4684 12540
rect 4684 12484 4740 12540
rect 4740 12484 4744 12540
rect 4680 12480 4744 12484
rect 10360 12540 10424 12544
rect 10360 12484 10364 12540
rect 10364 12484 10420 12540
rect 10420 12484 10424 12540
rect 10360 12480 10424 12484
rect 10440 12540 10504 12544
rect 10440 12484 10444 12540
rect 10444 12484 10500 12540
rect 10500 12484 10504 12540
rect 10440 12480 10504 12484
rect 10520 12540 10584 12544
rect 10520 12484 10524 12540
rect 10524 12484 10580 12540
rect 10580 12484 10584 12540
rect 10520 12480 10584 12484
rect 10600 12540 10664 12544
rect 10600 12484 10604 12540
rect 10604 12484 10660 12540
rect 10660 12484 10664 12540
rect 10600 12480 10664 12484
rect 10680 12540 10744 12544
rect 10680 12484 10684 12540
rect 10684 12484 10740 12540
rect 10740 12484 10744 12540
rect 10680 12480 10744 12484
rect 16360 12540 16424 12544
rect 16360 12484 16364 12540
rect 16364 12484 16420 12540
rect 16420 12484 16424 12540
rect 16360 12480 16424 12484
rect 16440 12540 16504 12544
rect 16440 12484 16444 12540
rect 16444 12484 16500 12540
rect 16500 12484 16504 12540
rect 16440 12480 16504 12484
rect 16520 12540 16584 12544
rect 16520 12484 16524 12540
rect 16524 12484 16580 12540
rect 16580 12484 16584 12540
rect 16520 12480 16584 12484
rect 16600 12540 16664 12544
rect 16600 12484 16604 12540
rect 16604 12484 16660 12540
rect 16660 12484 16664 12540
rect 16600 12480 16664 12484
rect 16680 12540 16744 12544
rect 16680 12484 16684 12540
rect 16684 12484 16740 12540
rect 16740 12484 16744 12540
rect 16680 12480 16744 12484
rect 22360 12540 22424 12544
rect 22360 12484 22364 12540
rect 22364 12484 22420 12540
rect 22420 12484 22424 12540
rect 22360 12480 22424 12484
rect 22440 12540 22504 12544
rect 22440 12484 22444 12540
rect 22444 12484 22500 12540
rect 22500 12484 22504 12540
rect 22440 12480 22504 12484
rect 22520 12540 22584 12544
rect 22520 12484 22524 12540
rect 22524 12484 22580 12540
rect 22580 12484 22584 12540
rect 22520 12480 22584 12484
rect 22600 12540 22664 12544
rect 22600 12484 22604 12540
rect 22604 12484 22660 12540
rect 22660 12484 22664 12540
rect 22600 12480 22664 12484
rect 22680 12540 22744 12544
rect 22680 12484 22684 12540
rect 22684 12484 22740 12540
rect 22740 12484 22744 12540
rect 22680 12480 22744 12484
rect 12940 12140 13004 12204
rect 10916 12004 10980 12068
rect 1360 11996 1424 12000
rect 1360 11940 1364 11996
rect 1364 11940 1420 11996
rect 1420 11940 1424 11996
rect 1360 11936 1424 11940
rect 1440 11996 1504 12000
rect 1440 11940 1444 11996
rect 1444 11940 1500 11996
rect 1500 11940 1504 11996
rect 1440 11936 1504 11940
rect 1520 11996 1584 12000
rect 1520 11940 1524 11996
rect 1524 11940 1580 11996
rect 1580 11940 1584 11996
rect 1520 11936 1584 11940
rect 1600 11996 1664 12000
rect 1600 11940 1604 11996
rect 1604 11940 1660 11996
rect 1660 11940 1664 11996
rect 1600 11936 1664 11940
rect 1680 11996 1744 12000
rect 1680 11940 1684 11996
rect 1684 11940 1740 11996
rect 1740 11940 1744 11996
rect 1680 11936 1744 11940
rect 7360 11996 7424 12000
rect 7360 11940 7364 11996
rect 7364 11940 7420 11996
rect 7420 11940 7424 11996
rect 7360 11936 7424 11940
rect 7440 11996 7504 12000
rect 7440 11940 7444 11996
rect 7444 11940 7500 11996
rect 7500 11940 7504 11996
rect 7440 11936 7504 11940
rect 7520 11996 7584 12000
rect 7520 11940 7524 11996
rect 7524 11940 7580 11996
rect 7580 11940 7584 11996
rect 7520 11936 7584 11940
rect 7600 11996 7664 12000
rect 7600 11940 7604 11996
rect 7604 11940 7660 11996
rect 7660 11940 7664 11996
rect 7600 11936 7664 11940
rect 7680 11996 7744 12000
rect 7680 11940 7684 11996
rect 7684 11940 7740 11996
rect 7740 11940 7744 11996
rect 7680 11936 7744 11940
rect 13360 11996 13424 12000
rect 13360 11940 13364 11996
rect 13364 11940 13420 11996
rect 13420 11940 13424 11996
rect 13360 11936 13424 11940
rect 13440 11996 13504 12000
rect 13440 11940 13444 11996
rect 13444 11940 13500 11996
rect 13500 11940 13504 11996
rect 13440 11936 13504 11940
rect 13520 11996 13584 12000
rect 13520 11940 13524 11996
rect 13524 11940 13580 11996
rect 13580 11940 13584 11996
rect 13520 11936 13584 11940
rect 13600 11996 13664 12000
rect 13600 11940 13604 11996
rect 13604 11940 13660 11996
rect 13660 11940 13664 11996
rect 13600 11936 13664 11940
rect 13680 11996 13744 12000
rect 13680 11940 13684 11996
rect 13684 11940 13740 11996
rect 13740 11940 13744 11996
rect 13680 11936 13744 11940
rect 19360 11996 19424 12000
rect 19360 11940 19364 11996
rect 19364 11940 19420 11996
rect 19420 11940 19424 11996
rect 19360 11936 19424 11940
rect 19440 11996 19504 12000
rect 19440 11940 19444 11996
rect 19444 11940 19500 11996
rect 19500 11940 19504 11996
rect 19440 11936 19504 11940
rect 19520 11996 19584 12000
rect 19520 11940 19524 11996
rect 19524 11940 19580 11996
rect 19580 11940 19584 11996
rect 19520 11936 19584 11940
rect 19600 11996 19664 12000
rect 19600 11940 19604 11996
rect 19604 11940 19660 11996
rect 19660 11940 19664 11996
rect 19600 11936 19664 11940
rect 19680 11996 19744 12000
rect 19680 11940 19684 11996
rect 19684 11940 19740 11996
rect 19740 11940 19744 11996
rect 19680 11936 19744 11940
rect 11284 11732 11348 11796
rect 20668 12200 20732 12204
rect 20668 12144 20682 12200
rect 20682 12144 20732 12200
rect 20668 12140 20732 12144
rect 10180 11596 10244 11660
rect 11284 11596 11348 11660
rect 12572 11520 12636 11524
rect 12572 11464 12586 11520
rect 12586 11464 12636 11520
rect 12572 11460 12636 11464
rect 4360 11452 4424 11456
rect 4360 11396 4364 11452
rect 4364 11396 4420 11452
rect 4420 11396 4424 11452
rect 4360 11392 4424 11396
rect 4440 11452 4504 11456
rect 4440 11396 4444 11452
rect 4444 11396 4500 11452
rect 4500 11396 4504 11452
rect 4440 11392 4504 11396
rect 4520 11452 4584 11456
rect 4520 11396 4524 11452
rect 4524 11396 4580 11452
rect 4580 11396 4584 11452
rect 4520 11392 4584 11396
rect 4600 11452 4664 11456
rect 4600 11396 4604 11452
rect 4604 11396 4660 11452
rect 4660 11396 4664 11452
rect 4600 11392 4664 11396
rect 4680 11452 4744 11456
rect 4680 11396 4684 11452
rect 4684 11396 4740 11452
rect 4740 11396 4744 11452
rect 4680 11392 4744 11396
rect 10360 11452 10424 11456
rect 10360 11396 10364 11452
rect 10364 11396 10420 11452
rect 10420 11396 10424 11452
rect 10360 11392 10424 11396
rect 10440 11452 10504 11456
rect 10440 11396 10444 11452
rect 10444 11396 10500 11452
rect 10500 11396 10504 11452
rect 10440 11392 10504 11396
rect 10520 11452 10584 11456
rect 10520 11396 10524 11452
rect 10524 11396 10580 11452
rect 10580 11396 10584 11452
rect 10520 11392 10584 11396
rect 10600 11452 10664 11456
rect 10600 11396 10604 11452
rect 10604 11396 10660 11452
rect 10660 11396 10664 11452
rect 10600 11392 10664 11396
rect 10680 11452 10744 11456
rect 10680 11396 10684 11452
rect 10684 11396 10740 11452
rect 10740 11396 10744 11452
rect 10680 11392 10744 11396
rect 16360 11452 16424 11456
rect 16360 11396 16364 11452
rect 16364 11396 16420 11452
rect 16420 11396 16424 11452
rect 16360 11392 16424 11396
rect 16440 11452 16504 11456
rect 16440 11396 16444 11452
rect 16444 11396 16500 11452
rect 16500 11396 16504 11452
rect 16440 11392 16504 11396
rect 16520 11452 16584 11456
rect 16520 11396 16524 11452
rect 16524 11396 16580 11452
rect 16580 11396 16584 11452
rect 16520 11392 16584 11396
rect 16600 11452 16664 11456
rect 16600 11396 16604 11452
rect 16604 11396 16660 11452
rect 16660 11396 16664 11452
rect 16600 11392 16664 11396
rect 16680 11452 16744 11456
rect 16680 11396 16684 11452
rect 16684 11396 16740 11452
rect 16740 11396 16744 11452
rect 16680 11392 16744 11396
rect 22360 11452 22424 11456
rect 22360 11396 22364 11452
rect 22364 11396 22420 11452
rect 22420 11396 22424 11452
rect 22360 11392 22424 11396
rect 22440 11452 22504 11456
rect 22440 11396 22444 11452
rect 22444 11396 22500 11452
rect 22500 11396 22504 11452
rect 22440 11392 22504 11396
rect 22520 11452 22584 11456
rect 22520 11396 22524 11452
rect 22524 11396 22580 11452
rect 22580 11396 22584 11452
rect 22520 11392 22584 11396
rect 22600 11452 22664 11456
rect 22600 11396 22604 11452
rect 22604 11396 22660 11452
rect 22660 11396 22664 11452
rect 22600 11392 22664 11396
rect 22680 11452 22744 11456
rect 22680 11396 22684 11452
rect 22684 11396 22740 11452
rect 22740 11396 22744 11452
rect 22680 11392 22744 11396
rect 5028 11052 5092 11116
rect 12020 11052 12084 11116
rect 7972 10916 8036 10980
rect 1360 10908 1424 10912
rect 1360 10852 1364 10908
rect 1364 10852 1420 10908
rect 1420 10852 1424 10908
rect 1360 10848 1424 10852
rect 1440 10908 1504 10912
rect 1440 10852 1444 10908
rect 1444 10852 1500 10908
rect 1500 10852 1504 10908
rect 1440 10848 1504 10852
rect 1520 10908 1584 10912
rect 1520 10852 1524 10908
rect 1524 10852 1580 10908
rect 1580 10852 1584 10908
rect 1520 10848 1584 10852
rect 1600 10908 1664 10912
rect 1600 10852 1604 10908
rect 1604 10852 1660 10908
rect 1660 10852 1664 10908
rect 1600 10848 1664 10852
rect 1680 10908 1744 10912
rect 1680 10852 1684 10908
rect 1684 10852 1740 10908
rect 1740 10852 1744 10908
rect 1680 10848 1744 10852
rect 7360 10908 7424 10912
rect 7360 10852 7364 10908
rect 7364 10852 7420 10908
rect 7420 10852 7424 10908
rect 7360 10848 7424 10852
rect 7440 10908 7504 10912
rect 7440 10852 7444 10908
rect 7444 10852 7500 10908
rect 7500 10852 7504 10908
rect 7440 10848 7504 10852
rect 7520 10908 7584 10912
rect 7520 10852 7524 10908
rect 7524 10852 7580 10908
rect 7580 10852 7584 10908
rect 7520 10848 7584 10852
rect 7600 10908 7664 10912
rect 7600 10852 7604 10908
rect 7604 10852 7660 10908
rect 7660 10852 7664 10908
rect 7600 10848 7664 10852
rect 7680 10908 7744 10912
rect 7680 10852 7684 10908
rect 7684 10852 7740 10908
rect 7740 10852 7744 10908
rect 7680 10848 7744 10852
rect 13360 10908 13424 10912
rect 13360 10852 13364 10908
rect 13364 10852 13420 10908
rect 13420 10852 13424 10908
rect 13360 10848 13424 10852
rect 13440 10908 13504 10912
rect 13440 10852 13444 10908
rect 13444 10852 13500 10908
rect 13500 10852 13504 10908
rect 13440 10848 13504 10852
rect 13520 10908 13584 10912
rect 13520 10852 13524 10908
rect 13524 10852 13580 10908
rect 13580 10852 13584 10908
rect 13520 10848 13584 10852
rect 13600 10908 13664 10912
rect 13600 10852 13604 10908
rect 13604 10852 13660 10908
rect 13660 10852 13664 10908
rect 13600 10848 13664 10852
rect 13680 10908 13744 10912
rect 13680 10852 13684 10908
rect 13684 10852 13740 10908
rect 13740 10852 13744 10908
rect 13680 10848 13744 10852
rect 19360 10908 19424 10912
rect 19360 10852 19364 10908
rect 19364 10852 19420 10908
rect 19420 10852 19424 10908
rect 19360 10848 19424 10852
rect 19440 10908 19504 10912
rect 19440 10852 19444 10908
rect 19444 10852 19500 10908
rect 19500 10852 19504 10908
rect 19440 10848 19504 10852
rect 19520 10908 19584 10912
rect 19520 10852 19524 10908
rect 19524 10852 19580 10908
rect 19580 10852 19584 10908
rect 19520 10848 19584 10852
rect 19600 10908 19664 10912
rect 19600 10852 19604 10908
rect 19604 10852 19660 10908
rect 19660 10852 19664 10908
rect 19600 10848 19664 10852
rect 19680 10908 19744 10912
rect 19680 10852 19684 10908
rect 19684 10852 19740 10908
rect 19740 10852 19744 10908
rect 19680 10848 19744 10852
rect 6684 10644 6748 10708
rect 19196 10704 19260 10708
rect 19196 10648 19246 10704
rect 19246 10648 19260 10704
rect 19196 10644 19260 10648
rect 4360 10364 4424 10368
rect 4360 10308 4364 10364
rect 4364 10308 4420 10364
rect 4420 10308 4424 10364
rect 4360 10304 4424 10308
rect 4440 10364 4504 10368
rect 4440 10308 4444 10364
rect 4444 10308 4500 10364
rect 4500 10308 4504 10364
rect 4440 10304 4504 10308
rect 4520 10364 4584 10368
rect 4520 10308 4524 10364
rect 4524 10308 4580 10364
rect 4580 10308 4584 10364
rect 4520 10304 4584 10308
rect 4600 10364 4664 10368
rect 4600 10308 4604 10364
rect 4604 10308 4660 10364
rect 4660 10308 4664 10364
rect 4600 10304 4664 10308
rect 4680 10364 4744 10368
rect 4680 10308 4684 10364
rect 4684 10308 4740 10364
rect 4740 10308 4744 10364
rect 4680 10304 4744 10308
rect 10360 10364 10424 10368
rect 10360 10308 10364 10364
rect 10364 10308 10420 10364
rect 10420 10308 10424 10364
rect 10360 10304 10424 10308
rect 10440 10364 10504 10368
rect 10440 10308 10444 10364
rect 10444 10308 10500 10364
rect 10500 10308 10504 10364
rect 10440 10304 10504 10308
rect 10520 10364 10584 10368
rect 10520 10308 10524 10364
rect 10524 10308 10580 10364
rect 10580 10308 10584 10364
rect 10520 10304 10584 10308
rect 10600 10364 10664 10368
rect 10600 10308 10604 10364
rect 10604 10308 10660 10364
rect 10660 10308 10664 10364
rect 10600 10304 10664 10308
rect 10680 10364 10744 10368
rect 10680 10308 10684 10364
rect 10684 10308 10740 10364
rect 10740 10308 10744 10364
rect 10680 10304 10744 10308
rect 12388 10508 12452 10572
rect 13124 10508 13188 10572
rect 16360 10364 16424 10368
rect 16360 10308 16364 10364
rect 16364 10308 16420 10364
rect 16420 10308 16424 10364
rect 16360 10304 16424 10308
rect 16440 10364 16504 10368
rect 16440 10308 16444 10364
rect 16444 10308 16500 10364
rect 16500 10308 16504 10364
rect 16440 10304 16504 10308
rect 16520 10364 16584 10368
rect 16520 10308 16524 10364
rect 16524 10308 16580 10364
rect 16580 10308 16584 10364
rect 16520 10304 16584 10308
rect 16600 10364 16664 10368
rect 16600 10308 16604 10364
rect 16604 10308 16660 10364
rect 16660 10308 16664 10364
rect 16600 10304 16664 10308
rect 16680 10364 16744 10368
rect 16680 10308 16684 10364
rect 16684 10308 16740 10364
rect 16740 10308 16744 10364
rect 16680 10304 16744 10308
rect 22360 10364 22424 10368
rect 22360 10308 22364 10364
rect 22364 10308 22420 10364
rect 22420 10308 22424 10364
rect 22360 10304 22424 10308
rect 22440 10364 22504 10368
rect 22440 10308 22444 10364
rect 22444 10308 22500 10364
rect 22500 10308 22504 10364
rect 22440 10304 22504 10308
rect 22520 10364 22584 10368
rect 22520 10308 22524 10364
rect 22524 10308 22580 10364
rect 22580 10308 22584 10364
rect 22520 10304 22584 10308
rect 22600 10364 22664 10368
rect 22600 10308 22604 10364
rect 22604 10308 22660 10364
rect 22660 10308 22664 10364
rect 22600 10304 22664 10308
rect 22680 10364 22744 10368
rect 22680 10308 22684 10364
rect 22684 10308 22740 10364
rect 22740 10308 22744 10364
rect 22680 10304 22744 10308
rect 18828 9964 18892 10028
rect 19932 9964 19996 10028
rect 1360 9820 1424 9824
rect 1360 9764 1364 9820
rect 1364 9764 1420 9820
rect 1420 9764 1424 9820
rect 1360 9760 1424 9764
rect 1440 9820 1504 9824
rect 1440 9764 1444 9820
rect 1444 9764 1500 9820
rect 1500 9764 1504 9820
rect 1440 9760 1504 9764
rect 1520 9820 1584 9824
rect 1520 9764 1524 9820
rect 1524 9764 1580 9820
rect 1580 9764 1584 9820
rect 1520 9760 1584 9764
rect 1600 9820 1664 9824
rect 1600 9764 1604 9820
rect 1604 9764 1660 9820
rect 1660 9764 1664 9820
rect 1600 9760 1664 9764
rect 1680 9820 1744 9824
rect 1680 9764 1684 9820
rect 1684 9764 1740 9820
rect 1740 9764 1744 9820
rect 1680 9760 1744 9764
rect 7360 9820 7424 9824
rect 7360 9764 7364 9820
rect 7364 9764 7420 9820
rect 7420 9764 7424 9820
rect 7360 9760 7424 9764
rect 7440 9820 7504 9824
rect 7440 9764 7444 9820
rect 7444 9764 7500 9820
rect 7500 9764 7504 9820
rect 7440 9760 7504 9764
rect 7520 9820 7584 9824
rect 7520 9764 7524 9820
rect 7524 9764 7580 9820
rect 7580 9764 7584 9820
rect 7520 9760 7584 9764
rect 7600 9820 7664 9824
rect 7600 9764 7604 9820
rect 7604 9764 7660 9820
rect 7660 9764 7664 9820
rect 7600 9760 7664 9764
rect 7680 9820 7744 9824
rect 7680 9764 7684 9820
rect 7684 9764 7740 9820
rect 7740 9764 7744 9820
rect 7680 9760 7744 9764
rect 9628 9692 9692 9756
rect 13360 9820 13424 9824
rect 13360 9764 13364 9820
rect 13364 9764 13420 9820
rect 13420 9764 13424 9820
rect 13360 9760 13424 9764
rect 13440 9820 13504 9824
rect 13440 9764 13444 9820
rect 13444 9764 13500 9820
rect 13500 9764 13504 9820
rect 13440 9760 13504 9764
rect 13520 9820 13584 9824
rect 13520 9764 13524 9820
rect 13524 9764 13580 9820
rect 13580 9764 13584 9820
rect 13520 9760 13584 9764
rect 13600 9820 13664 9824
rect 13600 9764 13604 9820
rect 13604 9764 13660 9820
rect 13660 9764 13664 9820
rect 13600 9760 13664 9764
rect 13680 9820 13744 9824
rect 13680 9764 13684 9820
rect 13684 9764 13740 9820
rect 13740 9764 13744 9820
rect 13680 9760 13744 9764
rect 19360 9820 19424 9824
rect 19360 9764 19364 9820
rect 19364 9764 19420 9820
rect 19420 9764 19424 9820
rect 19360 9760 19424 9764
rect 19440 9820 19504 9824
rect 19440 9764 19444 9820
rect 19444 9764 19500 9820
rect 19500 9764 19504 9820
rect 19440 9760 19504 9764
rect 19520 9820 19584 9824
rect 19520 9764 19524 9820
rect 19524 9764 19580 9820
rect 19580 9764 19584 9820
rect 19520 9760 19584 9764
rect 19600 9820 19664 9824
rect 19600 9764 19604 9820
rect 19604 9764 19660 9820
rect 19660 9764 19664 9820
rect 19600 9760 19664 9764
rect 19680 9820 19744 9824
rect 19680 9764 19684 9820
rect 19684 9764 19740 9820
rect 19740 9764 19744 9820
rect 19680 9760 19744 9764
rect 18276 9752 18340 9756
rect 18276 9696 18290 9752
rect 18290 9696 18340 9752
rect 18276 9692 18340 9696
rect 13124 9556 13188 9620
rect 4360 9276 4424 9280
rect 4360 9220 4364 9276
rect 4364 9220 4420 9276
rect 4420 9220 4424 9276
rect 4360 9216 4424 9220
rect 4440 9276 4504 9280
rect 4440 9220 4444 9276
rect 4444 9220 4500 9276
rect 4500 9220 4504 9276
rect 4440 9216 4504 9220
rect 4520 9276 4584 9280
rect 4520 9220 4524 9276
rect 4524 9220 4580 9276
rect 4580 9220 4584 9276
rect 4520 9216 4584 9220
rect 4600 9276 4664 9280
rect 4600 9220 4604 9276
rect 4604 9220 4660 9276
rect 4660 9220 4664 9276
rect 4600 9216 4664 9220
rect 4680 9276 4744 9280
rect 4680 9220 4684 9276
rect 4684 9220 4740 9276
rect 4740 9220 4744 9276
rect 4680 9216 4744 9220
rect 10360 9276 10424 9280
rect 10360 9220 10364 9276
rect 10364 9220 10420 9276
rect 10420 9220 10424 9276
rect 10360 9216 10424 9220
rect 10440 9276 10504 9280
rect 10440 9220 10444 9276
rect 10444 9220 10500 9276
rect 10500 9220 10504 9276
rect 10440 9216 10504 9220
rect 10520 9276 10584 9280
rect 10520 9220 10524 9276
rect 10524 9220 10580 9276
rect 10580 9220 10584 9276
rect 10520 9216 10584 9220
rect 10600 9276 10664 9280
rect 10600 9220 10604 9276
rect 10604 9220 10660 9276
rect 10660 9220 10664 9276
rect 10600 9216 10664 9220
rect 10680 9276 10744 9280
rect 10680 9220 10684 9276
rect 10684 9220 10740 9276
rect 10740 9220 10744 9276
rect 10680 9216 10744 9220
rect 7052 9148 7116 9212
rect 10916 9148 10980 9212
rect 14964 9012 15028 9076
rect 16360 9276 16424 9280
rect 16360 9220 16364 9276
rect 16364 9220 16420 9276
rect 16420 9220 16424 9276
rect 16360 9216 16424 9220
rect 16440 9276 16504 9280
rect 16440 9220 16444 9276
rect 16444 9220 16500 9276
rect 16500 9220 16504 9276
rect 16440 9216 16504 9220
rect 16520 9276 16584 9280
rect 16520 9220 16524 9276
rect 16524 9220 16580 9276
rect 16580 9220 16584 9276
rect 16520 9216 16584 9220
rect 16600 9276 16664 9280
rect 16600 9220 16604 9276
rect 16604 9220 16660 9276
rect 16660 9220 16664 9276
rect 16600 9216 16664 9220
rect 16680 9276 16744 9280
rect 16680 9220 16684 9276
rect 16684 9220 16740 9276
rect 16740 9220 16744 9276
rect 16680 9216 16744 9220
rect 22360 9276 22424 9280
rect 22360 9220 22364 9276
rect 22364 9220 22420 9276
rect 22420 9220 22424 9276
rect 22360 9216 22424 9220
rect 22440 9276 22504 9280
rect 22440 9220 22444 9276
rect 22444 9220 22500 9276
rect 22500 9220 22504 9276
rect 22440 9216 22504 9220
rect 22520 9276 22584 9280
rect 22520 9220 22524 9276
rect 22524 9220 22580 9276
rect 22580 9220 22584 9276
rect 22520 9216 22584 9220
rect 22600 9276 22664 9280
rect 22600 9220 22604 9276
rect 22604 9220 22660 9276
rect 22660 9220 22664 9276
rect 22600 9216 22664 9220
rect 22680 9276 22744 9280
rect 22680 9220 22684 9276
rect 22684 9220 22740 9276
rect 22740 9220 22744 9276
rect 22680 9216 22744 9220
rect 20300 9148 20364 9212
rect 18276 8936 18340 8940
rect 18276 8880 18290 8936
rect 18290 8880 18340 8936
rect 18276 8876 18340 8880
rect 13124 8740 13188 8804
rect 1360 8732 1424 8736
rect 1360 8676 1364 8732
rect 1364 8676 1420 8732
rect 1420 8676 1424 8732
rect 1360 8672 1424 8676
rect 1440 8732 1504 8736
rect 1440 8676 1444 8732
rect 1444 8676 1500 8732
rect 1500 8676 1504 8732
rect 1440 8672 1504 8676
rect 1520 8732 1584 8736
rect 1520 8676 1524 8732
rect 1524 8676 1580 8732
rect 1580 8676 1584 8732
rect 1520 8672 1584 8676
rect 1600 8732 1664 8736
rect 1600 8676 1604 8732
rect 1604 8676 1660 8732
rect 1660 8676 1664 8732
rect 1600 8672 1664 8676
rect 1680 8732 1744 8736
rect 1680 8676 1684 8732
rect 1684 8676 1740 8732
rect 1740 8676 1744 8732
rect 1680 8672 1744 8676
rect 7360 8732 7424 8736
rect 7360 8676 7364 8732
rect 7364 8676 7420 8732
rect 7420 8676 7424 8732
rect 7360 8672 7424 8676
rect 7440 8732 7504 8736
rect 7440 8676 7444 8732
rect 7444 8676 7500 8732
rect 7500 8676 7504 8732
rect 7440 8672 7504 8676
rect 7520 8732 7584 8736
rect 7520 8676 7524 8732
rect 7524 8676 7580 8732
rect 7580 8676 7584 8732
rect 7520 8672 7584 8676
rect 7600 8732 7664 8736
rect 7600 8676 7604 8732
rect 7604 8676 7660 8732
rect 7660 8676 7664 8732
rect 7600 8672 7664 8676
rect 7680 8732 7744 8736
rect 7680 8676 7684 8732
rect 7684 8676 7740 8732
rect 7740 8676 7744 8732
rect 7680 8672 7744 8676
rect 13360 8732 13424 8736
rect 13360 8676 13364 8732
rect 13364 8676 13420 8732
rect 13420 8676 13424 8732
rect 13360 8672 13424 8676
rect 13440 8732 13504 8736
rect 13440 8676 13444 8732
rect 13444 8676 13500 8732
rect 13500 8676 13504 8732
rect 13440 8672 13504 8676
rect 13520 8732 13584 8736
rect 13520 8676 13524 8732
rect 13524 8676 13580 8732
rect 13580 8676 13584 8732
rect 13520 8672 13584 8676
rect 13600 8732 13664 8736
rect 13600 8676 13604 8732
rect 13604 8676 13660 8732
rect 13660 8676 13664 8732
rect 13600 8672 13664 8676
rect 13680 8732 13744 8736
rect 13680 8676 13684 8732
rect 13684 8676 13740 8732
rect 13740 8676 13744 8732
rect 13680 8672 13744 8676
rect 19360 8732 19424 8736
rect 19360 8676 19364 8732
rect 19364 8676 19420 8732
rect 19420 8676 19424 8732
rect 19360 8672 19424 8676
rect 19440 8732 19504 8736
rect 19440 8676 19444 8732
rect 19444 8676 19500 8732
rect 19500 8676 19504 8732
rect 19440 8672 19504 8676
rect 19520 8732 19584 8736
rect 19520 8676 19524 8732
rect 19524 8676 19580 8732
rect 19580 8676 19584 8732
rect 19520 8672 19584 8676
rect 19600 8732 19664 8736
rect 19600 8676 19604 8732
rect 19604 8676 19660 8732
rect 19660 8676 19664 8732
rect 19600 8672 19664 8676
rect 19680 8732 19744 8736
rect 19680 8676 19684 8732
rect 19684 8676 19740 8732
rect 19740 8676 19744 8732
rect 19680 8672 19744 8676
rect 5764 8664 5828 8668
rect 5764 8608 5778 8664
rect 5778 8608 5828 8664
rect 5764 8604 5828 8608
rect 9260 8604 9324 8668
rect 18092 8604 18156 8668
rect 5396 8332 5460 8396
rect 12572 8196 12636 8260
rect 15148 8196 15212 8260
rect 4360 8188 4424 8192
rect 4360 8132 4364 8188
rect 4364 8132 4420 8188
rect 4420 8132 4424 8188
rect 4360 8128 4424 8132
rect 4440 8188 4504 8192
rect 4440 8132 4444 8188
rect 4444 8132 4500 8188
rect 4500 8132 4504 8188
rect 4440 8128 4504 8132
rect 4520 8188 4584 8192
rect 4520 8132 4524 8188
rect 4524 8132 4580 8188
rect 4580 8132 4584 8188
rect 4520 8128 4584 8132
rect 4600 8188 4664 8192
rect 4600 8132 4604 8188
rect 4604 8132 4660 8188
rect 4660 8132 4664 8188
rect 4600 8128 4664 8132
rect 4680 8188 4744 8192
rect 4680 8132 4684 8188
rect 4684 8132 4740 8188
rect 4740 8132 4744 8188
rect 4680 8128 4744 8132
rect 10360 8188 10424 8192
rect 10360 8132 10364 8188
rect 10364 8132 10420 8188
rect 10420 8132 10424 8188
rect 10360 8128 10424 8132
rect 10440 8188 10504 8192
rect 10440 8132 10444 8188
rect 10444 8132 10500 8188
rect 10500 8132 10504 8188
rect 10440 8128 10504 8132
rect 10520 8188 10584 8192
rect 10520 8132 10524 8188
rect 10524 8132 10580 8188
rect 10580 8132 10584 8188
rect 10520 8128 10584 8132
rect 10600 8188 10664 8192
rect 10600 8132 10604 8188
rect 10604 8132 10660 8188
rect 10660 8132 10664 8188
rect 10600 8128 10664 8132
rect 10680 8188 10744 8192
rect 10680 8132 10684 8188
rect 10684 8132 10740 8188
rect 10740 8132 10744 8188
rect 10680 8128 10744 8132
rect 16360 8188 16424 8192
rect 16360 8132 16364 8188
rect 16364 8132 16420 8188
rect 16420 8132 16424 8188
rect 16360 8128 16424 8132
rect 16440 8188 16504 8192
rect 16440 8132 16444 8188
rect 16444 8132 16500 8188
rect 16500 8132 16504 8188
rect 16440 8128 16504 8132
rect 16520 8188 16584 8192
rect 16520 8132 16524 8188
rect 16524 8132 16580 8188
rect 16580 8132 16584 8188
rect 16520 8128 16584 8132
rect 16600 8188 16664 8192
rect 16600 8132 16604 8188
rect 16604 8132 16660 8188
rect 16660 8132 16664 8188
rect 16600 8128 16664 8132
rect 16680 8188 16744 8192
rect 16680 8132 16684 8188
rect 16684 8132 16740 8188
rect 16740 8132 16744 8188
rect 16680 8128 16744 8132
rect 22360 8188 22424 8192
rect 22360 8132 22364 8188
rect 22364 8132 22420 8188
rect 22420 8132 22424 8188
rect 22360 8128 22424 8132
rect 22440 8188 22504 8192
rect 22440 8132 22444 8188
rect 22444 8132 22500 8188
rect 22500 8132 22504 8188
rect 22440 8128 22504 8132
rect 22520 8188 22584 8192
rect 22520 8132 22524 8188
rect 22524 8132 22580 8188
rect 22580 8132 22584 8188
rect 22520 8128 22584 8132
rect 22600 8188 22664 8192
rect 22600 8132 22604 8188
rect 22604 8132 22660 8188
rect 22660 8132 22664 8188
rect 22600 8128 22664 8132
rect 22680 8188 22744 8192
rect 22680 8132 22684 8188
rect 22684 8132 22740 8188
rect 22740 8132 22744 8188
rect 22680 8128 22744 8132
rect 3188 7984 3252 7988
rect 3188 7928 3202 7984
rect 3202 7928 3252 7984
rect 3188 7924 3252 7928
rect 9260 7924 9324 7988
rect 1360 7644 1424 7648
rect 1360 7588 1364 7644
rect 1364 7588 1420 7644
rect 1420 7588 1424 7644
rect 1360 7584 1424 7588
rect 1440 7644 1504 7648
rect 1440 7588 1444 7644
rect 1444 7588 1500 7644
rect 1500 7588 1504 7644
rect 1440 7584 1504 7588
rect 1520 7644 1584 7648
rect 1520 7588 1524 7644
rect 1524 7588 1580 7644
rect 1580 7588 1584 7644
rect 1520 7584 1584 7588
rect 1600 7644 1664 7648
rect 1600 7588 1604 7644
rect 1604 7588 1660 7644
rect 1660 7588 1664 7644
rect 1600 7584 1664 7588
rect 1680 7644 1744 7648
rect 1680 7588 1684 7644
rect 1684 7588 1740 7644
rect 1740 7588 1744 7644
rect 1680 7584 1744 7588
rect 7360 7644 7424 7648
rect 7360 7588 7364 7644
rect 7364 7588 7420 7644
rect 7420 7588 7424 7644
rect 7360 7584 7424 7588
rect 7440 7644 7504 7648
rect 7440 7588 7444 7644
rect 7444 7588 7500 7644
rect 7500 7588 7504 7644
rect 7440 7584 7504 7588
rect 7520 7644 7584 7648
rect 7520 7588 7524 7644
rect 7524 7588 7580 7644
rect 7580 7588 7584 7644
rect 7520 7584 7584 7588
rect 7600 7644 7664 7648
rect 7600 7588 7604 7644
rect 7604 7588 7660 7644
rect 7660 7588 7664 7644
rect 7600 7584 7664 7588
rect 7680 7644 7744 7648
rect 7680 7588 7684 7644
rect 7684 7588 7740 7644
rect 7740 7588 7744 7644
rect 7680 7584 7744 7588
rect 13360 7644 13424 7648
rect 13360 7588 13364 7644
rect 13364 7588 13420 7644
rect 13420 7588 13424 7644
rect 13360 7584 13424 7588
rect 13440 7644 13504 7648
rect 13440 7588 13444 7644
rect 13444 7588 13500 7644
rect 13500 7588 13504 7644
rect 13440 7584 13504 7588
rect 13520 7644 13584 7648
rect 13520 7588 13524 7644
rect 13524 7588 13580 7644
rect 13580 7588 13584 7644
rect 13520 7584 13584 7588
rect 13600 7644 13664 7648
rect 13600 7588 13604 7644
rect 13604 7588 13660 7644
rect 13660 7588 13664 7644
rect 13600 7584 13664 7588
rect 13680 7644 13744 7648
rect 13680 7588 13684 7644
rect 13684 7588 13740 7644
rect 13740 7588 13744 7644
rect 13680 7584 13744 7588
rect 19360 7644 19424 7648
rect 19360 7588 19364 7644
rect 19364 7588 19420 7644
rect 19420 7588 19424 7644
rect 19360 7584 19424 7588
rect 19440 7644 19504 7648
rect 19440 7588 19444 7644
rect 19444 7588 19500 7644
rect 19500 7588 19504 7644
rect 19440 7584 19504 7588
rect 19520 7644 19584 7648
rect 19520 7588 19524 7644
rect 19524 7588 19580 7644
rect 19580 7588 19584 7644
rect 19520 7584 19584 7588
rect 19600 7644 19664 7648
rect 19600 7588 19604 7644
rect 19604 7588 19660 7644
rect 19660 7588 19664 7644
rect 19600 7584 19664 7588
rect 19680 7644 19744 7648
rect 19680 7588 19684 7644
rect 19684 7588 19740 7644
rect 19740 7588 19744 7644
rect 19680 7584 19744 7588
rect 20300 7380 20364 7444
rect 12020 7108 12084 7172
rect 4360 7100 4424 7104
rect 4360 7044 4364 7100
rect 4364 7044 4420 7100
rect 4420 7044 4424 7100
rect 4360 7040 4424 7044
rect 4440 7100 4504 7104
rect 4440 7044 4444 7100
rect 4444 7044 4500 7100
rect 4500 7044 4504 7100
rect 4440 7040 4504 7044
rect 4520 7100 4584 7104
rect 4520 7044 4524 7100
rect 4524 7044 4580 7100
rect 4580 7044 4584 7100
rect 4520 7040 4584 7044
rect 4600 7100 4664 7104
rect 4600 7044 4604 7100
rect 4604 7044 4660 7100
rect 4660 7044 4664 7100
rect 4600 7040 4664 7044
rect 4680 7100 4744 7104
rect 4680 7044 4684 7100
rect 4684 7044 4740 7100
rect 4740 7044 4744 7100
rect 4680 7040 4744 7044
rect 10360 7100 10424 7104
rect 10360 7044 10364 7100
rect 10364 7044 10420 7100
rect 10420 7044 10424 7100
rect 10360 7040 10424 7044
rect 10440 7100 10504 7104
rect 10440 7044 10444 7100
rect 10444 7044 10500 7100
rect 10500 7044 10504 7100
rect 10440 7040 10504 7044
rect 10520 7100 10584 7104
rect 10520 7044 10524 7100
rect 10524 7044 10580 7100
rect 10580 7044 10584 7100
rect 10520 7040 10584 7044
rect 10600 7100 10664 7104
rect 10600 7044 10604 7100
rect 10604 7044 10660 7100
rect 10660 7044 10664 7100
rect 10600 7040 10664 7044
rect 10680 7100 10744 7104
rect 10680 7044 10684 7100
rect 10684 7044 10740 7100
rect 10740 7044 10744 7100
rect 10680 7040 10744 7044
rect 16360 7100 16424 7104
rect 16360 7044 16364 7100
rect 16364 7044 16420 7100
rect 16420 7044 16424 7100
rect 16360 7040 16424 7044
rect 16440 7100 16504 7104
rect 16440 7044 16444 7100
rect 16444 7044 16500 7100
rect 16500 7044 16504 7100
rect 16440 7040 16504 7044
rect 16520 7100 16584 7104
rect 16520 7044 16524 7100
rect 16524 7044 16580 7100
rect 16580 7044 16584 7100
rect 16520 7040 16584 7044
rect 16600 7100 16664 7104
rect 16600 7044 16604 7100
rect 16604 7044 16660 7100
rect 16660 7044 16664 7100
rect 16600 7040 16664 7044
rect 16680 7100 16744 7104
rect 16680 7044 16684 7100
rect 16684 7044 16740 7100
rect 16740 7044 16744 7100
rect 16680 7040 16744 7044
rect 22360 7100 22424 7104
rect 22360 7044 22364 7100
rect 22364 7044 22420 7100
rect 22420 7044 22424 7100
rect 22360 7040 22424 7044
rect 22440 7100 22504 7104
rect 22440 7044 22444 7100
rect 22444 7044 22500 7100
rect 22500 7044 22504 7100
rect 22440 7040 22504 7044
rect 22520 7100 22584 7104
rect 22520 7044 22524 7100
rect 22524 7044 22580 7100
rect 22580 7044 22584 7100
rect 22520 7040 22584 7044
rect 22600 7100 22664 7104
rect 22600 7044 22604 7100
rect 22604 7044 22660 7100
rect 22660 7044 22664 7100
rect 22600 7040 22664 7044
rect 22680 7100 22744 7104
rect 22680 7044 22684 7100
rect 22684 7044 22740 7100
rect 22740 7044 22744 7100
rect 22680 7040 22744 7044
rect 5948 6972 6012 7036
rect 6684 6972 6748 7036
rect 11100 6836 11164 6900
rect 1360 6556 1424 6560
rect 1360 6500 1364 6556
rect 1364 6500 1420 6556
rect 1420 6500 1424 6556
rect 1360 6496 1424 6500
rect 1440 6556 1504 6560
rect 1440 6500 1444 6556
rect 1444 6500 1500 6556
rect 1500 6500 1504 6556
rect 1440 6496 1504 6500
rect 1520 6556 1584 6560
rect 1520 6500 1524 6556
rect 1524 6500 1580 6556
rect 1580 6500 1584 6556
rect 1520 6496 1584 6500
rect 1600 6556 1664 6560
rect 1600 6500 1604 6556
rect 1604 6500 1660 6556
rect 1660 6500 1664 6556
rect 1600 6496 1664 6500
rect 1680 6556 1744 6560
rect 1680 6500 1684 6556
rect 1684 6500 1740 6556
rect 1740 6500 1744 6556
rect 1680 6496 1744 6500
rect 7360 6556 7424 6560
rect 7360 6500 7364 6556
rect 7364 6500 7420 6556
rect 7420 6500 7424 6556
rect 7360 6496 7424 6500
rect 7440 6556 7504 6560
rect 7440 6500 7444 6556
rect 7444 6500 7500 6556
rect 7500 6500 7504 6556
rect 7440 6496 7504 6500
rect 7520 6556 7584 6560
rect 7520 6500 7524 6556
rect 7524 6500 7580 6556
rect 7580 6500 7584 6556
rect 7520 6496 7584 6500
rect 7600 6556 7664 6560
rect 7600 6500 7604 6556
rect 7604 6500 7660 6556
rect 7660 6500 7664 6556
rect 7600 6496 7664 6500
rect 7680 6556 7744 6560
rect 7680 6500 7684 6556
rect 7684 6500 7740 6556
rect 7740 6500 7744 6556
rect 7680 6496 7744 6500
rect 13360 6556 13424 6560
rect 13360 6500 13364 6556
rect 13364 6500 13420 6556
rect 13420 6500 13424 6556
rect 13360 6496 13424 6500
rect 13440 6556 13504 6560
rect 13440 6500 13444 6556
rect 13444 6500 13500 6556
rect 13500 6500 13504 6556
rect 13440 6496 13504 6500
rect 13520 6556 13584 6560
rect 13520 6500 13524 6556
rect 13524 6500 13580 6556
rect 13580 6500 13584 6556
rect 13520 6496 13584 6500
rect 13600 6556 13664 6560
rect 13600 6500 13604 6556
rect 13604 6500 13660 6556
rect 13660 6500 13664 6556
rect 13600 6496 13664 6500
rect 13680 6556 13744 6560
rect 13680 6500 13684 6556
rect 13684 6500 13740 6556
rect 13740 6500 13744 6556
rect 13680 6496 13744 6500
rect 19360 6556 19424 6560
rect 19360 6500 19364 6556
rect 19364 6500 19420 6556
rect 19420 6500 19424 6556
rect 19360 6496 19424 6500
rect 19440 6556 19504 6560
rect 19440 6500 19444 6556
rect 19444 6500 19500 6556
rect 19500 6500 19504 6556
rect 19440 6496 19504 6500
rect 19520 6556 19584 6560
rect 19520 6500 19524 6556
rect 19524 6500 19580 6556
rect 19580 6500 19584 6556
rect 19520 6496 19584 6500
rect 19600 6556 19664 6560
rect 19600 6500 19604 6556
rect 19604 6500 19660 6556
rect 19660 6500 19664 6556
rect 19600 6496 19664 6500
rect 19680 6556 19744 6560
rect 19680 6500 19684 6556
rect 19684 6500 19740 6556
rect 19740 6500 19744 6556
rect 19680 6496 19744 6500
rect 7052 6428 7116 6492
rect 5948 6292 6012 6356
rect 19932 6292 19996 6356
rect 4360 6012 4424 6016
rect 4360 5956 4364 6012
rect 4364 5956 4420 6012
rect 4420 5956 4424 6012
rect 4360 5952 4424 5956
rect 4440 6012 4504 6016
rect 4440 5956 4444 6012
rect 4444 5956 4500 6012
rect 4500 5956 4504 6012
rect 4440 5952 4504 5956
rect 4520 6012 4584 6016
rect 4520 5956 4524 6012
rect 4524 5956 4580 6012
rect 4580 5956 4584 6012
rect 4520 5952 4584 5956
rect 4600 6012 4664 6016
rect 4600 5956 4604 6012
rect 4604 5956 4660 6012
rect 4660 5956 4664 6012
rect 4600 5952 4664 5956
rect 4680 6012 4744 6016
rect 4680 5956 4684 6012
rect 4684 5956 4740 6012
rect 4740 5956 4744 6012
rect 4680 5952 4744 5956
rect 10360 6012 10424 6016
rect 10360 5956 10364 6012
rect 10364 5956 10420 6012
rect 10420 5956 10424 6012
rect 10360 5952 10424 5956
rect 10440 6012 10504 6016
rect 10440 5956 10444 6012
rect 10444 5956 10500 6012
rect 10500 5956 10504 6012
rect 10440 5952 10504 5956
rect 10520 6012 10584 6016
rect 10520 5956 10524 6012
rect 10524 5956 10580 6012
rect 10580 5956 10584 6012
rect 10520 5952 10584 5956
rect 10600 6012 10664 6016
rect 10600 5956 10604 6012
rect 10604 5956 10660 6012
rect 10660 5956 10664 6012
rect 10600 5952 10664 5956
rect 10680 6012 10744 6016
rect 10680 5956 10684 6012
rect 10684 5956 10740 6012
rect 10740 5956 10744 6012
rect 10680 5952 10744 5956
rect 16360 6012 16424 6016
rect 16360 5956 16364 6012
rect 16364 5956 16420 6012
rect 16420 5956 16424 6012
rect 16360 5952 16424 5956
rect 16440 6012 16504 6016
rect 16440 5956 16444 6012
rect 16444 5956 16500 6012
rect 16500 5956 16504 6012
rect 16440 5952 16504 5956
rect 16520 6012 16584 6016
rect 16520 5956 16524 6012
rect 16524 5956 16580 6012
rect 16580 5956 16584 6012
rect 16520 5952 16584 5956
rect 16600 6012 16664 6016
rect 16600 5956 16604 6012
rect 16604 5956 16660 6012
rect 16660 5956 16664 6012
rect 16600 5952 16664 5956
rect 16680 6012 16744 6016
rect 16680 5956 16684 6012
rect 16684 5956 16740 6012
rect 16740 5956 16744 6012
rect 16680 5952 16744 5956
rect 22360 6012 22424 6016
rect 22360 5956 22364 6012
rect 22364 5956 22420 6012
rect 22420 5956 22424 6012
rect 22360 5952 22424 5956
rect 22440 6012 22504 6016
rect 22440 5956 22444 6012
rect 22444 5956 22500 6012
rect 22500 5956 22504 6012
rect 22440 5952 22504 5956
rect 22520 6012 22584 6016
rect 22520 5956 22524 6012
rect 22524 5956 22580 6012
rect 22580 5956 22584 6012
rect 22520 5952 22584 5956
rect 22600 6012 22664 6016
rect 22600 5956 22604 6012
rect 22604 5956 22660 6012
rect 22660 5956 22664 6012
rect 22600 5952 22664 5956
rect 22680 6012 22744 6016
rect 22680 5956 22684 6012
rect 22684 5956 22740 6012
rect 22740 5956 22744 6012
rect 22680 5952 22744 5956
rect 10180 5884 10244 5948
rect 15700 5748 15764 5812
rect 20852 5612 20916 5676
rect 7972 5476 8036 5540
rect 10916 5476 10980 5540
rect 1360 5468 1424 5472
rect 1360 5412 1364 5468
rect 1364 5412 1420 5468
rect 1420 5412 1424 5468
rect 1360 5408 1424 5412
rect 1440 5468 1504 5472
rect 1440 5412 1444 5468
rect 1444 5412 1500 5468
rect 1500 5412 1504 5468
rect 1440 5408 1504 5412
rect 1520 5468 1584 5472
rect 1520 5412 1524 5468
rect 1524 5412 1580 5468
rect 1580 5412 1584 5468
rect 1520 5408 1584 5412
rect 1600 5468 1664 5472
rect 1600 5412 1604 5468
rect 1604 5412 1660 5468
rect 1660 5412 1664 5468
rect 1600 5408 1664 5412
rect 1680 5468 1744 5472
rect 1680 5412 1684 5468
rect 1684 5412 1740 5468
rect 1740 5412 1744 5468
rect 1680 5408 1744 5412
rect 7360 5468 7424 5472
rect 7360 5412 7364 5468
rect 7364 5412 7420 5468
rect 7420 5412 7424 5468
rect 7360 5408 7424 5412
rect 7440 5468 7504 5472
rect 7440 5412 7444 5468
rect 7444 5412 7500 5468
rect 7500 5412 7504 5468
rect 7440 5408 7504 5412
rect 7520 5468 7584 5472
rect 7520 5412 7524 5468
rect 7524 5412 7580 5468
rect 7580 5412 7584 5468
rect 7520 5408 7584 5412
rect 7600 5468 7664 5472
rect 7600 5412 7604 5468
rect 7604 5412 7660 5468
rect 7660 5412 7664 5468
rect 7600 5408 7664 5412
rect 7680 5468 7744 5472
rect 7680 5412 7684 5468
rect 7684 5412 7740 5468
rect 7740 5412 7744 5468
rect 7680 5408 7744 5412
rect 13360 5468 13424 5472
rect 13360 5412 13364 5468
rect 13364 5412 13420 5468
rect 13420 5412 13424 5468
rect 13360 5408 13424 5412
rect 13440 5468 13504 5472
rect 13440 5412 13444 5468
rect 13444 5412 13500 5468
rect 13500 5412 13504 5468
rect 13440 5408 13504 5412
rect 13520 5468 13584 5472
rect 13520 5412 13524 5468
rect 13524 5412 13580 5468
rect 13580 5412 13584 5468
rect 13520 5408 13584 5412
rect 13600 5468 13664 5472
rect 13600 5412 13604 5468
rect 13604 5412 13660 5468
rect 13660 5412 13664 5468
rect 13600 5408 13664 5412
rect 13680 5468 13744 5472
rect 13680 5412 13684 5468
rect 13684 5412 13740 5468
rect 13740 5412 13744 5468
rect 13680 5408 13744 5412
rect 19360 5468 19424 5472
rect 19360 5412 19364 5468
rect 19364 5412 19420 5468
rect 19420 5412 19424 5468
rect 19360 5408 19424 5412
rect 19440 5468 19504 5472
rect 19440 5412 19444 5468
rect 19444 5412 19500 5468
rect 19500 5412 19504 5468
rect 19440 5408 19504 5412
rect 19520 5468 19584 5472
rect 19520 5412 19524 5468
rect 19524 5412 19580 5468
rect 19580 5412 19584 5468
rect 19520 5408 19584 5412
rect 19600 5468 19664 5472
rect 19600 5412 19604 5468
rect 19604 5412 19660 5468
rect 19660 5412 19664 5468
rect 19600 5408 19664 5412
rect 19680 5468 19744 5472
rect 19680 5412 19684 5468
rect 19684 5412 19740 5468
rect 19740 5412 19744 5468
rect 19680 5408 19744 5412
rect 9628 5204 9692 5268
rect 15148 5204 15212 5268
rect 19012 5204 19076 5268
rect 3740 4720 3804 4724
rect 3740 4664 3754 4720
rect 3754 4664 3804 4720
rect 3740 4660 3804 4664
rect 4360 4924 4424 4928
rect 4360 4868 4364 4924
rect 4364 4868 4420 4924
rect 4420 4868 4424 4924
rect 4360 4864 4424 4868
rect 4440 4924 4504 4928
rect 4440 4868 4444 4924
rect 4444 4868 4500 4924
rect 4500 4868 4504 4924
rect 4440 4864 4504 4868
rect 4520 4924 4584 4928
rect 4520 4868 4524 4924
rect 4524 4868 4580 4924
rect 4580 4868 4584 4924
rect 4520 4864 4584 4868
rect 4600 4924 4664 4928
rect 4600 4868 4604 4924
rect 4604 4868 4660 4924
rect 4660 4868 4664 4924
rect 4600 4864 4664 4868
rect 4680 4924 4744 4928
rect 4680 4868 4684 4924
rect 4684 4868 4740 4924
rect 4740 4868 4744 4924
rect 4680 4864 4744 4868
rect 10360 4924 10424 4928
rect 10360 4868 10364 4924
rect 10364 4868 10420 4924
rect 10420 4868 10424 4924
rect 10360 4864 10424 4868
rect 10440 4924 10504 4928
rect 10440 4868 10444 4924
rect 10444 4868 10500 4924
rect 10500 4868 10504 4924
rect 10440 4864 10504 4868
rect 10520 4924 10584 4928
rect 10520 4868 10524 4924
rect 10524 4868 10580 4924
rect 10580 4868 10584 4924
rect 10520 4864 10584 4868
rect 10600 4924 10664 4928
rect 10600 4868 10604 4924
rect 10604 4868 10660 4924
rect 10660 4868 10664 4924
rect 10600 4864 10664 4868
rect 10680 4924 10744 4928
rect 10680 4868 10684 4924
rect 10684 4868 10740 4924
rect 10740 4868 10744 4924
rect 10680 4864 10744 4868
rect 16360 4924 16424 4928
rect 16360 4868 16364 4924
rect 16364 4868 16420 4924
rect 16420 4868 16424 4924
rect 16360 4864 16424 4868
rect 16440 4924 16504 4928
rect 16440 4868 16444 4924
rect 16444 4868 16500 4924
rect 16500 4868 16504 4924
rect 16440 4864 16504 4868
rect 16520 4924 16584 4928
rect 16520 4868 16524 4924
rect 16524 4868 16580 4924
rect 16580 4868 16584 4924
rect 16520 4864 16584 4868
rect 16600 4924 16664 4928
rect 16600 4868 16604 4924
rect 16604 4868 16660 4924
rect 16660 4868 16664 4924
rect 16600 4864 16664 4868
rect 16680 4924 16744 4928
rect 16680 4868 16684 4924
rect 16684 4868 16740 4924
rect 16740 4868 16744 4924
rect 16680 4864 16744 4868
rect 22360 4924 22424 4928
rect 22360 4868 22364 4924
rect 22364 4868 22420 4924
rect 22420 4868 22424 4924
rect 22360 4864 22424 4868
rect 22440 4924 22504 4928
rect 22440 4868 22444 4924
rect 22444 4868 22500 4924
rect 22500 4868 22504 4924
rect 22440 4864 22504 4868
rect 22520 4924 22584 4928
rect 22520 4868 22524 4924
rect 22524 4868 22580 4924
rect 22580 4868 22584 4924
rect 22520 4864 22584 4868
rect 22600 4924 22664 4928
rect 22600 4868 22604 4924
rect 22604 4868 22660 4924
rect 22660 4868 22664 4924
rect 22600 4864 22664 4868
rect 22680 4924 22744 4928
rect 22680 4868 22684 4924
rect 22684 4868 22740 4924
rect 22740 4868 22744 4924
rect 22680 4864 22744 4868
rect 1360 4380 1424 4384
rect 1360 4324 1364 4380
rect 1364 4324 1420 4380
rect 1420 4324 1424 4380
rect 1360 4320 1424 4324
rect 1440 4380 1504 4384
rect 1440 4324 1444 4380
rect 1444 4324 1500 4380
rect 1500 4324 1504 4380
rect 1440 4320 1504 4324
rect 1520 4380 1584 4384
rect 1520 4324 1524 4380
rect 1524 4324 1580 4380
rect 1580 4324 1584 4380
rect 1520 4320 1584 4324
rect 1600 4380 1664 4384
rect 1600 4324 1604 4380
rect 1604 4324 1660 4380
rect 1660 4324 1664 4380
rect 1600 4320 1664 4324
rect 1680 4380 1744 4384
rect 1680 4324 1684 4380
rect 1684 4324 1740 4380
rect 1740 4324 1744 4380
rect 1680 4320 1744 4324
rect 7360 4380 7424 4384
rect 7360 4324 7364 4380
rect 7364 4324 7420 4380
rect 7420 4324 7424 4380
rect 7360 4320 7424 4324
rect 7440 4380 7504 4384
rect 7440 4324 7444 4380
rect 7444 4324 7500 4380
rect 7500 4324 7504 4380
rect 7440 4320 7504 4324
rect 7520 4380 7584 4384
rect 7520 4324 7524 4380
rect 7524 4324 7580 4380
rect 7580 4324 7584 4380
rect 7520 4320 7584 4324
rect 7600 4380 7664 4384
rect 7600 4324 7604 4380
rect 7604 4324 7660 4380
rect 7660 4324 7664 4380
rect 7600 4320 7664 4324
rect 7680 4380 7744 4384
rect 7680 4324 7684 4380
rect 7684 4324 7740 4380
rect 7740 4324 7744 4380
rect 7680 4320 7744 4324
rect 13360 4380 13424 4384
rect 13360 4324 13364 4380
rect 13364 4324 13420 4380
rect 13420 4324 13424 4380
rect 13360 4320 13424 4324
rect 13440 4380 13504 4384
rect 13440 4324 13444 4380
rect 13444 4324 13500 4380
rect 13500 4324 13504 4380
rect 13440 4320 13504 4324
rect 13520 4380 13584 4384
rect 13520 4324 13524 4380
rect 13524 4324 13580 4380
rect 13580 4324 13584 4380
rect 13520 4320 13584 4324
rect 13600 4380 13664 4384
rect 13600 4324 13604 4380
rect 13604 4324 13660 4380
rect 13660 4324 13664 4380
rect 13600 4320 13664 4324
rect 13680 4380 13744 4384
rect 13680 4324 13684 4380
rect 13684 4324 13740 4380
rect 13740 4324 13744 4380
rect 13680 4320 13744 4324
rect 19360 4380 19424 4384
rect 19360 4324 19364 4380
rect 19364 4324 19420 4380
rect 19420 4324 19424 4380
rect 19360 4320 19424 4324
rect 19440 4380 19504 4384
rect 19440 4324 19444 4380
rect 19444 4324 19500 4380
rect 19500 4324 19504 4380
rect 19440 4320 19504 4324
rect 19520 4380 19584 4384
rect 19520 4324 19524 4380
rect 19524 4324 19580 4380
rect 19580 4324 19584 4380
rect 19520 4320 19584 4324
rect 19600 4380 19664 4384
rect 19600 4324 19604 4380
rect 19604 4324 19660 4380
rect 19660 4324 19664 4380
rect 19600 4320 19664 4324
rect 19680 4380 19744 4384
rect 19680 4324 19684 4380
rect 19684 4324 19740 4380
rect 19740 4324 19744 4380
rect 19680 4320 19744 4324
rect 9996 4116 10060 4180
rect 21588 4116 21652 4180
rect 3924 3980 3988 4044
rect 21036 3980 21100 4044
rect 4360 3836 4424 3840
rect 4360 3780 4364 3836
rect 4364 3780 4420 3836
rect 4420 3780 4424 3836
rect 4360 3776 4424 3780
rect 4440 3836 4504 3840
rect 4440 3780 4444 3836
rect 4444 3780 4500 3836
rect 4500 3780 4504 3836
rect 4440 3776 4504 3780
rect 4520 3836 4584 3840
rect 4520 3780 4524 3836
rect 4524 3780 4580 3836
rect 4580 3780 4584 3836
rect 4520 3776 4584 3780
rect 4600 3836 4664 3840
rect 4600 3780 4604 3836
rect 4604 3780 4660 3836
rect 4660 3780 4664 3836
rect 4600 3776 4664 3780
rect 4680 3836 4744 3840
rect 4680 3780 4684 3836
rect 4684 3780 4740 3836
rect 4740 3780 4744 3836
rect 4680 3776 4744 3780
rect 10360 3836 10424 3840
rect 10360 3780 10364 3836
rect 10364 3780 10420 3836
rect 10420 3780 10424 3836
rect 10360 3776 10424 3780
rect 10440 3836 10504 3840
rect 10440 3780 10444 3836
rect 10444 3780 10500 3836
rect 10500 3780 10504 3836
rect 10440 3776 10504 3780
rect 10520 3836 10584 3840
rect 10520 3780 10524 3836
rect 10524 3780 10580 3836
rect 10580 3780 10584 3836
rect 10520 3776 10584 3780
rect 10600 3836 10664 3840
rect 10600 3780 10604 3836
rect 10604 3780 10660 3836
rect 10660 3780 10664 3836
rect 10600 3776 10664 3780
rect 10680 3836 10744 3840
rect 10680 3780 10684 3836
rect 10684 3780 10740 3836
rect 10740 3780 10744 3836
rect 10680 3776 10744 3780
rect 16360 3836 16424 3840
rect 16360 3780 16364 3836
rect 16364 3780 16420 3836
rect 16420 3780 16424 3836
rect 16360 3776 16424 3780
rect 16440 3836 16504 3840
rect 16440 3780 16444 3836
rect 16444 3780 16500 3836
rect 16500 3780 16504 3836
rect 16440 3776 16504 3780
rect 16520 3836 16584 3840
rect 16520 3780 16524 3836
rect 16524 3780 16580 3836
rect 16580 3780 16584 3836
rect 16520 3776 16584 3780
rect 16600 3836 16664 3840
rect 16600 3780 16604 3836
rect 16604 3780 16660 3836
rect 16660 3780 16664 3836
rect 16600 3776 16664 3780
rect 16680 3836 16744 3840
rect 16680 3780 16684 3836
rect 16684 3780 16740 3836
rect 16740 3780 16744 3836
rect 16680 3776 16744 3780
rect 22360 3836 22424 3840
rect 22360 3780 22364 3836
rect 22364 3780 22420 3836
rect 22420 3780 22424 3836
rect 22360 3776 22424 3780
rect 22440 3836 22504 3840
rect 22440 3780 22444 3836
rect 22444 3780 22500 3836
rect 22500 3780 22504 3836
rect 22440 3776 22504 3780
rect 22520 3836 22584 3840
rect 22520 3780 22524 3836
rect 22524 3780 22580 3836
rect 22580 3780 22584 3836
rect 22520 3776 22584 3780
rect 22600 3836 22664 3840
rect 22600 3780 22604 3836
rect 22604 3780 22660 3836
rect 22660 3780 22664 3836
rect 22600 3776 22664 3780
rect 22680 3836 22744 3840
rect 22680 3780 22684 3836
rect 22684 3780 22740 3836
rect 22740 3780 22744 3836
rect 22680 3776 22744 3780
rect 20116 3572 20180 3636
rect 21036 3632 21100 3636
rect 21036 3576 21086 3632
rect 21086 3576 21100 3632
rect 21036 3572 21100 3576
rect 11284 3436 11348 3500
rect 1360 3292 1424 3296
rect 1360 3236 1364 3292
rect 1364 3236 1420 3292
rect 1420 3236 1424 3292
rect 1360 3232 1424 3236
rect 1440 3292 1504 3296
rect 1440 3236 1444 3292
rect 1444 3236 1500 3292
rect 1500 3236 1504 3292
rect 1440 3232 1504 3236
rect 1520 3292 1584 3296
rect 1520 3236 1524 3292
rect 1524 3236 1580 3292
rect 1580 3236 1584 3292
rect 1520 3232 1584 3236
rect 1600 3292 1664 3296
rect 1600 3236 1604 3292
rect 1604 3236 1660 3292
rect 1660 3236 1664 3292
rect 1600 3232 1664 3236
rect 1680 3292 1744 3296
rect 1680 3236 1684 3292
rect 1684 3236 1740 3292
rect 1740 3236 1744 3292
rect 1680 3232 1744 3236
rect 7360 3292 7424 3296
rect 7360 3236 7364 3292
rect 7364 3236 7420 3292
rect 7420 3236 7424 3292
rect 7360 3232 7424 3236
rect 7440 3292 7504 3296
rect 7440 3236 7444 3292
rect 7444 3236 7500 3292
rect 7500 3236 7504 3292
rect 7440 3232 7504 3236
rect 7520 3292 7584 3296
rect 7520 3236 7524 3292
rect 7524 3236 7580 3292
rect 7580 3236 7584 3292
rect 7520 3232 7584 3236
rect 7600 3292 7664 3296
rect 7600 3236 7604 3292
rect 7604 3236 7660 3292
rect 7660 3236 7664 3292
rect 7600 3232 7664 3236
rect 7680 3292 7744 3296
rect 7680 3236 7684 3292
rect 7684 3236 7740 3292
rect 7740 3236 7744 3292
rect 7680 3232 7744 3236
rect 13360 3292 13424 3296
rect 13360 3236 13364 3292
rect 13364 3236 13420 3292
rect 13420 3236 13424 3292
rect 13360 3232 13424 3236
rect 13440 3292 13504 3296
rect 13440 3236 13444 3292
rect 13444 3236 13500 3292
rect 13500 3236 13504 3292
rect 13440 3232 13504 3236
rect 13520 3292 13584 3296
rect 13520 3236 13524 3292
rect 13524 3236 13580 3292
rect 13580 3236 13584 3292
rect 13520 3232 13584 3236
rect 13600 3292 13664 3296
rect 13600 3236 13604 3292
rect 13604 3236 13660 3292
rect 13660 3236 13664 3292
rect 13600 3232 13664 3236
rect 13680 3292 13744 3296
rect 13680 3236 13684 3292
rect 13684 3236 13740 3292
rect 13740 3236 13744 3292
rect 13680 3232 13744 3236
rect 19360 3292 19424 3296
rect 19360 3236 19364 3292
rect 19364 3236 19420 3292
rect 19420 3236 19424 3292
rect 19360 3232 19424 3236
rect 19440 3292 19504 3296
rect 19440 3236 19444 3292
rect 19444 3236 19500 3292
rect 19500 3236 19504 3292
rect 19440 3232 19504 3236
rect 19520 3292 19584 3296
rect 19520 3236 19524 3292
rect 19524 3236 19580 3292
rect 19580 3236 19584 3292
rect 19520 3232 19584 3236
rect 19600 3292 19664 3296
rect 19600 3236 19604 3292
rect 19604 3236 19660 3292
rect 19660 3236 19664 3292
rect 19600 3232 19664 3236
rect 19680 3292 19744 3296
rect 19680 3236 19684 3292
rect 19684 3236 19740 3292
rect 19740 3236 19744 3292
rect 19680 3232 19744 3236
rect 5028 3088 5092 3092
rect 5028 3032 5042 3088
rect 5042 3032 5092 3088
rect 5028 3028 5092 3032
rect 11100 3028 11164 3092
rect 10916 2816 10980 2820
rect 10916 2760 10966 2816
rect 10966 2760 10980 2816
rect 10916 2756 10980 2760
rect 4360 2748 4424 2752
rect 4360 2692 4364 2748
rect 4364 2692 4420 2748
rect 4420 2692 4424 2748
rect 4360 2688 4424 2692
rect 4440 2748 4504 2752
rect 4440 2692 4444 2748
rect 4444 2692 4500 2748
rect 4500 2692 4504 2748
rect 4440 2688 4504 2692
rect 4520 2748 4584 2752
rect 4520 2692 4524 2748
rect 4524 2692 4580 2748
rect 4580 2692 4584 2748
rect 4520 2688 4584 2692
rect 4600 2748 4664 2752
rect 4600 2692 4604 2748
rect 4604 2692 4660 2748
rect 4660 2692 4664 2748
rect 4600 2688 4664 2692
rect 4680 2748 4744 2752
rect 4680 2692 4684 2748
rect 4684 2692 4740 2748
rect 4740 2692 4744 2748
rect 4680 2688 4744 2692
rect 10360 2748 10424 2752
rect 10360 2692 10364 2748
rect 10364 2692 10420 2748
rect 10420 2692 10424 2748
rect 10360 2688 10424 2692
rect 10440 2748 10504 2752
rect 10440 2692 10444 2748
rect 10444 2692 10500 2748
rect 10500 2692 10504 2748
rect 10440 2688 10504 2692
rect 10520 2748 10584 2752
rect 10520 2692 10524 2748
rect 10524 2692 10580 2748
rect 10580 2692 10584 2748
rect 10520 2688 10584 2692
rect 10600 2748 10664 2752
rect 10600 2692 10604 2748
rect 10604 2692 10660 2748
rect 10660 2692 10664 2748
rect 10600 2688 10664 2692
rect 10680 2748 10744 2752
rect 10680 2692 10684 2748
rect 10684 2692 10740 2748
rect 10740 2692 10744 2748
rect 10680 2688 10744 2692
rect 16360 2748 16424 2752
rect 16360 2692 16364 2748
rect 16364 2692 16420 2748
rect 16420 2692 16424 2748
rect 16360 2688 16424 2692
rect 16440 2748 16504 2752
rect 16440 2692 16444 2748
rect 16444 2692 16500 2748
rect 16500 2692 16504 2748
rect 16440 2688 16504 2692
rect 16520 2748 16584 2752
rect 16520 2692 16524 2748
rect 16524 2692 16580 2748
rect 16580 2692 16584 2748
rect 16520 2688 16584 2692
rect 16600 2748 16664 2752
rect 16600 2692 16604 2748
rect 16604 2692 16660 2748
rect 16660 2692 16664 2748
rect 16600 2688 16664 2692
rect 16680 2748 16744 2752
rect 16680 2692 16684 2748
rect 16684 2692 16740 2748
rect 16740 2692 16744 2748
rect 16680 2688 16744 2692
rect 22360 2748 22424 2752
rect 22360 2692 22364 2748
rect 22364 2692 22420 2748
rect 22420 2692 22424 2748
rect 22360 2688 22424 2692
rect 22440 2748 22504 2752
rect 22440 2692 22444 2748
rect 22444 2692 22500 2748
rect 22500 2692 22504 2748
rect 22440 2688 22504 2692
rect 22520 2748 22584 2752
rect 22520 2692 22524 2748
rect 22524 2692 22580 2748
rect 22580 2692 22584 2748
rect 22520 2688 22584 2692
rect 22600 2748 22664 2752
rect 22600 2692 22604 2748
rect 22604 2692 22660 2748
rect 22660 2692 22664 2748
rect 22600 2688 22664 2692
rect 22680 2748 22744 2752
rect 22680 2692 22684 2748
rect 22684 2692 22740 2748
rect 22740 2692 22744 2748
rect 22680 2688 22744 2692
rect 9444 2348 9508 2412
rect 10180 2408 10244 2412
rect 10180 2352 10230 2408
rect 10230 2352 10244 2408
rect 10180 2348 10244 2352
rect 1360 2204 1424 2208
rect 1360 2148 1364 2204
rect 1364 2148 1420 2204
rect 1420 2148 1424 2204
rect 1360 2144 1424 2148
rect 1440 2204 1504 2208
rect 1440 2148 1444 2204
rect 1444 2148 1500 2204
rect 1500 2148 1504 2204
rect 1440 2144 1504 2148
rect 1520 2204 1584 2208
rect 1520 2148 1524 2204
rect 1524 2148 1580 2204
rect 1580 2148 1584 2204
rect 1520 2144 1584 2148
rect 1600 2204 1664 2208
rect 1600 2148 1604 2204
rect 1604 2148 1660 2204
rect 1660 2148 1664 2204
rect 1600 2144 1664 2148
rect 1680 2204 1744 2208
rect 1680 2148 1684 2204
rect 1684 2148 1740 2204
rect 1740 2148 1744 2204
rect 1680 2144 1744 2148
rect 7360 2204 7424 2208
rect 7360 2148 7364 2204
rect 7364 2148 7420 2204
rect 7420 2148 7424 2204
rect 7360 2144 7424 2148
rect 7440 2204 7504 2208
rect 7440 2148 7444 2204
rect 7444 2148 7500 2204
rect 7500 2148 7504 2204
rect 7440 2144 7504 2148
rect 7520 2204 7584 2208
rect 7520 2148 7524 2204
rect 7524 2148 7580 2204
rect 7580 2148 7584 2204
rect 7520 2144 7584 2148
rect 7600 2204 7664 2208
rect 7600 2148 7604 2204
rect 7604 2148 7660 2204
rect 7660 2148 7664 2204
rect 7600 2144 7664 2148
rect 7680 2204 7744 2208
rect 7680 2148 7684 2204
rect 7684 2148 7740 2204
rect 7740 2148 7744 2204
rect 7680 2144 7744 2148
rect 13360 2204 13424 2208
rect 13360 2148 13364 2204
rect 13364 2148 13420 2204
rect 13420 2148 13424 2204
rect 13360 2144 13424 2148
rect 13440 2204 13504 2208
rect 13440 2148 13444 2204
rect 13444 2148 13500 2204
rect 13500 2148 13504 2204
rect 13440 2144 13504 2148
rect 13520 2204 13584 2208
rect 13520 2148 13524 2204
rect 13524 2148 13580 2204
rect 13580 2148 13584 2204
rect 13520 2144 13584 2148
rect 13600 2204 13664 2208
rect 13600 2148 13604 2204
rect 13604 2148 13660 2204
rect 13660 2148 13664 2204
rect 13600 2144 13664 2148
rect 13680 2204 13744 2208
rect 13680 2148 13684 2204
rect 13684 2148 13740 2204
rect 13740 2148 13744 2204
rect 13680 2144 13744 2148
rect 19360 2204 19424 2208
rect 19360 2148 19364 2204
rect 19364 2148 19420 2204
rect 19420 2148 19424 2204
rect 19360 2144 19424 2148
rect 19440 2204 19504 2208
rect 19440 2148 19444 2204
rect 19444 2148 19500 2204
rect 19500 2148 19504 2204
rect 19440 2144 19504 2148
rect 19520 2204 19584 2208
rect 19520 2148 19524 2204
rect 19524 2148 19580 2204
rect 19580 2148 19584 2204
rect 19520 2144 19584 2148
rect 19600 2204 19664 2208
rect 19600 2148 19604 2204
rect 19604 2148 19660 2204
rect 19660 2148 19664 2204
rect 19600 2144 19664 2148
rect 19680 2204 19744 2208
rect 19680 2148 19684 2204
rect 19684 2148 19740 2204
rect 19740 2148 19744 2204
rect 19680 2144 19744 2148
rect 9076 2076 9140 2140
rect 6500 1940 6564 2004
rect 18460 1940 18524 2004
rect 19932 1668 19996 1732
rect 4360 1660 4424 1664
rect 4360 1604 4364 1660
rect 4364 1604 4420 1660
rect 4420 1604 4424 1660
rect 4360 1600 4424 1604
rect 4440 1660 4504 1664
rect 4440 1604 4444 1660
rect 4444 1604 4500 1660
rect 4500 1604 4504 1660
rect 4440 1600 4504 1604
rect 4520 1660 4584 1664
rect 4520 1604 4524 1660
rect 4524 1604 4580 1660
rect 4580 1604 4584 1660
rect 4520 1600 4584 1604
rect 4600 1660 4664 1664
rect 4600 1604 4604 1660
rect 4604 1604 4660 1660
rect 4660 1604 4664 1660
rect 4600 1600 4664 1604
rect 4680 1660 4744 1664
rect 4680 1604 4684 1660
rect 4684 1604 4740 1660
rect 4740 1604 4744 1660
rect 4680 1600 4744 1604
rect 10360 1660 10424 1664
rect 10360 1604 10364 1660
rect 10364 1604 10420 1660
rect 10420 1604 10424 1660
rect 10360 1600 10424 1604
rect 10440 1660 10504 1664
rect 10440 1604 10444 1660
rect 10444 1604 10500 1660
rect 10500 1604 10504 1660
rect 10440 1600 10504 1604
rect 10520 1660 10584 1664
rect 10520 1604 10524 1660
rect 10524 1604 10580 1660
rect 10580 1604 10584 1660
rect 10520 1600 10584 1604
rect 10600 1660 10664 1664
rect 10600 1604 10604 1660
rect 10604 1604 10660 1660
rect 10660 1604 10664 1660
rect 10600 1600 10664 1604
rect 10680 1660 10744 1664
rect 10680 1604 10684 1660
rect 10684 1604 10740 1660
rect 10740 1604 10744 1660
rect 10680 1600 10744 1604
rect 16360 1660 16424 1664
rect 16360 1604 16364 1660
rect 16364 1604 16420 1660
rect 16420 1604 16424 1660
rect 16360 1600 16424 1604
rect 16440 1660 16504 1664
rect 16440 1604 16444 1660
rect 16444 1604 16500 1660
rect 16500 1604 16504 1660
rect 16440 1600 16504 1604
rect 16520 1660 16584 1664
rect 16520 1604 16524 1660
rect 16524 1604 16580 1660
rect 16580 1604 16584 1660
rect 16520 1600 16584 1604
rect 16600 1660 16664 1664
rect 16600 1604 16604 1660
rect 16604 1604 16660 1660
rect 16660 1604 16664 1660
rect 16600 1600 16664 1604
rect 16680 1660 16744 1664
rect 16680 1604 16684 1660
rect 16684 1604 16740 1660
rect 16740 1604 16744 1660
rect 16680 1600 16744 1604
rect 22360 1660 22424 1664
rect 22360 1604 22364 1660
rect 22364 1604 22420 1660
rect 22420 1604 22424 1660
rect 22360 1600 22424 1604
rect 22440 1660 22504 1664
rect 22440 1604 22444 1660
rect 22444 1604 22500 1660
rect 22500 1604 22504 1660
rect 22440 1600 22504 1604
rect 22520 1660 22584 1664
rect 22520 1604 22524 1660
rect 22524 1604 22580 1660
rect 22580 1604 22584 1660
rect 22520 1600 22584 1604
rect 22600 1660 22664 1664
rect 22600 1604 22604 1660
rect 22604 1604 22660 1660
rect 22660 1604 22664 1660
rect 22600 1600 22664 1604
rect 22680 1660 22744 1664
rect 22680 1604 22684 1660
rect 22684 1604 22740 1660
rect 22740 1604 22744 1660
rect 22680 1600 22744 1604
rect 5396 1592 5460 1596
rect 5396 1536 5446 1592
rect 5446 1536 5460 1592
rect 5396 1532 5460 1536
rect 6684 1456 6748 1460
rect 6684 1400 6734 1456
rect 6734 1400 6748 1456
rect 6684 1396 6748 1400
rect 9812 1320 9876 1324
rect 9812 1264 9862 1320
rect 9862 1264 9876 1320
rect 9812 1260 9876 1264
rect 11100 1260 11164 1324
rect 1360 1116 1424 1120
rect 1360 1060 1364 1116
rect 1364 1060 1420 1116
rect 1420 1060 1424 1116
rect 1360 1056 1424 1060
rect 1440 1116 1504 1120
rect 1440 1060 1444 1116
rect 1444 1060 1500 1116
rect 1500 1060 1504 1116
rect 1440 1056 1504 1060
rect 1520 1116 1584 1120
rect 1520 1060 1524 1116
rect 1524 1060 1580 1116
rect 1580 1060 1584 1116
rect 1520 1056 1584 1060
rect 1600 1116 1664 1120
rect 1600 1060 1604 1116
rect 1604 1060 1660 1116
rect 1660 1060 1664 1116
rect 1600 1056 1664 1060
rect 1680 1116 1744 1120
rect 1680 1060 1684 1116
rect 1684 1060 1740 1116
rect 1740 1060 1744 1116
rect 1680 1056 1744 1060
rect 7360 1116 7424 1120
rect 7360 1060 7364 1116
rect 7364 1060 7420 1116
rect 7420 1060 7424 1116
rect 7360 1056 7424 1060
rect 7440 1116 7504 1120
rect 7440 1060 7444 1116
rect 7444 1060 7500 1116
rect 7500 1060 7504 1116
rect 7440 1056 7504 1060
rect 7520 1116 7584 1120
rect 7520 1060 7524 1116
rect 7524 1060 7580 1116
rect 7580 1060 7584 1116
rect 7520 1056 7584 1060
rect 7600 1116 7664 1120
rect 7600 1060 7604 1116
rect 7604 1060 7660 1116
rect 7660 1060 7664 1116
rect 7600 1056 7664 1060
rect 7680 1116 7744 1120
rect 7680 1060 7684 1116
rect 7684 1060 7740 1116
rect 7740 1060 7744 1116
rect 7680 1056 7744 1060
rect 13360 1116 13424 1120
rect 13360 1060 13364 1116
rect 13364 1060 13420 1116
rect 13420 1060 13424 1116
rect 13360 1056 13424 1060
rect 13440 1116 13504 1120
rect 13440 1060 13444 1116
rect 13444 1060 13500 1116
rect 13500 1060 13504 1116
rect 13440 1056 13504 1060
rect 13520 1116 13584 1120
rect 13520 1060 13524 1116
rect 13524 1060 13580 1116
rect 13580 1060 13584 1116
rect 13520 1056 13584 1060
rect 13600 1116 13664 1120
rect 13600 1060 13604 1116
rect 13604 1060 13660 1116
rect 13660 1060 13664 1116
rect 13600 1056 13664 1060
rect 13680 1116 13744 1120
rect 13680 1060 13684 1116
rect 13684 1060 13740 1116
rect 13740 1060 13744 1116
rect 13680 1056 13744 1060
rect 19360 1116 19424 1120
rect 19360 1060 19364 1116
rect 19364 1060 19420 1116
rect 19420 1060 19424 1116
rect 19360 1056 19424 1060
rect 19440 1116 19504 1120
rect 19440 1060 19444 1116
rect 19444 1060 19500 1116
rect 19500 1060 19504 1116
rect 19440 1056 19504 1060
rect 19520 1116 19584 1120
rect 19520 1060 19524 1116
rect 19524 1060 19580 1116
rect 19580 1060 19584 1116
rect 19520 1056 19584 1060
rect 19600 1116 19664 1120
rect 19600 1060 19604 1116
rect 19604 1060 19660 1116
rect 19660 1060 19664 1116
rect 19600 1056 19664 1060
rect 19680 1116 19744 1120
rect 19680 1060 19684 1116
rect 19684 1060 19740 1116
rect 19740 1060 19744 1116
rect 19680 1056 19744 1060
rect 14412 988 14476 1052
rect 4360 572 4424 576
rect 4360 516 4364 572
rect 4364 516 4420 572
rect 4420 516 4424 572
rect 4360 512 4424 516
rect 4440 572 4504 576
rect 4440 516 4444 572
rect 4444 516 4500 572
rect 4500 516 4504 572
rect 4440 512 4504 516
rect 4520 572 4584 576
rect 4520 516 4524 572
rect 4524 516 4580 572
rect 4580 516 4584 572
rect 4520 512 4584 516
rect 4600 572 4664 576
rect 4600 516 4604 572
rect 4604 516 4660 572
rect 4660 516 4664 572
rect 4600 512 4664 516
rect 4680 572 4744 576
rect 4680 516 4684 572
rect 4684 516 4740 572
rect 4740 516 4744 572
rect 4680 512 4744 516
rect 10360 572 10424 576
rect 10360 516 10364 572
rect 10364 516 10420 572
rect 10420 516 10424 572
rect 10360 512 10424 516
rect 10440 572 10504 576
rect 10440 516 10444 572
rect 10444 516 10500 572
rect 10500 516 10504 572
rect 10440 512 10504 516
rect 10520 572 10584 576
rect 10520 516 10524 572
rect 10524 516 10580 572
rect 10580 516 10584 572
rect 10520 512 10584 516
rect 10600 572 10664 576
rect 10600 516 10604 572
rect 10604 516 10660 572
rect 10660 516 10664 572
rect 10600 512 10664 516
rect 10680 572 10744 576
rect 10680 516 10684 572
rect 10684 516 10740 572
rect 10740 516 10744 572
rect 10680 512 10744 516
rect 16360 572 16424 576
rect 16360 516 16364 572
rect 16364 516 16420 572
rect 16420 516 16424 572
rect 16360 512 16424 516
rect 16440 572 16504 576
rect 16440 516 16444 572
rect 16444 516 16500 572
rect 16500 516 16504 572
rect 16440 512 16504 516
rect 16520 572 16584 576
rect 16520 516 16524 572
rect 16524 516 16580 572
rect 16580 516 16584 572
rect 16520 512 16584 516
rect 16600 572 16664 576
rect 16600 516 16604 572
rect 16604 516 16660 572
rect 16660 516 16664 572
rect 16600 512 16664 516
rect 16680 572 16744 576
rect 16680 516 16684 572
rect 16684 516 16740 572
rect 16740 516 16744 572
rect 16680 512 16744 516
rect 22360 572 22424 576
rect 22360 516 22364 572
rect 22364 516 22420 572
rect 22420 516 22424 572
rect 22360 512 22424 516
rect 22440 572 22504 576
rect 22440 516 22444 572
rect 22444 516 22500 572
rect 22500 516 22504 572
rect 22440 512 22504 516
rect 22520 572 22584 576
rect 22520 516 22524 572
rect 22524 516 22580 572
rect 22580 516 22584 572
rect 22520 512 22584 516
rect 22600 572 22664 576
rect 22600 516 22604 572
rect 22604 516 22660 572
rect 22660 516 22664 572
rect 22600 512 22664 516
rect 22680 572 22744 576
rect 22680 516 22684 572
rect 22684 516 22740 572
rect 22740 516 22744 572
rect 22680 512 22744 516
rect 11100 308 11164 372
rect 19932 308 19996 372
<< metal4 >>
rect 1352 22880 1752 23440
rect 1352 22816 1360 22880
rect 1424 22816 1440 22880
rect 1504 22816 1520 22880
rect 1584 22816 1600 22880
rect 1664 22816 1680 22880
rect 1744 22816 1752 22880
rect 1352 21792 1752 22816
rect 4352 23424 4752 23440
rect 4352 23360 4360 23424
rect 4424 23360 4440 23424
rect 4504 23360 4520 23424
rect 4584 23360 4600 23424
rect 4664 23360 4680 23424
rect 4744 23360 4752 23424
rect 3187 22404 3253 22405
rect 3187 22340 3188 22404
rect 3252 22340 3253 22404
rect 3187 22339 3253 22340
rect 1352 21728 1360 21792
rect 1424 21728 1440 21792
rect 1504 21728 1520 21792
rect 1584 21728 1600 21792
rect 1664 21728 1680 21792
rect 1744 21728 1752 21792
rect 1352 20704 1752 21728
rect 1352 20640 1360 20704
rect 1424 20640 1440 20704
rect 1504 20640 1520 20704
rect 1584 20640 1600 20704
rect 1664 20640 1680 20704
rect 1744 20640 1752 20704
rect 1352 19616 1752 20640
rect 1352 19552 1360 19616
rect 1424 19552 1440 19616
rect 1504 19552 1520 19616
rect 1584 19552 1600 19616
rect 1664 19552 1680 19616
rect 1744 19552 1752 19616
rect 1352 18528 1752 19552
rect 1352 18464 1360 18528
rect 1424 18464 1440 18528
rect 1504 18464 1520 18528
rect 1584 18464 1600 18528
rect 1664 18464 1680 18528
rect 1744 18464 1752 18528
rect 1352 17440 1752 18464
rect 1352 17376 1360 17440
rect 1424 17376 1440 17440
rect 1504 17376 1520 17440
rect 1584 17376 1600 17440
rect 1664 17376 1680 17440
rect 1744 17376 1752 17440
rect 1352 16352 1752 17376
rect 1352 16288 1360 16352
rect 1424 16288 1440 16352
rect 1504 16288 1520 16352
rect 1584 16288 1600 16352
rect 1664 16288 1680 16352
rect 1744 16288 1752 16352
rect 1352 15264 1752 16288
rect 1352 15200 1360 15264
rect 1424 15200 1440 15264
rect 1504 15200 1520 15264
rect 1584 15200 1600 15264
rect 1664 15200 1680 15264
rect 1744 15200 1752 15264
rect 1352 14176 1752 15200
rect 1352 14112 1360 14176
rect 1424 14112 1440 14176
rect 1504 14112 1520 14176
rect 1584 14112 1600 14176
rect 1664 14112 1680 14176
rect 1744 14112 1752 14176
rect 1352 13088 1752 14112
rect 1352 13024 1360 13088
rect 1424 13024 1440 13088
rect 1504 13024 1520 13088
rect 1584 13024 1600 13088
rect 1664 13024 1680 13088
rect 1744 13024 1752 13088
rect 1352 12000 1752 13024
rect 1352 11936 1360 12000
rect 1424 11936 1440 12000
rect 1504 11936 1520 12000
rect 1584 11936 1600 12000
rect 1664 11936 1680 12000
rect 1744 11936 1752 12000
rect 1352 10912 1752 11936
rect 1352 10848 1360 10912
rect 1424 10848 1440 10912
rect 1504 10848 1520 10912
rect 1584 10848 1600 10912
rect 1664 10848 1680 10912
rect 1744 10848 1752 10912
rect 1352 9824 1752 10848
rect 1352 9760 1360 9824
rect 1424 9760 1440 9824
rect 1504 9760 1520 9824
rect 1584 9760 1600 9824
rect 1664 9760 1680 9824
rect 1744 9760 1752 9824
rect 1352 8736 1752 9760
rect 1352 8672 1360 8736
rect 1424 8672 1440 8736
rect 1504 8672 1520 8736
rect 1584 8672 1600 8736
rect 1664 8672 1680 8736
rect 1744 8672 1752 8736
rect 1352 7648 1752 8672
rect 3190 7989 3250 22339
rect 4352 22336 4752 23360
rect 7352 22880 7752 23440
rect 7352 22816 7360 22880
rect 7424 22816 7440 22880
rect 7504 22816 7520 22880
rect 7584 22816 7600 22880
rect 7664 22816 7680 22880
rect 7744 22816 7752 22880
rect 6499 22404 6565 22405
rect 6499 22340 6500 22404
rect 6564 22340 6565 22404
rect 6499 22339 6565 22340
rect 4352 22272 4360 22336
rect 4424 22272 4440 22336
rect 4504 22272 4520 22336
rect 4584 22272 4600 22336
rect 4664 22272 4680 22336
rect 4744 22272 4752 22336
rect 3923 22132 3989 22133
rect 3923 22068 3924 22132
rect 3988 22068 3989 22132
rect 3923 22067 3989 22068
rect 3739 15468 3805 15469
rect 3739 15404 3740 15468
rect 3804 15404 3805 15468
rect 3739 15403 3805 15404
rect 3187 7988 3253 7989
rect 3187 7924 3188 7988
rect 3252 7924 3253 7988
rect 3187 7923 3253 7924
rect 1352 7584 1360 7648
rect 1424 7584 1440 7648
rect 1504 7584 1520 7648
rect 1584 7584 1600 7648
rect 1664 7584 1680 7648
rect 1744 7584 1752 7648
rect 1352 6560 1752 7584
rect 1352 6496 1360 6560
rect 1424 6496 1440 6560
rect 1504 6496 1520 6560
rect 1584 6496 1600 6560
rect 1664 6496 1680 6560
rect 1744 6496 1752 6560
rect 1352 5472 1752 6496
rect 1352 5408 1360 5472
rect 1424 5408 1440 5472
rect 1504 5408 1520 5472
rect 1584 5408 1600 5472
rect 1664 5408 1680 5472
rect 1744 5408 1752 5472
rect 1352 4384 1752 5408
rect 3742 4725 3802 15403
rect 3739 4724 3805 4725
rect 3739 4660 3740 4724
rect 3804 4660 3805 4724
rect 3739 4659 3805 4660
rect 1352 4320 1360 4384
rect 1424 4320 1440 4384
rect 1504 4320 1520 4384
rect 1584 4320 1600 4384
rect 1664 4320 1680 4384
rect 1744 4320 1752 4384
rect 1352 3296 1752 4320
rect 3926 4045 3986 22067
rect 4352 21248 4752 22272
rect 4352 21184 4360 21248
rect 4424 21184 4440 21248
rect 4504 21184 4520 21248
rect 4584 21184 4600 21248
rect 4664 21184 4680 21248
rect 4744 21184 4752 21248
rect 4352 20160 4752 21184
rect 4352 20096 4360 20160
rect 4424 20096 4440 20160
rect 4504 20096 4520 20160
rect 4584 20096 4600 20160
rect 4664 20096 4680 20160
rect 4744 20096 4752 20160
rect 4352 19072 4752 20096
rect 4352 19008 4360 19072
rect 4424 19008 4440 19072
rect 4504 19008 4520 19072
rect 4584 19008 4600 19072
rect 4664 19008 4680 19072
rect 4744 19008 4752 19072
rect 4352 17984 4752 19008
rect 4352 17920 4360 17984
rect 4424 17920 4440 17984
rect 4504 17920 4520 17984
rect 4584 17920 4600 17984
rect 4664 17920 4680 17984
rect 4744 17920 4752 17984
rect 4352 16896 4752 17920
rect 5763 17100 5829 17101
rect 5763 17036 5764 17100
rect 5828 17036 5829 17100
rect 5763 17035 5829 17036
rect 4352 16832 4360 16896
rect 4424 16832 4440 16896
rect 4504 16832 4520 16896
rect 4584 16832 4600 16896
rect 4664 16832 4680 16896
rect 4744 16832 4752 16896
rect 4352 15808 4752 16832
rect 4352 15744 4360 15808
rect 4424 15744 4440 15808
rect 4504 15744 4520 15808
rect 4584 15744 4600 15808
rect 4664 15744 4680 15808
rect 4744 15744 4752 15808
rect 4352 14720 4752 15744
rect 4352 14656 4360 14720
rect 4424 14656 4440 14720
rect 4504 14656 4520 14720
rect 4584 14656 4600 14720
rect 4664 14656 4680 14720
rect 4744 14656 4752 14720
rect 4352 13632 4752 14656
rect 4352 13568 4360 13632
rect 4424 13568 4440 13632
rect 4504 13568 4520 13632
rect 4584 13568 4600 13632
rect 4664 13568 4680 13632
rect 4744 13568 4752 13632
rect 4352 12544 4752 13568
rect 4352 12480 4360 12544
rect 4424 12480 4440 12544
rect 4504 12480 4520 12544
rect 4584 12480 4600 12544
rect 4664 12480 4680 12544
rect 4744 12480 4752 12544
rect 4352 11456 4752 12480
rect 4352 11392 4360 11456
rect 4424 11392 4440 11456
rect 4504 11392 4520 11456
rect 4584 11392 4600 11456
rect 4664 11392 4680 11456
rect 4744 11392 4752 11456
rect 4352 10368 4752 11392
rect 5027 11116 5093 11117
rect 5027 11052 5028 11116
rect 5092 11052 5093 11116
rect 5027 11051 5093 11052
rect 4352 10304 4360 10368
rect 4424 10304 4440 10368
rect 4504 10304 4520 10368
rect 4584 10304 4600 10368
rect 4664 10304 4680 10368
rect 4744 10304 4752 10368
rect 4352 9280 4752 10304
rect 4352 9216 4360 9280
rect 4424 9216 4440 9280
rect 4504 9216 4520 9280
rect 4584 9216 4600 9280
rect 4664 9216 4680 9280
rect 4744 9216 4752 9280
rect 4352 8192 4752 9216
rect 4352 8128 4360 8192
rect 4424 8128 4440 8192
rect 4504 8128 4520 8192
rect 4584 8128 4600 8192
rect 4664 8128 4680 8192
rect 4744 8128 4752 8192
rect 4352 7104 4752 8128
rect 4352 7040 4360 7104
rect 4424 7040 4440 7104
rect 4504 7040 4520 7104
rect 4584 7040 4600 7104
rect 4664 7040 4680 7104
rect 4744 7040 4752 7104
rect 4352 6016 4752 7040
rect 4352 5952 4360 6016
rect 4424 5952 4440 6016
rect 4504 5952 4520 6016
rect 4584 5952 4600 6016
rect 4664 5952 4680 6016
rect 4744 5952 4752 6016
rect 4352 4928 4752 5952
rect 4352 4864 4360 4928
rect 4424 4864 4440 4928
rect 4504 4864 4520 4928
rect 4584 4864 4600 4928
rect 4664 4864 4680 4928
rect 4744 4864 4752 4928
rect 3923 4044 3989 4045
rect 3923 3980 3924 4044
rect 3988 3980 3989 4044
rect 3923 3979 3989 3980
rect 1352 3232 1360 3296
rect 1424 3232 1440 3296
rect 1504 3232 1520 3296
rect 1584 3232 1600 3296
rect 1664 3232 1680 3296
rect 1744 3232 1752 3296
rect 1352 2208 1752 3232
rect 1352 2144 1360 2208
rect 1424 2144 1440 2208
rect 1504 2144 1520 2208
rect 1584 2144 1600 2208
rect 1664 2144 1680 2208
rect 1744 2144 1752 2208
rect 1352 1120 1752 2144
rect 1352 1056 1360 1120
rect 1424 1056 1440 1120
rect 1504 1056 1520 1120
rect 1584 1056 1600 1120
rect 1664 1056 1680 1120
rect 1744 1056 1752 1120
rect 1352 496 1752 1056
rect 4352 3840 4752 4864
rect 4352 3776 4360 3840
rect 4424 3776 4440 3840
rect 4504 3776 4520 3840
rect 4584 3776 4600 3840
rect 4664 3776 4680 3840
rect 4744 3776 4752 3840
rect 4352 2752 4752 3776
rect 5030 3093 5090 11051
rect 5766 8669 5826 17035
rect 5947 13836 6013 13837
rect 5947 13772 5948 13836
rect 6012 13772 6013 13836
rect 5947 13771 6013 13772
rect 5763 8668 5829 8669
rect 5763 8604 5764 8668
rect 5828 8604 5829 8668
rect 5763 8603 5829 8604
rect 5395 8396 5461 8397
rect 5395 8332 5396 8396
rect 5460 8332 5461 8396
rect 5395 8331 5461 8332
rect 5027 3092 5093 3093
rect 5027 3028 5028 3092
rect 5092 3028 5093 3092
rect 5027 3027 5093 3028
rect 4352 2688 4360 2752
rect 4424 2688 4440 2752
rect 4504 2688 4520 2752
rect 4584 2688 4600 2752
rect 4664 2688 4680 2752
rect 4744 2688 4752 2752
rect 4352 1664 4752 2688
rect 4352 1600 4360 1664
rect 4424 1600 4440 1664
rect 4504 1600 4520 1664
rect 4584 1600 4600 1664
rect 4664 1600 4680 1664
rect 4744 1600 4752 1664
rect 4352 576 4752 1600
rect 5398 1597 5458 8331
rect 5950 7037 6010 13771
rect 5947 7036 6013 7037
rect 5947 6972 5948 7036
rect 6012 6972 6013 7036
rect 5947 6971 6013 6972
rect 5950 6357 6010 6971
rect 5947 6356 6013 6357
rect 5947 6292 5948 6356
rect 6012 6292 6013 6356
rect 5947 6291 6013 6292
rect 6502 2005 6562 22339
rect 7352 21792 7752 22816
rect 10352 23424 10752 23440
rect 10352 23360 10360 23424
rect 10424 23360 10440 23424
rect 10504 23360 10520 23424
rect 10584 23360 10600 23424
rect 10664 23360 10680 23424
rect 10744 23360 10752 23424
rect 9995 22540 10061 22541
rect 9995 22476 9996 22540
rect 10060 22476 10061 22540
rect 9995 22475 10061 22476
rect 9811 21860 9877 21861
rect 9811 21796 9812 21860
rect 9876 21796 9877 21860
rect 9811 21795 9877 21796
rect 7352 21728 7360 21792
rect 7424 21728 7440 21792
rect 7504 21728 7520 21792
rect 7584 21728 7600 21792
rect 7664 21728 7680 21792
rect 7744 21728 7752 21792
rect 6683 20772 6749 20773
rect 6683 20708 6684 20772
rect 6748 20708 6749 20772
rect 6683 20707 6749 20708
rect 6686 10709 6746 20707
rect 7352 20704 7752 21728
rect 7352 20640 7360 20704
rect 7424 20640 7440 20704
rect 7504 20640 7520 20704
rect 7584 20640 7600 20704
rect 7664 20640 7680 20704
rect 7744 20640 7752 20704
rect 7352 19616 7752 20640
rect 7352 19552 7360 19616
rect 7424 19552 7440 19616
rect 7504 19552 7520 19616
rect 7584 19552 7600 19616
rect 7664 19552 7680 19616
rect 7744 19552 7752 19616
rect 7352 18528 7752 19552
rect 7352 18464 7360 18528
rect 7424 18464 7440 18528
rect 7504 18464 7520 18528
rect 7584 18464 7600 18528
rect 7664 18464 7680 18528
rect 7744 18464 7752 18528
rect 7352 17440 7752 18464
rect 9443 18188 9509 18189
rect 9443 18186 9444 18188
rect 9262 18126 9444 18186
rect 7971 17916 8037 17917
rect 7971 17852 7972 17916
rect 8036 17852 8037 17916
rect 7971 17851 8037 17852
rect 7352 17376 7360 17440
rect 7424 17376 7440 17440
rect 7504 17376 7520 17440
rect 7584 17376 7600 17440
rect 7664 17376 7680 17440
rect 7744 17376 7752 17440
rect 7352 16352 7752 17376
rect 7352 16288 7360 16352
rect 7424 16288 7440 16352
rect 7504 16288 7520 16352
rect 7584 16288 7600 16352
rect 7664 16288 7680 16352
rect 7744 16288 7752 16352
rect 7352 15264 7752 16288
rect 7352 15200 7360 15264
rect 7424 15200 7440 15264
rect 7504 15200 7520 15264
rect 7584 15200 7600 15264
rect 7664 15200 7680 15264
rect 7744 15200 7752 15264
rect 7352 14176 7752 15200
rect 7352 14112 7360 14176
rect 7424 14112 7440 14176
rect 7504 14112 7520 14176
rect 7584 14112 7600 14176
rect 7664 14112 7680 14176
rect 7744 14112 7752 14176
rect 7352 13088 7752 14112
rect 7974 13565 8034 17851
rect 9075 13700 9141 13701
rect 9075 13636 9076 13700
rect 9140 13636 9141 13700
rect 9075 13635 9141 13636
rect 7971 13564 8037 13565
rect 7971 13500 7972 13564
rect 8036 13500 8037 13564
rect 7971 13499 8037 13500
rect 7352 13024 7360 13088
rect 7424 13024 7440 13088
rect 7504 13024 7520 13088
rect 7584 13024 7600 13088
rect 7664 13024 7680 13088
rect 7744 13024 7752 13088
rect 7352 12000 7752 13024
rect 7352 11936 7360 12000
rect 7424 11936 7440 12000
rect 7504 11936 7520 12000
rect 7584 11936 7600 12000
rect 7664 11936 7680 12000
rect 7744 11936 7752 12000
rect 7352 10912 7752 11936
rect 7971 10980 8037 10981
rect 7971 10916 7972 10980
rect 8036 10916 8037 10980
rect 7971 10915 8037 10916
rect 7352 10848 7360 10912
rect 7424 10848 7440 10912
rect 7504 10848 7520 10912
rect 7584 10848 7600 10912
rect 7664 10848 7680 10912
rect 7744 10848 7752 10912
rect 6683 10708 6749 10709
rect 6683 10644 6684 10708
rect 6748 10644 6749 10708
rect 6683 10643 6749 10644
rect 7352 9824 7752 10848
rect 7352 9760 7360 9824
rect 7424 9760 7440 9824
rect 7504 9760 7520 9824
rect 7584 9760 7600 9824
rect 7664 9760 7680 9824
rect 7744 9760 7752 9824
rect 7051 9212 7117 9213
rect 7051 9148 7052 9212
rect 7116 9148 7117 9212
rect 7051 9147 7117 9148
rect 6683 7036 6749 7037
rect 6683 6972 6684 7036
rect 6748 6972 6749 7036
rect 6683 6971 6749 6972
rect 6499 2004 6565 2005
rect 6499 1940 6500 2004
rect 6564 1940 6565 2004
rect 6499 1939 6565 1940
rect 5395 1596 5461 1597
rect 5395 1532 5396 1596
rect 5460 1532 5461 1596
rect 5395 1531 5461 1532
rect 6686 1461 6746 6971
rect 7054 6493 7114 9147
rect 7352 8736 7752 9760
rect 7352 8672 7360 8736
rect 7424 8672 7440 8736
rect 7504 8672 7520 8736
rect 7584 8672 7600 8736
rect 7664 8672 7680 8736
rect 7744 8672 7752 8736
rect 7352 7648 7752 8672
rect 7352 7584 7360 7648
rect 7424 7584 7440 7648
rect 7504 7584 7520 7648
rect 7584 7584 7600 7648
rect 7664 7584 7680 7648
rect 7744 7584 7752 7648
rect 7352 6560 7752 7584
rect 7352 6496 7360 6560
rect 7424 6496 7440 6560
rect 7504 6496 7520 6560
rect 7584 6496 7600 6560
rect 7664 6496 7680 6560
rect 7744 6496 7752 6560
rect 7051 6492 7117 6493
rect 7051 6428 7052 6492
rect 7116 6428 7117 6492
rect 7051 6427 7117 6428
rect 7352 5472 7752 6496
rect 7974 5541 8034 10915
rect 7971 5540 8037 5541
rect 7971 5476 7972 5540
rect 8036 5476 8037 5540
rect 7971 5475 8037 5476
rect 7352 5408 7360 5472
rect 7424 5408 7440 5472
rect 7504 5408 7520 5472
rect 7584 5408 7600 5472
rect 7664 5408 7680 5472
rect 7744 5408 7752 5472
rect 7352 4384 7752 5408
rect 7352 4320 7360 4384
rect 7424 4320 7440 4384
rect 7504 4320 7520 4384
rect 7584 4320 7600 4384
rect 7664 4320 7680 4384
rect 7744 4320 7752 4384
rect 7352 3296 7752 4320
rect 7352 3232 7360 3296
rect 7424 3232 7440 3296
rect 7504 3232 7520 3296
rect 7584 3232 7600 3296
rect 7664 3232 7680 3296
rect 7744 3232 7752 3296
rect 7352 2208 7752 3232
rect 7352 2144 7360 2208
rect 7424 2144 7440 2208
rect 7504 2144 7520 2208
rect 7584 2144 7600 2208
rect 7664 2144 7680 2208
rect 7744 2144 7752 2208
rect 6683 1460 6749 1461
rect 6683 1396 6684 1460
rect 6748 1396 6749 1460
rect 6683 1395 6749 1396
rect 4352 512 4360 576
rect 4424 512 4440 576
rect 4504 512 4520 576
rect 4584 512 4600 576
rect 4664 512 4680 576
rect 4744 512 4752 576
rect 4352 496 4752 512
rect 7352 1120 7752 2144
rect 9078 2141 9138 13635
rect 9262 12885 9322 18126
rect 9443 18124 9444 18126
rect 9508 18124 9509 18188
rect 9443 18123 9509 18124
rect 9443 17236 9509 17237
rect 9443 17172 9444 17236
rect 9508 17172 9509 17236
rect 9443 17171 9509 17172
rect 9259 12884 9325 12885
rect 9259 12820 9260 12884
rect 9324 12820 9325 12884
rect 9259 12819 9325 12820
rect 9259 8668 9325 8669
rect 9259 8604 9260 8668
rect 9324 8604 9325 8668
rect 9259 8603 9325 8604
rect 9262 7989 9322 8603
rect 9259 7988 9325 7989
rect 9259 7924 9260 7988
rect 9324 7924 9325 7988
rect 9259 7923 9325 7924
rect 9446 2413 9506 17171
rect 9627 9756 9693 9757
rect 9627 9692 9628 9756
rect 9692 9692 9693 9756
rect 9627 9691 9693 9692
rect 9630 5269 9690 9691
rect 9627 5268 9693 5269
rect 9627 5204 9628 5268
rect 9692 5204 9693 5268
rect 9627 5203 9693 5204
rect 9443 2412 9509 2413
rect 9443 2348 9444 2412
rect 9508 2348 9509 2412
rect 9443 2347 9509 2348
rect 9075 2140 9141 2141
rect 9075 2076 9076 2140
rect 9140 2076 9141 2140
rect 9075 2075 9141 2076
rect 9814 1325 9874 21795
rect 9998 4181 10058 22475
rect 10352 22336 10752 23360
rect 13352 22880 13752 23440
rect 13352 22816 13360 22880
rect 13424 22816 13440 22880
rect 13504 22816 13520 22880
rect 13584 22816 13600 22880
rect 13664 22816 13680 22880
rect 13744 22816 13752 22880
rect 11651 22676 11717 22677
rect 11651 22612 11652 22676
rect 11716 22612 11717 22676
rect 11651 22611 11717 22612
rect 10352 22272 10360 22336
rect 10424 22272 10440 22336
rect 10504 22272 10520 22336
rect 10584 22272 10600 22336
rect 10664 22272 10680 22336
rect 10744 22272 10752 22336
rect 10352 21248 10752 22272
rect 10352 21184 10360 21248
rect 10424 21184 10440 21248
rect 10504 21184 10520 21248
rect 10584 21184 10600 21248
rect 10664 21184 10680 21248
rect 10744 21184 10752 21248
rect 10352 20160 10752 21184
rect 10352 20096 10360 20160
rect 10424 20096 10440 20160
rect 10504 20096 10520 20160
rect 10584 20096 10600 20160
rect 10664 20096 10680 20160
rect 10744 20096 10752 20160
rect 10179 19140 10245 19141
rect 10179 19076 10180 19140
rect 10244 19076 10245 19140
rect 10179 19075 10245 19076
rect 10182 11661 10242 19075
rect 10352 19072 10752 20096
rect 10352 19008 10360 19072
rect 10424 19008 10440 19072
rect 10504 19008 10520 19072
rect 10584 19008 10600 19072
rect 10664 19008 10680 19072
rect 10744 19008 10752 19072
rect 10352 17984 10752 19008
rect 10352 17920 10360 17984
rect 10424 17920 10440 17984
rect 10504 17920 10520 17984
rect 10584 17920 10600 17984
rect 10664 17920 10680 17984
rect 10744 17920 10752 17984
rect 10352 16896 10752 17920
rect 10352 16832 10360 16896
rect 10424 16832 10440 16896
rect 10504 16832 10520 16896
rect 10584 16832 10600 16896
rect 10664 16832 10680 16896
rect 10744 16832 10752 16896
rect 10352 15808 10752 16832
rect 10352 15744 10360 15808
rect 10424 15744 10440 15808
rect 10504 15744 10520 15808
rect 10584 15744 10600 15808
rect 10664 15744 10680 15808
rect 10744 15744 10752 15808
rect 10352 14720 10752 15744
rect 11283 15332 11349 15333
rect 11283 15268 11284 15332
rect 11348 15268 11349 15332
rect 11283 15267 11349 15268
rect 10915 15060 10981 15061
rect 10915 14996 10916 15060
rect 10980 14996 10981 15060
rect 10915 14995 10981 14996
rect 10352 14656 10360 14720
rect 10424 14656 10440 14720
rect 10504 14656 10520 14720
rect 10584 14656 10600 14720
rect 10664 14656 10680 14720
rect 10744 14656 10752 14720
rect 10352 13632 10752 14656
rect 10352 13568 10360 13632
rect 10424 13568 10440 13632
rect 10504 13568 10520 13632
rect 10584 13568 10600 13632
rect 10664 13568 10680 13632
rect 10744 13568 10752 13632
rect 10352 12544 10752 13568
rect 10352 12480 10360 12544
rect 10424 12480 10440 12544
rect 10504 12480 10520 12544
rect 10584 12480 10600 12544
rect 10664 12480 10680 12544
rect 10744 12480 10752 12544
rect 10179 11660 10245 11661
rect 10179 11596 10180 11660
rect 10244 11596 10245 11660
rect 10179 11595 10245 11596
rect 10352 11456 10752 12480
rect 10918 12069 10978 14995
rect 10915 12068 10981 12069
rect 10915 12004 10916 12068
rect 10980 12004 10981 12068
rect 10915 12003 10981 12004
rect 11286 11797 11346 15267
rect 11654 13293 11714 22611
rect 13352 21792 13752 22816
rect 16352 23424 16752 23440
rect 16352 23360 16360 23424
rect 16424 23360 16440 23424
rect 16504 23360 16520 23424
rect 16584 23360 16600 23424
rect 16664 23360 16680 23424
rect 16744 23360 16752 23424
rect 16352 22336 16752 23360
rect 16352 22272 16360 22336
rect 16424 22272 16440 22336
rect 16504 22272 16520 22336
rect 16584 22272 16600 22336
rect 16664 22272 16680 22336
rect 16744 22272 16752 22336
rect 14411 21860 14477 21861
rect 14411 21796 14412 21860
rect 14476 21796 14477 21860
rect 14411 21795 14477 21796
rect 13352 21728 13360 21792
rect 13424 21728 13440 21792
rect 13504 21728 13520 21792
rect 13584 21728 13600 21792
rect 13664 21728 13680 21792
rect 13744 21728 13752 21792
rect 12755 20772 12821 20773
rect 12755 20708 12756 20772
rect 12820 20708 12821 20772
rect 12755 20707 12821 20708
rect 11835 17644 11901 17645
rect 11835 17580 11836 17644
rect 11900 17580 11901 17644
rect 11835 17579 11901 17580
rect 11838 14653 11898 17579
rect 11835 14652 11901 14653
rect 11835 14588 11836 14652
rect 11900 14588 11901 14652
rect 11835 14587 11901 14588
rect 12758 13429 12818 20707
rect 13352 20704 13752 21728
rect 13352 20640 13360 20704
rect 13424 20640 13440 20704
rect 13504 20640 13520 20704
rect 13584 20640 13600 20704
rect 13664 20640 13680 20704
rect 13744 20640 13752 20704
rect 13352 19616 13752 20640
rect 13352 19552 13360 19616
rect 13424 19552 13440 19616
rect 13504 19552 13520 19616
rect 13584 19552 13600 19616
rect 13664 19552 13680 19616
rect 13744 19552 13752 19616
rect 13352 18528 13752 19552
rect 13352 18464 13360 18528
rect 13424 18464 13440 18528
rect 13504 18464 13520 18528
rect 13584 18464 13600 18528
rect 13664 18464 13680 18528
rect 13744 18464 13752 18528
rect 13352 17440 13752 18464
rect 13352 17376 13360 17440
rect 13424 17376 13440 17440
rect 13504 17376 13520 17440
rect 13584 17376 13600 17440
rect 13664 17376 13680 17440
rect 13744 17376 13752 17440
rect 13352 16352 13752 17376
rect 13352 16288 13360 16352
rect 13424 16288 13440 16352
rect 13504 16288 13520 16352
rect 13584 16288 13600 16352
rect 13664 16288 13680 16352
rect 13744 16288 13752 16352
rect 13352 15264 13752 16288
rect 13352 15200 13360 15264
rect 13424 15200 13440 15264
rect 13504 15200 13520 15264
rect 13584 15200 13600 15264
rect 13664 15200 13680 15264
rect 13744 15200 13752 15264
rect 12939 14244 13005 14245
rect 12939 14180 12940 14244
rect 13004 14180 13005 14244
rect 12939 14179 13005 14180
rect 12755 13428 12821 13429
rect 12755 13364 12756 13428
rect 12820 13364 12821 13428
rect 12755 13363 12821 13364
rect 11651 13292 11717 13293
rect 11651 13228 11652 13292
rect 11716 13228 11717 13292
rect 11651 13227 11717 13228
rect 12571 12612 12637 12613
rect 12571 12548 12572 12612
rect 12636 12548 12637 12612
rect 12571 12547 12637 12548
rect 11283 11796 11349 11797
rect 11283 11732 11284 11796
rect 11348 11732 11349 11796
rect 11283 11731 11349 11732
rect 11283 11660 11349 11661
rect 11283 11596 11284 11660
rect 11348 11596 11349 11660
rect 11283 11595 11349 11596
rect 10352 11392 10360 11456
rect 10424 11392 10440 11456
rect 10504 11392 10520 11456
rect 10584 11392 10600 11456
rect 10664 11392 10680 11456
rect 10744 11392 10752 11456
rect 10352 10368 10752 11392
rect 10352 10304 10360 10368
rect 10424 10304 10440 10368
rect 10504 10304 10520 10368
rect 10584 10304 10600 10368
rect 10664 10304 10680 10368
rect 10744 10304 10752 10368
rect 10352 9280 10752 10304
rect 10352 9216 10360 9280
rect 10424 9216 10440 9280
rect 10504 9216 10520 9280
rect 10584 9216 10600 9280
rect 10664 9216 10680 9280
rect 10744 9216 10752 9280
rect 10352 8192 10752 9216
rect 10915 9212 10981 9213
rect 10915 9148 10916 9212
rect 10980 9148 10981 9212
rect 10915 9147 10981 9148
rect 10352 8128 10360 8192
rect 10424 8128 10440 8192
rect 10504 8128 10520 8192
rect 10584 8128 10600 8192
rect 10664 8128 10680 8192
rect 10744 8128 10752 8192
rect 10352 7104 10752 8128
rect 10352 7040 10360 7104
rect 10424 7040 10440 7104
rect 10504 7040 10520 7104
rect 10584 7040 10600 7104
rect 10664 7040 10680 7104
rect 10744 7040 10752 7104
rect 10352 6016 10752 7040
rect 10352 5952 10360 6016
rect 10424 5952 10440 6016
rect 10504 5952 10520 6016
rect 10584 5952 10600 6016
rect 10664 5952 10680 6016
rect 10744 5952 10752 6016
rect 10179 5948 10245 5949
rect 10179 5884 10180 5948
rect 10244 5884 10245 5948
rect 10179 5883 10245 5884
rect 9995 4180 10061 4181
rect 9995 4116 9996 4180
rect 10060 4116 10061 4180
rect 9995 4115 10061 4116
rect 10182 2413 10242 5883
rect 10352 4928 10752 5952
rect 10918 5541 10978 9147
rect 11099 6900 11165 6901
rect 11099 6836 11100 6900
rect 11164 6836 11165 6900
rect 11099 6835 11165 6836
rect 10915 5540 10981 5541
rect 10915 5476 10916 5540
rect 10980 5476 10981 5540
rect 10915 5475 10981 5476
rect 10352 4864 10360 4928
rect 10424 4864 10440 4928
rect 10504 4864 10520 4928
rect 10584 4864 10600 4928
rect 10664 4864 10680 4928
rect 10744 4864 10752 4928
rect 10352 3840 10752 4864
rect 10352 3776 10360 3840
rect 10424 3776 10440 3840
rect 10504 3776 10520 3840
rect 10584 3776 10600 3840
rect 10664 3776 10680 3840
rect 10744 3776 10752 3840
rect 10352 2752 10752 3776
rect 10918 2821 10978 5475
rect 11102 3093 11162 6835
rect 11286 3501 11346 11595
rect 12574 11525 12634 12547
rect 12942 12205 13002 14179
rect 13352 14176 13752 15200
rect 13352 14112 13360 14176
rect 13424 14112 13440 14176
rect 13504 14112 13520 14176
rect 13584 14112 13600 14176
rect 13664 14112 13680 14176
rect 13744 14112 13752 14176
rect 13123 13156 13189 13157
rect 13123 13092 13124 13156
rect 13188 13092 13189 13156
rect 13123 13091 13189 13092
rect 12939 12204 13005 12205
rect 12939 12140 12940 12204
rect 13004 12140 13005 12204
rect 12939 12139 13005 12140
rect 12571 11524 12637 11525
rect 12571 11460 12572 11524
rect 12636 11460 12637 11524
rect 12571 11459 12637 11460
rect 12019 11116 12085 11117
rect 12019 11052 12020 11116
rect 12084 11052 12085 11116
rect 12019 11051 12085 11052
rect 12022 7173 12082 11051
rect 13126 10573 13186 13091
rect 13352 13088 13752 14112
rect 13352 13024 13360 13088
rect 13424 13024 13440 13088
rect 13504 13024 13520 13088
rect 13584 13024 13600 13088
rect 13664 13024 13680 13088
rect 13744 13024 13752 13088
rect 13352 12000 13752 13024
rect 13352 11936 13360 12000
rect 13424 11936 13440 12000
rect 13504 11936 13520 12000
rect 13584 11936 13600 12000
rect 13664 11936 13680 12000
rect 13744 11936 13752 12000
rect 13352 10912 13752 11936
rect 13352 10848 13360 10912
rect 13424 10848 13440 10912
rect 13504 10848 13520 10912
rect 13584 10848 13600 10912
rect 13664 10848 13680 10912
rect 13744 10848 13752 10912
rect 12387 10572 12453 10573
rect 12387 10508 12388 10572
rect 12452 10570 12453 10572
rect 13123 10572 13189 10573
rect 12452 10510 12634 10570
rect 12452 10508 12453 10510
rect 12387 10507 12453 10508
rect 12574 8261 12634 10510
rect 13123 10508 13124 10572
rect 13188 10508 13189 10572
rect 13123 10507 13189 10508
rect 13352 9824 13752 10848
rect 13352 9760 13360 9824
rect 13424 9760 13440 9824
rect 13504 9760 13520 9824
rect 13584 9760 13600 9824
rect 13664 9760 13680 9824
rect 13744 9760 13752 9824
rect 13123 9620 13189 9621
rect 13123 9556 13124 9620
rect 13188 9556 13189 9620
rect 13123 9555 13189 9556
rect 13126 8805 13186 9555
rect 13123 8804 13189 8805
rect 13123 8740 13124 8804
rect 13188 8740 13189 8804
rect 13123 8739 13189 8740
rect 13352 8736 13752 9760
rect 13352 8672 13360 8736
rect 13424 8672 13440 8736
rect 13504 8672 13520 8736
rect 13584 8672 13600 8736
rect 13664 8672 13680 8736
rect 13744 8672 13752 8736
rect 12571 8260 12637 8261
rect 12571 8196 12572 8260
rect 12636 8196 12637 8260
rect 12571 8195 12637 8196
rect 13352 7648 13752 8672
rect 13352 7584 13360 7648
rect 13424 7584 13440 7648
rect 13504 7584 13520 7648
rect 13584 7584 13600 7648
rect 13664 7584 13680 7648
rect 13744 7584 13752 7648
rect 12019 7172 12085 7173
rect 12019 7108 12020 7172
rect 12084 7108 12085 7172
rect 12019 7107 12085 7108
rect 13352 6560 13752 7584
rect 13352 6496 13360 6560
rect 13424 6496 13440 6560
rect 13504 6496 13520 6560
rect 13584 6496 13600 6560
rect 13664 6496 13680 6560
rect 13744 6496 13752 6560
rect 13352 5472 13752 6496
rect 13352 5408 13360 5472
rect 13424 5408 13440 5472
rect 13504 5408 13520 5472
rect 13584 5408 13600 5472
rect 13664 5408 13680 5472
rect 13744 5408 13752 5472
rect 13352 4384 13752 5408
rect 13352 4320 13360 4384
rect 13424 4320 13440 4384
rect 13504 4320 13520 4384
rect 13584 4320 13600 4384
rect 13664 4320 13680 4384
rect 13744 4320 13752 4384
rect 11283 3500 11349 3501
rect 11283 3436 11284 3500
rect 11348 3436 11349 3500
rect 11283 3435 11349 3436
rect 13352 3296 13752 4320
rect 13352 3232 13360 3296
rect 13424 3232 13440 3296
rect 13504 3232 13520 3296
rect 13584 3232 13600 3296
rect 13664 3232 13680 3296
rect 13744 3232 13752 3296
rect 11099 3092 11165 3093
rect 11099 3028 11100 3092
rect 11164 3028 11165 3092
rect 11099 3027 11165 3028
rect 10915 2820 10981 2821
rect 10915 2756 10916 2820
rect 10980 2756 10981 2820
rect 10915 2755 10981 2756
rect 10352 2688 10360 2752
rect 10424 2688 10440 2752
rect 10504 2688 10520 2752
rect 10584 2688 10600 2752
rect 10664 2688 10680 2752
rect 10744 2688 10752 2752
rect 10179 2412 10245 2413
rect 10179 2348 10180 2412
rect 10244 2348 10245 2412
rect 10179 2347 10245 2348
rect 10352 1664 10752 2688
rect 10352 1600 10360 1664
rect 10424 1600 10440 1664
rect 10504 1600 10520 1664
rect 10584 1600 10600 1664
rect 10664 1600 10680 1664
rect 10744 1600 10752 1664
rect 9811 1324 9877 1325
rect 9811 1260 9812 1324
rect 9876 1260 9877 1324
rect 9811 1259 9877 1260
rect 7352 1056 7360 1120
rect 7424 1056 7440 1120
rect 7504 1056 7520 1120
rect 7584 1056 7600 1120
rect 7664 1056 7680 1120
rect 7744 1056 7752 1120
rect 7352 496 7752 1056
rect 10352 576 10752 1600
rect 13352 2208 13752 3232
rect 13352 2144 13360 2208
rect 13424 2144 13440 2208
rect 13504 2144 13520 2208
rect 13584 2144 13600 2208
rect 13664 2144 13680 2208
rect 13744 2144 13752 2208
rect 11099 1324 11165 1325
rect 11099 1260 11100 1324
rect 11164 1260 11165 1324
rect 11099 1259 11165 1260
rect 10352 512 10360 576
rect 10424 512 10440 576
rect 10504 512 10520 576
rect 10584 512 10600 576
rect 10664 512 10680 576
rect 10744 512 10752 576
rect 10352 496 10752 512
rect 11102 373 11162 1259
rect 13352 1120 13752 2144
rect 13352 1056 13360 1120
rect 13424 1056 13440 1120
rect 13504 1056 13520 1120
rect 13584 1056 13600 1120
rect 13664 1056 13680 1120
rect 13744 1056 13752 1120
rect 13352 496 13752 1056
rect 14414 1053 14474 21795
rect 16352 21248 16752 22272
rect 16352 21184 16360 21248
rect 16424 21184 16440 21248
rect 16504 21184 16520 21248
rect 16584 21184 16600 21248
rect 16664 21184 16680 21248
rect 16744 21184 16752 21248
rect 16352 20160 16752 21184
rect 16352 20096 16360 20160
rect 16424 20096 16440 20160
rect 16504 20096 16520 20160
rect 16584 20096 16600 20160
rect 16664 20096 16680 20160
rect 16744 20096 16752 20160
rect 15699 19276 15765 19277
rect 15699 19212 15700 19276
rect 15764 19212 15765 19276
rect 15699 19211 15765 19212
rect 14963 18052 15029 18053
rect 14963 17988 14964 18052
rect 15028 17988 15029 18052
rect 14963 17987 15029 17988
rect 14966 9077 15026 17987
rect 14963 9076 15029 9077
rect 14963 9012 14964 9076
rect 15028 9012 15029 9076
rect 14963 9011 15029 9012
rect 15147 8260 15213 8261
rect 15147 8196 15148 8260
rect 15212 8196 15213 8260
rect 15147 8195 15213 8196
rect 15150 5269 15210 8195
rect 15702 5813 15762 19211
rect 16352 19072 16752 20096
rect 19352 22880 19752 23440
rect 22352 23424 22752 23440
rect 22352 23360 22360 23424
rect 22424 23360 22440 23424
rect 22504 23360 22520 23424
rect 22584 23360 22600 23424
rect 22664 23360 22680 23424
rect 22744 23360 22752 23424
rect 21587 22948 21653 22949
rect 21587 22884 21588 22948
rect 21652 22884 21653 22948
rect 21587 22883 21653 22884
rect 19352 22816 19360 22880
rect 19424 22816 19440 22880
rect 19504 22816 19520 22880
rect 19584 22816 19600 22880
rect 19664 22816 19680 22880
rect 19744 22816 19752 22880
rect 19352 21792 19752 22816
rect 21219 22268 21285 22269
rect 21219 22204 21220 22268
rect 21284 22204 21285 22268
rect 21219 22203 21285 22204
rect 19352 21728 19360 21792
rect 19424 21728 19440 21792
rect 19504 21728 19520 21792
rect 19584 21728 19600 21792
rect 19664 21728 19680 21792
rect 19744 21728 19752 21792
rect 19352 20704 19752 21728
rect 21035 20908 21101 20909
rect 21035 20844 21036 20908
rect 21100 20844 21101 20908
rect 21035 20843 21101 20844
rect 19352 20640 19360 20704
rect 19424 20640 19440 20704
rect 19504 20640 19520 20704
rect 19584 20640 19600 20704
rect 19664 20640 19680 20704
rect 19744 20640 19752 20704
rect 18827 19684 18893 19685
rect 18827 19620 18828 19684
rect 18892 19620 18893 19684
rect 18827 19619 18893 19620
rect 16352 19008 16360 19072
rect 16424 19008 16440 19072
rect 16504 19008 16520 19072
rect 16584 19008 16600 19072
rect 16664 19008 16680 19072
rect 16744 19008 16752 19072
rect 16352 17984 16752 19008
rect 16352 17920 16360 17984
rect 16424 17920 16440 17984
rect 16504 17920 16520 17984
rect 16584 17920 16600 17984
rect 16664 17920 16680 17984
rect 16744 17920 16752 17984
rect 16352 16896 16752 17920
rect 16352 16832 16360 16896
rect 16424 16832 16440 16896
rect 16504 16832 16520 16896
rect 16584 16832 16600 16896
rect 16664 16832 16680 16896
rect 16744 16832 16752 16896
rect 16352 15808 16752 16832
rect 16352 15744 16360 15808
rect 16424 15744 16440 15808
rect 16504 15744 16520 15808
rect 16584 15744 16600 15808
rect 16664 15744 16680 15808
rect 16744 15744 16752 15808
rect 16352 14720 16752 15744
rect 18091 15604 18157 15605
rect 18091 15540 18092 15604
rect 18156 15540 18157 15604
rect 18091 15539 18157 15540
rect 16352 14656 16360 14720
rect 16424 14656 16440 14720
rect 16504 14656 16520 14720
rect 16584 14656 16600 14720
rect 16664 14656 16680 14720
rect 16744 14656 16752 14720
rect 16352 13632 16752 14656
rect 16352 13568 16360 13632
rect 16424 13568 16440 13632
rect 16504 13568 16520 13632
rect 16584 13568 16600 13632
rect 16664 13568 16680 13632
rect 16744 13568 16752 13632
rect 16352 12544 16752 13568
rect 16352 12480 16360 12544
rect 16424 12480 16440 12544
rect 16504 12480 16520 12544
rect 16584 12480 16600 12544
rect 16664 12480 16680 12544
rect 16744 12480 16752 12544
rect 16352 11456 16752 12480
rect 16352 11392 16360 11456
rect 16424 11392 16440 11456
rect 16504 11392 16520 11456
rect 16584 11392 16600 11456
rect 16664 11392 16680 11456
rect 16744 11392 16752 11456
rect 16352 10368 16752 11392
rect 16352 10304 16360 10368
rect 16424 10304 16440 10368
rect 16504 10304 16520 10368
rect 16584 10304 16600 10368
rect 16664 10304 16680 10368
rect 16744 10304 16752 10368
rect 16352 9280 16752 10304
rect 16352 9216 16360 9280
rect 16424 9216 16440 9280
rect 16504 9216 16520 9280
rect 16584 9216 16600 9280
rect 16664 9216 16680 9280
rect 16744 9216 16752 9280
rect 16352 8192 16752 9216
rect 18094 8669 18154 15539
rect 18459 13292 18525 13293
rect 18459 13228 18460 13292
rect 18524 13228 18525 13292
rect 18459 13227 18525 13228
rect 18275 9756 18341 9757
rect 18275 9692 18276 9756
rect 18340 9692 18341 9756
rect 18275 9691 18341 9692
rect 18278 8941 18338 9691
rect 18275 8940 18341 8941
rect 18275 8876 18276 8940
rect 18340 8876 18341 8940
rect 18275 8875 18341 8876
rect 18091 8668 18157 8669
rect 18091 8604 18092 8668
rect 18156 8604 18157 8668
rect 18091 8603 18157 8604
rect 16352 8128 16360 8192
rect 16424 8128 16440 8192
rect 16504 8128 16520 8192
rect 16584 8128 16600 8192
rect 16664 8128 16680 8192
rect 16744 8128 16752 8192
rect 16352 7104 16752 8128
rect 16352 7040 16360 7104
rect 16424 7040 16440 7104
rect 16504 7040 16520 7104
rect 16584 7040 16600 7104
rect 16664 7040 16680 7104
rect 16744 7040 16752 7104
rect 16352 6016 16752 7040
rect 16352 5952 16360 6016
rect 16424 5952 16440 6016
rect 16504 5952 16520 6016
rect 16584 5952 16600 6016
rect 16664 5952 16680 6016
rect 16744 5952 16752 6016
rect 15699 5812 15765 5813
rect 15699 5748 15700 5812
rect 15764 5748 15765 5812
rect 15699 5747 15765 5748
rect 15147 5268 15213 5269
rect 15147 5204 15148 5268
rect 15212 5204 15213 5268
rect 15147 5203 15213 5204
rect 16352 4928 16752 5952
rect 16352 4864 16360 4928
rect 16424 4864 16440 4928
rect 16504 4864 16520 4928
rect 16584 4864 16600 4928
rect 16664 4864 16680 4928
rect 16744 4864 16752 4928
rect 16352 3840 16752 4864
rect 16352 3776 16360 3840
rect 16424 3776 16440 3840
rect 16504 3776 16520 3840
rect 16584 3776 16600 3840
rect 16664 3776 16680 3840
rect 16744 3776 16752 3840
rect 16352 2752 16752 3776
rect 16352 2688 16360 2752
rect 16424 2688 16440 2752
rect 16504 2688 16520 2752
rect 16584 2688 16600 2752
rect 16664 2688 16680 2752
rect 16744 2688 16752 2752
rect 16352 1664 16752 2688
rect 18462 2005 18522 13227
rect 18830 10029 18890 19619
rect 19352 19616 19752 20640
rect 19352 19552 19360 19616
rect 19424 19552 19440 19616
rect 19504 19552 19520 19616
rect 19584 19552 19600 19616
rect 19664 19552 19680 19616
rect 19744 19552 19752 19616
rect 19011 19412 19077 19413
rect 19011 19348 19012 19412
rect 19076 19348 19077 19412
rect 19011 19347 19077 19348
rect 18827 10028 18893 10029
rect 18827 9964 18828 10028
rect 18892 9964 18893 10028
rect 18827 9963 18893 9964
rect 19014 5269 19074 19347
rect 19352 18528 19752 19552
rect 19931 18596 19997 18597
rect 19931 18532 19932 18596
rect 19996 18532 19997 18596
rect 19931 18531 19997 18532
rect 19352 18464 19360 18528
rect 19424 18464 19440 18528
rect 19504 18464 19520 18528
rect 19584 18464 19600 18528
rect 19664 18464 19680 18528
rect 19744 18464 19752 18528
rect 19352 17440 19752 18464
rect 19352 17376 19360 17440
rect 19424 17376 19440 17440
rect 19504 17376 19520 17440
rect 19584 17376 19600 17440
rect 19664 17376 19680 17440
rect 19744 17376 19752 17440
rect 19352 16352 19752 17376
rect 19352 16288 19360 16352
rect 19424 16288 19440 16352
rect 19504 16288 19520 16352
rect 19584 16288 19600 16352
rect 19664 16288 19680 16352
rect 19744 16288 19752 16352
rect 19352 15264 19752 16288
rect 19352 15200 19360 15264
rect 19424 15200 19440 15264
rect 19504 15200 19520 15264
rect 19584 15200 19600 15264
rect 19664 15200 19680 15264
rect 19744 15200 19752 15264
rect 19195 14516 19261 14517
rect 19195 14452 19196 14516
rect 19260 14452 19261 14516
rect 19195 14451 19261 14452
rect 19198 10709 19258 14451
rect 19352 14176 19752 15200
rect 19352 14112 19360 14176
rect 19424 14112 19440 14176
rect 19504 14112 19520 14176
rect 19584 14112 19600 14176
rect 19664 14112 19680 14176
rect 19744 14112 19752 14176
rect 19352 13088 19752 14112
rect 19352 13024 19360 13088
rect 19424 13024 19440 13088
rect 19504 13024 19520 13088
rect 19584 13024 19600 13088
rect 19664 13024 19680 13088
rect 19744 13024 19752 13088
rect 19352 12000 19752 13024
rect 19934 12450 19994 18531
rect 20667 18052 20733 18053
rect 20667 17988 20668 18052
rect 20732 17988 20733 18052
rect 20667 17987 20733 17988
rect 19934 12390 20178 12450
rect 19352 11936 19360 12000
rect 19424 11936 19440 12000
rect 19504 11936 19520 12000
rect 19584 11936 19600 12000
rect 19664 11936 19680 12000
rect 19744 11936 19752 12000
rect 19352 10912 19752 11936
rect 19352 10848 19360 10912
rect 19424 10848 19440 10912
rect 19504 10848 19520 10912
rect 19584 10848 19600 10912
rect 19664 10848 19680 10912
rect 19744 10848 19752 10912
rect 19195 10708 19261 10709
rect 19195 10644 19196 10708
rect 19260 10644 19261 10708
rect 19195 10643 19261 10644
rect 19352 9824 19752 10848
rect 19931 10028 19997 10029
rect 19931 9964 19932 10028
rect 19996 9964 19997 10028
rect 19931 9963 19997 9964
rect 19352 9760 19360 9824
rect 19424 9760 19440 9824
rect 19504 9760 19520 9824
rect 19584 9760 19600 9824
rect 19664 9760 19680 9824
rect 19744 9760 19752 9824
rect 19352 8736 19752 9760
rect 19352 8672 19360 8736
rect 19424 8672 19440 8736
rect 19504 8672 19520 8736
rect 19584 8672 19600 8736
rect 19664 8672 19680 8736
rect 19744 8672 19752 8736
rect 19352 7648 19752 8672
rect 19352 7584 19360 7648
rect 19424 7584 19440 7648
rect 19504 7584 19520 7648
rect 19584 7584 19600 7648
rect 19664 7584 19680 7648
rect 19744 7584 19752 7648
rect 19352 6560 19752 7584
rect 19352 6496 19360 6560
rect 19424 6496 19440 6560
rect 19504 6496 19520 6560
rect 19584 6496 19600 6560
rect 19664 6496 19680 6560
rect 19744 6496 19752 6560
rect 19352 5472 19752 6496
rect 19934 6357 19994 9963
rect 19931 6356 19997 6357
rect 19931 6292 19932 6356
rect 19996 6292 19997 6356
rect 19931 6291 19997 6292
rect 19352 5408 19360 5472
rect 19424 5408 19440 5472
rect 19504 5408 19520 5472
rect 19584 5408 19600 5472
rect 19664 5408 19680 5472
rect 19744 5408 19752 5472
rect 19011 5268 19077 5269
rect 19011 5204 19012 5268
rect 19076 5204 19077 5268
rect 19011 5203 19077 5204
rect 19352 4384 19752 5408
rect 19352 4320 19360 4384
rect 19424 4320 19440 4384
rect 19504 4320 19520 4384
rect 19584 4320 19600 4384
rect 19664 4320 19680 4384
rect 19744 4320 19752 4384
rect 19352 3296 19752 4320
rect 20118 3637 20178 12390
rect 20670 12205 20730 17987
rect 21038 17645 21098 20843
rect 21222 19277 21282 22203
rect 21219 19276 21285 19277
rect 21219 19212 21220 19276
rect 21284 19212 21285 19276
rect 21219 19211 21285 19212
rect 21035 17644 21101 17645
rect 21035 17580 21036 17644
rect 21100 17580 21101 17644
rect 21035 17579 21101 17580
rect 20851 12884 20917 12885
rect 20851 12820 20852 12884
rect 20916 12820 20917 12884
rect 20851 12819 20917 12820
rect 20667 12204 20733 12205
rect 20667 12140 20668 12204
rect 20732 12140 20733 12204
rect 20667 12139 20733 12140
rect 20299 9212 20365 9213
rect 20299 9148 20300 9212
rect 20364 9148 20365 9212
rect 20299 9147 20365 9148
rect 20302 7445 20362 9147
rect 20299 7444 20365 7445
rect 20299 7380 20300 7444
rect 20364 7380 20365 7444
rect 20299 7379 20365 7380
rect 20854 5677 20914 12819
rect 20851 5676 20917 5677
rect 20851 5612 20852 5676
rect 20916 5612 20917 5676
rect 20851 5611 20917 5612
rect 21038 4045 21098 17579
rect 21222 12885 21282 19211
rect 21590 18053 21650 22883
rect 22352 22336 22752 23360
rect 22352 22272 22360 22336
rect 22424 22272 22440 22336
rect 22504 22272 22520 22336
rect 22584 22272 22600 22336
rect 22664 22272 22680 22336
rect 22744 22272 22752 22336
rect 22352 21248 22752 22272
rect 22352 21184 22360 21248
rect 22424 21184 22440 21248
rect 22504 21184 22520 21248
rect 22584 21184 22600 21248
rect 22664 21184 22680 21248
rect 22744 21184 22752 21248
rect 22352 20160 22752 21184
rect 22352 20096 22360 20160
rect 22424 20096 22440 20160
rect 22504 20096 22520 20160
rect 22584 20096 22600 20160
rect 22664 20096 22680 20160
rect 22744 20096 22752 20160
rect 22352 19072 22752 20096
rect 22352 19008 22360 19072
rect 22424 19008 22440 19072
rect 22504 19008 22520 19072
rect 22584 19008 22600 19072
rect 22664 19008 22680 19072
rect 22744 19008 22752 19072
rect 21587 18052 21653 18053
rect 21587 17988 21588 18052
rect 21652 17988 21653 18052
rect 21587 17987 21653 17988
rect 21219 12884 21285 12885
rect 21219 12820 21220 12884
rect 21284 12820 21285 12884
rect 21219 12819 21285 12820
rect 21590 4181 21650 17987
rect 22352 17984 22752 19008
rect 22352 17920 22360 17984
rect 22424 17920 22440 17984
rect 22504 17920 22520 17984
rect 22584 17920 22600 17984
rect 22664 17920 22680 17984
rect 22744 17920 22752 17984
rect 22352 16896 22752 17920
rect 22352 16832 22360 16896
rect 22424 16832 22440 16896
rect 22504 16832 22520 16896
rect 22584 16832 22600 16896
rect 22664 16832 22680 16896
rect 22744 16832 22752 16896
rect 22352 15808 22752 16832
rect 22352 15744 22360 15808
rect 22424 15744 22440 15808
rect 22504 15744 22520 15808
rect 22584 15744 22600 15808
rect 22664 15744 22680 15808
rect 22744 15744 22752 15808
rect 22352 14720 22752 15744
rect 22352 14656 22360 14720
rect 22424 14656 22440 14720
rect 22504 14656 22520 14720
rect 22584 14656 22600 14720
rect 22664 14656 22680 14720
rect 22744 14656 22752 14720
rect 22352 13632 22752 14656
rect 22352 13568 22360 13632
rect 22424 13568 22440 13632
rect 22504 13568 22520 13632
rect 22584 13568 22600 13632
rect 22664 13568 22680 13632
rect 22744 13568 22752 13632
rect 22352 12544 22752 13568
rect 22352 12480 22360 12544
rect 22424 12480 22440 12544
rect 22504 12480 22520 12544
rect 22584 12480 22600 12544
rect 22664 12480 22680 12544
rect 22744 12480 22752 12544
rect 22352 11456 22752 12480
rect 22352 11392 22360 11456
rect 22424 11392 22440 11456
rect 22504 11392 22520 11456
rect 22584 11392 22600 11456
rect 22664 11392 22680 11456
rect 22744 11392 22752 11456
rect 22352 10368 22752 11392
rect 22352 10304 22360 10368
rect 22424 10304 22440 10368
rect 22504 10304 22520 10368
rect 22584 10304 22600 10368
rect 22664 10304 22680 10368
rect 22744 10304 22752 10368
rect 22352 9280 22752 10304
rect 22352 9216 22360 9280
rect 22424 9216 22440 9280
rect 22504 9216 22520 9280
rect 22584 9216 22600 9280
rect 22664 9216 22680 9280
rect 22744 9216 22752 9280
rect 22352 8192 22752 9216
rect 22352 8128 22360 8192
rect 22424 8128 22440 8192
rect 22504 8128 22520 8192
rect 22584 8128 22600 8192
rect 22664 8128 22680 8192
rect 22744 8128 22752 8192
rect 22352 7104 22752 8128
rect 22352 7040 22360 7104
rect 22424 7040 22440 7104
rect 22504 7040 22520 7104
rect 22584 7040 22600 7104
rect 22664 7040 22680 7104
rect 22744 7040 22752 7104
rect 22352 6016 22752 7040
rect 22352 5952 22360 6016
rect 22424 5952 22440 6016
rect 22504 5952 22520 6016
rect 22584 5952 22600 6016
rect 22664 5952 22680 6016
rect 22744 5952 22752 6016
rect 22352 4928 22752 5952
rect 22352 4864 22360 4928
rect 22424 4864 22440 4928
rect 22504 4864 22520 4928
rect 22584 4864 22600 4928
rect 22664 4864 22680 4928
rect 22744 4864 22752 4928
rect 21587 4180 21653 4181
rect 21587 4116 21588 4180
rect 21652 4116 21653 4180
rect 21587 4115 21653 4116
rect 21035 4044 21101 4045
rect 21035 3980 21036 4044
rect 21100 3980 21101 4044
rect 21035 3979 21101 3980
rect 21038 3637 21098 3979
rect 22352 3840 22752 4864
rect 22352 3776 22360 3840
rect 22424 3776 22440 3840
rect 22504 3776 22520 3840
rect 22584 3776 22600 3840
rect 22664 3776 22680 3840
rect 22744 3776 22752 3840
rect 20115 3636 20181 3637
rect 20115 3572 20116 3636
rect 20180 3572 20181 3636
rect 20115 3571 20181 3572
rect 21035 3636 21101 3637
rect 21035 3572 21036 3636
rect 21100 3572 21101 3636
rect 21035 3571 21101 3572
rect 19352 3232 19360 3296
rect 19424 3232 19440 3296
rect 19504 3232 19520 3296
rect 19584 3232 19600 3296
rect 19664 3232 19680 3296
rect 19744 3232 19752 3296
rect 19352 2208 19752 3232
rect 19352 2144 19360 2208
rect 19424 2144 19440 2208
rect 19504 2144 19520 2208
rect 19584 2144 19600 2208
rect 19664 2144 19680 2208
rect 19744 2144 19752 2208
rect 18459 2004 18525 2005
rect 18459 1940 18460 2004
rect 18524 1940 18525 2004
rect 18459 1939 18525 1940
rect 16352 1600 16360 1664
rect 16424 1600 16440 1664
rect 16504 1600 16520 1664
rect 16584 1600 16600 1664
rect 16664 1600 16680 1664
rect 16744 1600 16752 1664
rect 14411 1052 14477 1053
rect 14411 988 14412 1052
rect 14476 988 14477 1052
rect 14411 987 14477 988
rect 16352 576 16752 1600
rect 16352 512 16360 576
rect 16424 512 16440 576
rect 16504 512 16520 576
rect 16584 512 16600 576
rect 16664 512 16680 576
rect 16744 512 16752 576
rect 16352 496 16752 512
rect 19352 1120 19752 2144
rect 22352 2752 22752 3776
rect 22352 2688 22360 2752
rect 22424 2688 22440 2752
rect 22504 2688 22520 2752
rect 22584 2688 22600 2752
rect 22664 2688 22680 2752
rect 22744 2688 22752 2752
rect 19931 1732 19997 1733
rect 19931 1668 19932 1732
rect 19996 1668 19997 1732
rect 19931 1667 19997 1668
rect 19352 1056 19360 1120
rect 19424 1056 19440 1120
rect 19504 1056 19520 1120
rect 19584 1056 19600 1120
rect 19664 1056 19680 1120
rect 19744 1056 19752 1120
rect 19352 496 19752 1056
rect 19934 373 19994 1667
rect 22352 1664 22752 2688
rect 22352 1600 22360 1664
rect 22424 1600 22440 1664
rect 22504 1600 22520 1664
rect 22584 1600 22600 1664
rect 22664 1600 22680 1664
rect 22744 1600 22752 1664
rect 22352 576 22752 1600
rect 22352 512 22360 576
rect 22424 512 22440 576
rect 22504 512 22520 576
rect 22584 512 22600 576
rect 22664 512 22680 576
rect 22744 512 22752 576
rect 22352 496 22752 512
rect 11099 372 11165 373
rect 11099 308 11100 372
rect 11164 308 11165 372
rect 11099 307 11165 308
rect 19931 372 19997 373
rect 19931 308 19932 372
rect 19996 308 19997 372
rect 19931 307 19997 308
use sky130_fd_sc_hd__buf_1  _1187_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 5244 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1188_
timestamp 1723858470
transform 1 0 5060 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1189_
timestamp 1723858470
transform 1 0 3312 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1190_
timestamp 1723858470
transform 1 0 3772 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1191_
timestamp 1723858470
transform 1 0 5060 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1192_
timestamp 1723858470
transform 1 0 2392 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1193_
timestamp 1723858470
transform 1 0 6164 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1194_
timestamp 1723858470
transform -1 0 2944 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1195_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3312 0 1 7072
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  _1196_
timestamp 1723858470
transform 1 0 10304 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1197_
timestamp 1723858470
transform -1 0 11592 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1198_
timestamp 1723858470
transform -1 0 8280 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1199_
timestamp 1723858470
transform -1 0 7728 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1200_
timestamp 1723858470
transform -1 0 7176 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1201_
timestamp 1723858470
transform 1 0 4600 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1202_
timestamp 1723858470
transform 1 0 6532 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1203_
timestamp 1723858470
transform 1 0 3680 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1204_
timestamp 1723858470
transform -1 0 1932 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1205_
timestamp 1723858470
transform 1 0 5796 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1206_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 6440 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1207_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 4508 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1208_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 6164 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1209_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 6164 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1210_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5336 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1211_
timestamp 1723858470
transform 1 0 4692 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1212_
timestamp 1723858470
transform -1 0 4324 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1213_
timestamp 1723858470
transform 1 0 4416 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1214_
timestamp 1723858470
transform -1 0 4048 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1215_
timestamp 1723858470
transform 1 0 1840 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1216_
timestamp 1723858470
transform 1 0 2392 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1217_
timestamp 1723858470
transform -1 0 3404 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1218_
timestamp 1723858470
transform 1 0 3864 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1219_
timestamp 1723858470
transform -1 0 5152 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1220_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 4324 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _1221_
timestamp 1723858470
transform -1 0 6440 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1222_
timestamp 1723858470
transform -1 0 13800 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1223_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 11500 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1224_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 7728 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1225_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 5244 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _1226_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 4600 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_2  _1227_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 5060 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1228_
timestamp 1723858470
transform -1 0 23092 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1229_
timestamp 1723858470
transform -1 0 22264 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1230_
timestamp 1723858470
transform -1 0 21436 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1231_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 21988 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1232_
timestamp 1723858470
transform 1 0 20884 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1233_
timestamp 1723858470
transform 1 0 19044 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1234_
timestamp 1723858470
transform 1 0 20608 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1235_
timestamp 1723858470
transform -1 0 21528 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1236_
timestamp 1723858470
transform -1 0 19964 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1237_
timestamp 1723858470
transform -1 0 21620 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1238_
timestamp 1723858470
transform -1 0 21160 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1239_
timestamp 1723858470
transform 1 0 21252 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1240_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 22448 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1241_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 22172 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1242_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 22816 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1243_
timestamp 1723858470
transform 1 0 21620 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1244_
timestamp 1723858470
transform 1 0 22264 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1245_
timestamp 1723858470
transform 1 0 22172 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1246_
timestamp 1723858470
transform 1 0 22816 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1247_
timestamp 1723858470
transform 1 0 5336 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1248_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 8372 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1249_
timestamp 1723858470
transform -1 0 21436 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1250_
timestamp 1723858470
transform -1 0 20608 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1251_
timestamp 1723858470
transform -1 0 20976 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1252_
timestamp 1723858470
transform -1 0 20976 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1253_
timestamp 1723858470
transform -1 0 21988 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1254_
timestamp 1723858470
transform -1 0 21160 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1255_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 19504 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1256_
timestamp 1723858470
transform 1 0 20700 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1257_
timestamp 1723858470
transform -1 0 21252 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1258_
timestamp 1723858470
transform -1 0 20608 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1259_
timestamp 1723858470
transform 1 0 20884 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1260_
timestamp 1723858470
transform 1 0 20700 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1261_
timestamp 1723858470
transform 1 0 21252 0 -1 1632
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1262_
timestamp 1723858470
transform -1 0 5428 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1263_
timestamp 1723858470
transform -1 0 5152 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1264_
timestamp 1723858470
transform -1 0 8004 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1265_
timestamp 1723858470
transform 1 0 5520 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1266_
timestamp 1723858470
transform 1 0 6992 0 1 14688
box -38 -48 958 592
use sky130_fd_sc_hd__and4b_1  _1267_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 7084 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1268_
timestamp 1723858470
transform -1 0 8280 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1269_
timestamp 1723858470
transform 1 0 12052 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1270_
timestamp 1723858470
transform -1 0 12144 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1271_
timestamp 1723858470
transform -1 0 20240 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1272_
timestamp 1723858470
transform -1 0 20056 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1273_
timestamp 1723858470
transform -1 0 20884 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1274_
timestamp 1723858470
transform -1 0 20332 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1275_
timestamp 1723858470
transform 1 0 20240 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1276_
timestamp 1723858470
transform 1 0 14628 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1277_
timestamp 1723858470
transform -1 0 15732 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1278_
timestamp 1723858470
transform 1 0 15088 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1279_
timestamp 1723858470
transform -1 0 19596 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1280_
timestamp 1723858470
transform 1 0 20976 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1281_
timestamp 1723858470
transform -1 0 18584 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1282_
timestamp 1723858470
transform 1 0 19596 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1283_
timestamp 1723858470
transform -1 0 22816 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1284_
timestamp 1723858470
transform -1 0 22816 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1285_
timestamp 1723858470
transform -1 0 23000 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1286_
timestamp 1723858470
transform -1 0 22172 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1287_
timestamp 1723858470
transform -1 0 20148 0 -1 7072
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  _1288_
timestamp 1723858470
transform 1 0 15456 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1289_
timestamp 1723858470
transform -1 0 13432 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1290_
timestamp 1723858470
transform -1 0 11592 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1291_
timestamp 1723858470
transform -1 0 18216 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1292_
timestamp 1723858470
transform 1 0 15916 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1293_
timestamp 1723858470
transform -1 0 13156 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1294_
timestamp 1723858470
transform 1 0 3956 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1295_
timestamp 1723858470
transform -1 0 8372 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _1296_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 10856 0 1 14688
box -38 -48 1970 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1297_
timestamp 1723858470
transform 1 0 12788 0 -1 14688
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1298_
timestamp 1723858470
transform -1 0 22724 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1299_
timestamp 1723858470
transform -1 0 20332 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1300_
timestamp 1723858470
transform -1 0 19504 0 -1 19040
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _1301_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 19964 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1302_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 20516 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1303_
timestamp 1723858470
transform 1 0 13524 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1304_
timestamp 1723858470
transform -1 0 19688 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1305_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 20148 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1306_
timestamp 1723858470
transform 1 0 19596 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _1307_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 19964 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1308_
timestamp 1723858470
transform -1 0 22264 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1309_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 21528 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1310_
timestamp 1723858470
transform -1 0 20332 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1311_
timestamp 1723858470
transform -1 0 20056 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1312_
timestamp 1723858470
transform 1 0 19504 0 1 9248
box -38 -48 958 592
use sky130_fd_sc_hd__o21a_1  _1313_
timestamp 1723858470
transform 1 0 19964 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_2  _1314_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 21252 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _1315_
timestamp 1723858470
transform 1 0 9200 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1316_
timestamp 1723858470
transform -1 0 8372 0 -1 7072
box -38 -48 958 592
use sky130_fd_sc_hd__o31a_1  _1317_
timestamp 1723858470
transform -1 0 20332 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1318_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 20700 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1319_
timestamp 1723858470
transform -1 0 6072 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1320_
timestamp 1723858470
transform -1 0 12696 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1321_
timestamp 1723858470
transform 1 0 13616 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1322_
timestamp 1723858470
transform 1 0 13892 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1323_
timestamp 1723858470
transform 1 0 14076 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1324_
timestamp 1723858470
transform 1 0 15364 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1325_
timestamp 1723858470
transform 1 0 21804 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1326_
timestamp 1723858470
transform -1 0 21528 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _1327_
timestamp 1723858470
transform -1 0 20884 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1328_
timestamp 1723858470
transform 1 0 21896 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1329_
timestamp 1723858470
transform -1 0 21804 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1330_
timestamp 1723858470
transform 1 0 22080 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1331_
timestamp 1723858470
transform 1 0 8464 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1332_
timestamp 1723858470
transform -1 0 9292 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1333_
timestamp 1723858470
transform -1 0 11960 0 1 13600
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1334_
timestamp 1723858470
transform 1 0 12696 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1335_
timestamp 1723858470
transform -1 0 11868 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1336_
timestamp 1723858470
transform 1 0 2208 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1337_
timestamp 1723858470
transform -1 0 2392 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1338_
timestamp 1723858470
transform 1 0 1472 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1339_
timestamp 1723858470
transform 1 0 5428 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1340_
timestamp 1723858470
transform -1 0 6164 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1341_
timestamp 1723858470
transform 1 0 5796 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1342_
timestamp 1723858470
transform -1 0 11960 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1343_
timestamp 1723858470
transform -1 0 11776 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1344_
timestamp 1723858470
transform -1 0 14536 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1345_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 13616 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1346_
timestamp 1723858470
transform 1 0 13892 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1347_
timestamp 1723858470
transform 1 0 13984 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1348_
timestamp 1723858470
transform -1 0 15088 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1349_
timestamp 1723858470
transform 1 0 13524 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1350_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 13616 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1351_
timestamp 1723858470
transform -1 0 13248 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _1352_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 12052 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1353_
timestamp 1723858470
transform 1 0 3588 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1354_
timestamp 1723858470
transform -1 0 4232 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1355_
timestamp 1723858470
transform 1 0 3496 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1356_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5244 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_1  _1357_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 4876 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_2  _1358_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 2392 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1359_
timestamp 1723858470
transform -1 0 2116 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1360_
timestamp 1723858470
transform -1 0 1840 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1361_
timestamp 1723858470
transform 1 0 1840 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1362_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 2024 0 1 19040
box -38 -48 1234 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1363_
timestamp 1723858470
transform 1 0 2116 0 1 9248
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  _1364_
timestamp 1723858470
transform 1 0 2300 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1365_
timestamp 1723858470
transform -1 0 10856 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1366_
timestamp 1723858470
transform 1 0 2392 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1367_
timestamp 1723858470
transform -1 0 3128 0 1 7072
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1368_
timestamp 1723858470
transform -1 0 3772 0 -1 5984
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  _1369_
timestamp 1723858470
transform -1 0 13432 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1370_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 10580 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1371_
timestamp 1723858470
transform -1 0 12144 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1372_
timestamp 1723858470
transform 1 0 4692 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_2  _1373_
timestamp 1723858470
transform 1 0 4232 0 1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_1  _1374_
timestamp 1723858470
transform -1 0 5244 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1375_
timestamp 1723858470
transform 1 0 5796 0 -1 4896
box -38 -48 958 592
use sky130_fd_sc_hd__xor2_1  _1376_
timestamp 1723858470
transform 1 0 5796 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _1377_
timestamp 1723858470
transform -1 0 6992 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1378_
timestamp 1723858470
transform 1 0 6716 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1379_
timestamp 1723858470
transform 1 0 10120 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1380_
timestamp 1723858470
transform 1 0 9476 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1381_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 9936 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1382_
timestamp 1723858470
transform 1 0 11776 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1383_
timestamp 1723858470
transform 1 0 12236 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _1384_
timestamp 1723858470
transform 1 0 12880 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1385_
timestamp 1723858470
transform -1 0 12420 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1386_
timestamp 1723858470
transform -1 0 12052 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1387_
timestamp 1723858470
transform 1 0 13984 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1388_
timestamp 1723858470
transform 1 0 13984 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _1389_
timestamp 1723858470
transform 1 0 15088 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1390_
timestamp 1723858470
transform 1 0 17296 0 1 13600
box -38 -48 958 592
use sky130_fd_sc_hd__or3b_1  _1391_
timestamp 1723858470
transform 1 0 10396 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1392_
timestamp 1723858470
transform 1 0 14628 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _1393_
timestamp 1723858470
transform 1 0 17020 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1394_
timestamp 1723858470
transform 1 0 19780 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1395_
timestamp 1723858470
transform 1 0 19320 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1396_
timestamp 1723858470
transform 1 0 10948 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _1397_
timestamp 1723858470
transform 1 0 10580 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1398_
timestamp 1723858470
transform 1 0 10120 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1399_
timestamp 1723858470
transform 1 0 10948 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _1400_
timestamp 1723858470
transform 1 0 10120 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1401_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 1104 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1402_
timestamp 1723858470
transform 1 0 4140 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1403_
timestamp 1723858470
transform 1 0 4416 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1404_
timestamp 1723858470
transform -1 0 6348 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1405_
timestamp 1723858470
transform 1 0 1380 0 -1 19040
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _1406_
timestamp 1723858470
transform -1 0 9200 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1407_
timestamp 1723858470
transform 1 0 9016 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1408_
timestamp 1723858470
transform -1 0 10120 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1409_
timestamp 1723858470
transform 1 0 10948 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1410_
timestamp 1723858470
transform 1 0 9936 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1411_
timestamp 1723858470
transform -1 0 22540 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1412_
timestamp 1723858470
transform -1 0 21620 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1413_
timestamp 1723858470
transform -1 0 20976 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1414_
timestamp 1723858470
transform -1 0 21896 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1415_
timestamp 1723858470
transform 1 0 19412 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1416_
timestamp 1723858470
transform -1 0 20424 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1417_
timestamp 1723858470
transform -1 0 21896 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _1418_
timestamp 1723858470
transform 1 0 21160 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1419_
timestamp 1723858470
transform -1 0 7176 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1420_
timestamp 1723858470
transform 1 0 18032 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1421_
timestamp 1723858470
transform -1 0 23092 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1422_
timestamp 1723858470
transform -1 0 22540 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1423_
timestamp 1723858470
transform 1 0 22172 0 1 8160
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1424_
timestamp 1723858470
transform -1 0 22172 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1425_
timestamp 1723858470
transform 1 0 20884 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1426_
timestamp 1723858470
transform 1 0 21252 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1427_
timestamp 1723858470
transform 1 0 22724 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1428_
timestamp 1723858470
transform 1 0 5796 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1429_
timestamp 1723858470
transform -1 0 9016 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_2  _1430_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 8372 0 1 13600
box -38 -48 1694 592
use sky130_fd_sc_hd__a22o_1  _1431_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 18860 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1432_
timestamp 1723858470
transform 1 0 19320 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1433_
timestamp 1723858470
transform -1 0 21620 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1434_
timestamp 1723858470
transform -1 0 19412 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1435_
timestamp 1723858470
transform 1 0 20332 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1436_
timestamp 1723858470
transform 1 0 19872 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1437_
timestamp 1723858470
transform 1 0 20056 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1438_
timestamp 1723858470
transform 1 0 19688 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1439_
timestamp 1723858470
transform -1 0 20608 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1440_
timestamp 1723858470
transform -1 0 20332 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1441_
timestamp 1723858470
transform 1 0 18676 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1442_
timestamp 1723858470
transform -1 0 19228 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1443_
timestamp 1723858470
transform -1 0 20332 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1444_
timestamp 1723858470
transform -1 0 20148 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1445_
timestamp 1723858470
transform -1 0 14168 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1446_
timestamp 1723858470
transform -1 0 14628 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1447_
timestamp 1723858470
transform -1 0 18584 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__nand3_2  _1448_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 21160 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1449_
timestamp 1723858470
transform -1 0 12236 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1450_
timestamp 1723858470
transform -1 0 8280 0 1 8160
box -38 -48 958 592
use sky130_fd_sc_hd__xnor2_1  _1451_
timestamp 1723858470
transform 1 0 14444 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1452_
timestamp 1723858470
transform -1 0 20148 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1453_
timestamp 1723858470
transform -1 0 12328 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1454_
timestamp 1723858470
transform 1 0 7820 0 -1 9248
box -38 -48 958 592
use sky130_fd_sc_hd__o21a_1  _1455_
timestamp 1723858470
transform -1 0 16928 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1456_
timestamp 1723858470
transform 1 0 8372 0 1 8160
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1457_
timestamp 1723858470
transform 1 0 20884 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1458_
timestamp 1723858470
transform 1 0 21344 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1459_
timestamp 1723858470
transform 1 0 22080 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1460_
timestamp 1723858470
transform 1 0 17756 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1461_
timestamp 1723858470
transform 1 0 21620 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1462_
timestamp 1723858470
transform -1 0 22080 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1463_
timestamp 1723858470
transform 1 0 21436 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1464_
timestamp 1723858470
transform -1 0 22724 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1465_
timestamp 1723858470
transform -1 0 18584 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1466_
timestamp 1723858470
transform 1 0 18216 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1467_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 18492 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1468_
timestamp 1723858470
transform -1 0 19872 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1469_
timestamp 1723858470
transform 1 0 19688 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1470_
timestamp 1723858470
transform -1 0 19228 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _1471_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 18400 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1472_
timestamp 1723858470
transform 1 0 10212 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1473_
timestamp 1723858470
transform 1 0 17756 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1474_
timestamp 1723858470
transform 1 0 18492 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1475_
timestamp 1723858470
transform -1 0 21620 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _1476_
timestamp 1723858470
transform 1 0 18400 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1477_
timestamp 1723858470
transform -1 0 5336 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1478_
timestamp 1723858470
transform -1 0 21068 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1479_
timestamp 1723858470
transform 1 0 19136 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1480_
timestamp 1723858470
transform -1 0 16560 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1481_
timestamp 1723858470
transform 1 0 12972 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1482_
timestamp 1723858470
transform -1 0 13524 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1483_
timestamp 1723858470
transform 1 0 16100 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1484_
timestamp 1723858470
transform -1 0 21160 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1485_
timestamp 1723858470
transform 1 0 15088 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1486_
timestamp 1723858470
transform -1 0 17480 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1487_
timestamp 1723858470
transform 1 0 17480 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1488_
timestamp 1723858470
transform -1 0 17020 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1489_
timestamp 1723858470
transform 1 0 17756 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1490_
timestamp 1723858470
transform 1 0 20332 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1491_
timestamp 1723858470
transform 1 0 18676 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1492_
timestamp 1723858470
transform -1 0 19688 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1493_
timestamp 1723858470
transform 1 0 19228 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1494_
timestamp 1723858470
transform 1 0 19044 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _1495_
timestamp 1723858470
transform -1 0 16744 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1496_
timestamp 1723858470
transform 1 0 18124 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1497_
timestamp 1723858470
transform -1 0 16468 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1498_
timestamp 1723858470
transform -1 0 19136 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1499_
timestamp 1723858470
transform -1 0 18860 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1500_
timestamp 1723858470
transform -1 0 19596 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1501_
timestamp 1723858470
transform -1 0 19320 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1502_
timestamp 1723858470
transform 1 0 18216 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1503_
timestamp 1723858470
transform 1 0 17480 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1504_
timestamp 1723858470
transform 1 0 18676 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1505_
timestamp 1723858470
transform 1 0 20608 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1506_
timestamp 1723858470
transform -1 0 18952 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1507_
timestamp 1723858470
transform -1 0 18032 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1508_
timestamp 1723858470
transform -1 0 18860 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _1509_
timestamp 1723858470
transform 1 0 11224 0 -1 12512
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_2  _1510_
timestamp 1723858470
transform -1 0 12420 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1511_
timestamp 1723858470
transform -1 0 19228 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1512_
timestamp 1723858470
transform -1 0 13064 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1513_
timestamp 1723858470
transform 1 0 13340 0 -1 10336
box -38 -48 958 592
use sky130_fd_sc_hd__a211oi_1  _1514_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 18308 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1515_
timestamp 1723858470
transform 1 0 17848 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1516_
timestamp 1723858470
transform -1 0 17664 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1517_
timestamp 1723858470
transform 1 0 5796 0 -1 14688
box -38 -48 958 592
use sky130_fd_sc_hd__mux4_2  _1518_
timestamp 1723858470
transform 1 0 6624 0 1 13600
box -38 -48 1694 592
use sky130_fd_sc_hd__a22o_1  _1519_
timestamp 1723858470
transform 1 0 18216 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1520_
timestamp 1723858470
transform 1 0 18768 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1521_
timestamp 1723858470
transform 1 0 18676 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1522_
timestamp 1723858470
transform 1 0 17572 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1523_
timestamp 1723858470
transform -1 0 17940 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1524_
timestamp 1723858470
transform 1 0 17020 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1525_
timestamp 1723858470
transform -1 0 16744 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1526_
timestamp 1723858470
transform -1 0 22172 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1527_
timestamp 1723858470
transform 1 0 20700 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1528_
timestamp 1723858470
transform 1 0 20148 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _1529_
timestamp 1723858470
transform -1 0 16836 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1530_
timestamp 1723858470
transform -1 0 4600 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1531_
timestamp 1723858470
transform -1 0 12144 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1532_
timestamp 1723858470
transform -1 0 17940 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1533_
timestamp 1723858470
transform 1 0 18676 0 1 10336
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1534_
timestamp 1723858470
transform -1 0 19596 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1535_
timestamp 1723858470
transform 1 0 10948 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1536_
timestamp 1723858470
transform 1 0 12696 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1537_
timestamp 1723858470
transform 1 0 12236 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1538_
timestamp 1723858470
transform 1 0 12788 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1539_
timestamp 1723858470
transform 1 0 13708 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1540_
timestamp 1723858470
transform 1 0 17020 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1541_
timestamp 1723858470
transform 1 0 13984 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _1542_
timestamp 1723858470
transform 1 0 15088 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1543_
timestamp 1723858470
transform 1 0 14904 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1544_
timestamp 1723858470
transform -1 0 14904 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1545_
timestamp 1723858470
transform -1 0 14720 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1546_
timestamp 1723858470
transform -1 0 15088 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1547_
timestamp 1723858470
transform 1 0 15088 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1548_
timestamp 1723858470
transform -1 0 14904 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1549_
timestamp 1723858470
transform -1 0 15548 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1550_
timestamp 1723858470
transform -1 0 15272 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1551_
timestamp 1723858470
transform 1 0 18676 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1552_
timestamp 1723858470
transform -1 0 15364 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _1553_
timestamp 1723858470
transform 1 0 15640 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1554_
timestamp 1723858470
transform 1 0 13800 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1555_
timestamp 1723858470
transform 1 0 13340 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1556_
timestamp 1723858470
transform 1 0 13524 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _1557_
timestamp 1723858470
transform -1 0 19596 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1558_
timestamp 1723858470
transform 1 0 14628 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1559_
timestamp 1723858470
transform 1 0 14720 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1560_
timestamp 1723858470
transform 1 0 20148 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1561_
timestamp 1723858470
transform -1 0 17480 0 -1 11424
box -38 -48 958 592
use sky130_fd_sc_hd__o21a_1  _1562_
timestamp 1723858470
transform -1 0 15548 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1563_
timestamp 1723858470
transform 1 0 16100 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1564_
timestamp 1723858470
transform 1 0 16560 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1565_
timestamp 1723858470
transform -1 0 15916 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1566_
timestamp 1723858470
transform 1 0 14812 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1567_
timestamp 1723858470
transform -1 0 13340 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1568_
timestamp 1723858470
transform 1 0 13064 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1569_
timestamp 1723858470
transform -1 0 15640 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1570_
timestamp 1723858470
transform 1 0 14168 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1571_
timestamp 1723858470
transform -1 0 20056 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1572_
timestamp 1723858470
transform 1 0 3772 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1573_
timestamp 1723858470
transform 1 0 3864 0 1 4896
box -38 -48 958 592
use sky130_fd_sc_hd__mux4_2  _1574_
timestamp 1723858470
transform 1 0 6072 0 -1 13600
box -38 -48 1694 592
use sky130_fd_sc_hd__o22a_1  _1575_
timestamp 1723858470
transform 1 0 14536 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1576_
timestamp 1723858470
transform 1 0 14260 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1577_
timestamp 1723858470
transform 1 0 15640 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1578_
timestamp 1723858470
transform 1 0 14904 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1579_
timestamp 1723858470
transform -1 0 15364 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1580_
timestamp 1723858470
transform 1 0 14904 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1581_
timestamp 1723858470
transform 1 0 19780 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1582_
timestamp 1723858470
transform 1 0 14996 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1583_
timestamp 1723858470
transform -1 0 15180 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1584_
timestamp 1723858470
transform -1 0 15364 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1585_
timestamp 1723858470
transform -1 0 15456 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1586_
timestamp 1723858470
transform 1 0 20608 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _1587_
timestamp 1723858470
transform 1 0 14076 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1588_
timestamp 1723858470
transform -1 0 3496 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1589_
timestamp 1723858470
transform 1 0 19780 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1590_
timestamp 1723858470
transform -1 0 14444 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1591_
timestamp 1723858470
transform -1 0 12144 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1592_
timestamp 1723858470
transform -1 0 15088 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1593_
timestamp 1723858470
transform -1 0 6624 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1594_
timestamp 1723858470
transform -1 0 7268 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1595_
timestamp 1723858470
transform 1 0 6532 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1596_
timestamp 1723858470
transform 1 0 7544 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1597_
timestamp 1723858470
transform 1 0 6808 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1598_
timestamp 1723858470
transform 1 0 12144 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1599_
timestamp 1723858470
transform 1 0 8464 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1600_
timestamp 1723858470
transform 1 0 10488 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1601_
timestamp 1723858470
transform 1 0 9844 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1602_
timestamp 1723858470
transform 1 0 14444 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1603_
timestamp 1723858470
transform -1 0 13708 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1604_
timestamp 1723858470
transform 1 0 12788 0 -1 13600
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1605_
timestamp 1723858470
transform 1 0 8188 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1606_
timestamp 1723858470
transform -1 0 9200 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1607_
timestamp 1723858470
transform -1 0 8832 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1608_
timestamp 1723858470
transform -1 0 8924 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1609_
timestamp 1723858470
transform 1 0 8832 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1610_
timestamp 1723858470
transform -1 0 10488 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1611_
timestamp 1723858470
transform -1 0 10764 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1612_
timestamp 1723858470
transform -1 0 10304 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_2  _1613_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 13800 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1614_
timestamp 1723858470
transform 1 0 9384 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1615_
timestamp 1723858470
transform -1 0 9936 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1616_
timestamp 1723858470
transform -1 0 17204 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1617_
timestamp 1723858470
transform -1 0 10488 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1618_
timestamp 1723858470
transform -1 0 13064 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1619_
timestamp 1723858470
transform 1 0 11592 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1620_
timestamp 1723858470
transform 1 0 12420 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1621_
timestamp 1723858470
transform -1 0 11040 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1622_
timestamp 1723858470
transform -1 0 10396 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1623_
timestamp 1723858470
transform 1 0 13064 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1624_
timestamp 1723858470
transform -1 0 13616 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1625_
timestamp 1723858470
transform 1 0 10120 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1626_
timestamp 1723858470
transform -1 0 3956 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_2  _1627_
timestamp 1723858470
transform 1 0 4876 0 1 12512
box -38 -48 1694 592
use sky130_fd_sc_hd__or2_1  _1628_
timestamp 1723858470
transform 1 0 12052 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1629_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 12512 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1630_
timestamp 1723858470
transform 1 0 12512 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1631_
timestamp 1723858470
transform -1 0 20700 0 -1 5984
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1632_
timestamp 1723858470
transform -1 0 12972 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1633_
timestamp 1723858470
transform 1 0 11776 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1634_
timestamp 1723858470
transform 1 0 20424 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1635_
timestamp 1723858470
transform 1 0 11132 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1636_
timestamp 1723858470
transform -1 0 10672 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1637_
timestamp 1723858470
transform -1 0 12052 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1638_
timestamp 1723858470
transform -1 0 11408 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1639_
timestamp 1723858470
transform 1 0 20700 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _1640_
timestamp 1723858470
transform 1 0 11132 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1641_
timestamp 1723858470
transform -1 0 3128 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1642_
timestamp 1723858470
transform 1 0 15364 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1643_
timestamp 1723858470
transform 1 0 10212 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1644_
timestamp 1723858470
transform 1 0 15732 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1645_
timestamp 1723858470
transform -1 0 8648 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1646_
timestamp 1723858470
transform 1 0 10488 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  _1647_
timestamp 1723858470
transform 1 0 4508 0 1 14688
box -38 -48 1694 592
use sky130_fd_sc_hd__o22a_1  _1648_
timestamp 1723858470
transform 1 0 11500 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1649_
timestamp 1723858470
transform 1 0 11224 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1650_
timestamp 1723858470
transform -1 0 14904 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1651_
timestamp 1723858470
transform -1 0 12696 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1652_
timestamp 1723858470
transform -1 0 9660 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1653_
timestamp 1723858470
transform -1 0 9384 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1654_
timestamp 1723858470
transform 1 0 4692 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1655_
timestamp 1723858470
transform -1 0 3680 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1656_
timestamp 1723858470
transform 1 0 4600 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1657_
timestamp 1723858470
transform 1 0 5244 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1658_
timestamp 1723858470
transform 1 0 5060 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1659_
timestamp 1723858470
transform 1 0 6808 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1660_
timestamp 1723858470
transform 1 0 6624 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1661_
timestamp 1723858470
transform 1 0 8004 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1662_
timestamp 1723858470
transform -1 0 8004 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1663_
timestamp 1723858470
transform 1 0 8372 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1664_
timestamp 1723858470
transform -1 0 4324 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1665_
timestamp 1723858470
transform 1 0 4416 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1666_
timestamp 1723858470
transform -1 0 5520 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1667_
timestamp 1723858470
transform -1 0 4876 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1668_
timestamp 1723858470
transform 1 0 4692 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1669_
timestamp 1723858470
transform -1 0 5704 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1670_
timestamp 1723858470
transform 1 0 8372 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1671_
timestamp 1723858470
transform 1 0 5796 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1672_
timestamp 1723858470
transform 1 0 4324 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1673_
timestamp 1723858470
transform -1 0 5520 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1674_
timestamp 1723858470
transform -1 0 4876 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _1675_
timestamp 1723858470
transform 1 0 9660 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1676_
timestamp 1723858470
transform 1 0 5796 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1677_
timestamp 1723858470
transform 1 0 6992 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1678_
timestamp 1723858470
transform 1 0 6532 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1679_
timestamp 1723858470
transform 1 0 6900 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1680_
timestamp 1723858470
transform 1 0 11224 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1681_
timestamp 1723858470
transform -1 0 8096 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1682_
timestamp 1723858470
transform -1 0 9200 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1683_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 11868 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1684_
timestamp 1723858470
transform 1 0 11592 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1685_
timestamp 1723858470
transform -1 0 15916 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1686_
timestamp 1723858470
transform -1 0 12328 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1687_
timestamp 1723858470
transform 1 0 19136 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1688_
timestamp 1723858470
transform -1 0 12972 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1689_
timestamp 1723858470
transform 1 0 12328 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1690_
timestamp 1723858470
transform -1 0 12880 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1691_
timestamp 1723858470
transform -1 0 12328 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1692_
timestamp 1723858470
transform 1 0 20056 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _1693_
timestamp 1723858470
transform 1 0 12328 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1694_
timestamp 1723858470
transform 1 0 2024 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1695_
timestamp 1723858470
transform -1 0 20608 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1696_
timestamp 1723858470
transform -1 0 9936 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1697_
timestamp 1723858470
transform -1 0 11316 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1698_
timestamp 1723858470
transform -1 0 10764 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1699_
timestamp 1723858470
transform -1 0 13892 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1700_
timestamp 1723858470
transform -1 0 15180 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1701_
timestamp 1723858470
transform -1 0 6716 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1702_
timestamp 1723858470
transform 1 0 3128 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1703_
timestamp 1723858470
transform 1 0 4140 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1704_
timestamp 1723858470
transform 1 0 3404 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1705_
timestamp 1723858470
transform -1 0 4692 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1706_
timestamp 1723858470
transform 1 0 3680 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1707_
timestamp 1723858470
transform -1 0 5796 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1708_
timestamp 1723858470
transform 1 0 5796 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1709_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 8280 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1710_
timestamp 1723858470
transform 1 0 6624 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1711_
timestamp 1723858470
transform 1 0 7176 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1712_
timestamp 1723858470
transform 1 0 5520 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1713_
timestamp 1723858470
transform 1 0 4324 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1714_
timestamp 1723858470
transform -1 0 4140 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1715_
timestamp 1723858470
transform -1 0 5612 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1716_
timestamp 1723858470
transform 1 0 5520 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1717_
timestamp 1723858470
transform 1 0 5244 0 -1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _1718_
timestamp 1723858470
transform 1 0 6348 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1719_
timestamp 1723858470
transform 1 0 6532 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1720_
timestamp 1723858470
transform -1 0 4600 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1721_
timestamp 1723858470
transform 1 0 4784 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1722_
timestamp 1723858470
transform -1 0 4784 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_2  _1723_
timestamp 1723858470
transform 1 0 4876 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1724_
timestamp 1723858470
transform 1 0 4692 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1725_
timestamp 1723858470
transform -1 0 7544 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1726_
timestamp 1723858470
transform -1 0 7636 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1727_
timestamp 1723858470
transform 1 0 6992 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1728_
timestamp 1723858470
transform 1 0 7360 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1729_
timestamp 1723858470
transform 1 0 6992 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1730_
timestamp 1723858470
transform -1 0 7820 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1731_
timestamp 1723858470
transform -1 0 12420 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1732_
timestamp 1723858470
transform 1 0 14444 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1733_
timestamp 1723858470
transform -1 0 13432 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1734_
timestamp 1723858470
transform 1 0 5796 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1735_
timestamp 1723858470
transform -1 0 11132 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1736_
timestamp 1723858470
transform -1 0 18492 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1737_
timestamp 1723858470
transform 1 0 8372 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  _1738_
timestamp 1723858470
transform 1 0 4048 0 -1 14688
box -38 -48 1694 592
use sky130_fd_sc_hd__or2_1  _1739_
timestamp 1723858470
transform 1 0 9200 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1740_
timestamp 1723858470
transform 1 0 9568 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1741_
timestamp 1723858470
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _1742_
timestamp 1723858470
transform 1 0 8372 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1743_
timestamp 1723858470
transform -1 0 11224 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1744_
timestamp 1723858470
transform -1 0 8740 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1745_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 19964 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1746_
timestamp 1723858470
transform 1 0 9108 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1747_
timestamp 1723858470
transform -1 0 14168 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1748_
timestamp 1723858470
transform 1 0 13524 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1749_
timestamp 1723858470
transform 1 0 7820 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1750_
timestamp 1723858470
transform 1 0 18952 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1751_
timestamp 1723858470
transform -1 0 8280 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1752_
timestamp 1723858470
transform 1 0 7176 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1753_
timestamp 1723858470
transform 1 0 6072 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1754_
timestamp 1723858470
transform 1 0 4048 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1755_
timestamp 1723858470
transform -1 0 5244 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1756_
timestamp 1723858470
transform 1 0 4232 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1757_
timestamp 1723858470
transform 1 0 4416 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1758_
timestamp 1723858470
transform 1 0 4968 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1759_
timestamp 1723858470
transform 1 0 5888 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1760_
timestamp 1723858470
transform 1 0 6716 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1761_
timestamp 1723858470
transform 1 0 17480 0 -1 11424
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  _1762_
timestamp 1723858470
transform -1 0 6072 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1763_
timestamp 1723858470
transform 1 0 5888 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1764_
timestamp 1723858470
transform 1 0 2024 0 1 10336
box -38 -48 958 592
use sky130_fd_sc_hd__xnor2_1  _1765_
timestamp 1723858470
transform 1 0 2116 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1766_
timestamp 1723858470
transform 1 0 4140 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1767_
timestamp 1723858470
transform 1 0 3128 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1768_
timestamp 1723858470
transform 1 0 3772 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1769_
timestamp 1723858470
transform 1 0 4416 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1770_
timestamp 1723858470
transform 1 0 5796 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1771_
timestamp 1723858470
transform 1 0 3404 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1772_
timestamp 1723858470
transform -1 0 7360 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1773_
timestamp 1723858470
transform 1 0 6256 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1774_
timestamp 1723858470
transform -1 0 7452 0 -1 7072
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1775_
timestamp 1723858470
transform -1 0 7452 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1776_
timestamp 1723858470
transform -1 0 13616 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1777_
timestamp 1723858470
transform 1 0 9660 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1778_
timestamp 1723858470
transform -1 0 5520 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1779_
timestamp 1723858470
transform 1 0 7176 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1780_
timestamp 1723858470
transform -1 0 6900 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1781_
timestamp 1723858470
transform 1 0 9660 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1782_
timestamp 1723858470
transform 1 0 9108 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1783_
timestamp 1723858470
transform 1 0 8556 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _1784_
timestamp 1723858470
transform 1 0 8464 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1785_
timestamp 1723858470
transform 1 0 10028 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1786_
timestamp 1723858470
transform -1 0 10212 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1787_
timestamp 1723858470
transform 1 0 8740 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1788_
timestamp 1723858470
transform 1 0 9292 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1789_
timestamp 1723858470
transform -1 0 10672 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1790_
timestamp 1723858470
transform -1 0 9108 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1791_
timestamp 1723858470
transform 1 0 18400 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1792_
timestamp 1723858470
transform -1 0 8648 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1793_
timestamp 1723858470
transform 1 0 8280 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1794_
timestamp 1723858470
transform 1 0 21804 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1795_
timestamp 1723858470
transform 1 0 19964 0 1 7072
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1796_
timestamp 1723858470
transform -1 0 22724 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1797_
timestamp 1723858470
transform -1 0 21620 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1798_
timestamp 1723858470
transform -1 0 21068 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1799_
timestamp 1723858470
transform 1 0 21252 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1800_
timestamp 1723858470
transform 1 0 20516 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1801_
timestamp 1723858470
transform 1 0 19044 0 -1 14688
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1802_
timestamp 1723858470
transform -1 0 20884 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1803_
timestamp 1723858470
transform -1 0 14720 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1804_
timestamp 1723858470
transform 1 0 6256 0 1 8160
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1805_
timestamp 1723858470
transform 1 0 17664 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1806_
timestamp 1723858470
transform -1 0 18400 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1807_
timestamp 1723858470
transform -1 0 19596 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1808_
timestamp 1723858470
transform 1 0 21988 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__a211oi_1  _1809_
timestamp 1723858470
transform 1 0 21528 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1810_
timestamp 1723858470
transform -1 0 21896 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1811_
timestamp 1723858470
transform -1 0 21988 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1812_
timestamp 1723858470
transform 1 0 22172 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1813_
timestamp 1723858470
transform -1 0 16008 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1814_
timestamp 1723858470
transform 1 0 12880 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1815_
timestamp 1723858470
transform -1 0 18584 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1816_
timestamp 1723858470
transform 1 0 17664 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1817_
timestamp 1723858470
transform 1 0 16744 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1818_
timestamp 1723858470
transform -1 0 16192 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1819_
timestamp 1723858470
transform 1 0 16100 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1820_
timestamp 1723858470
transform 1 0 16744 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1821_
timestamp 1723858470
transform -1 0 17112 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1822_
timestamp 1723858470
transform 1 0 21988 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1823_
timestamp 1723858470
transform 1 0 22264 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1824_
timestamp 1723858470
transform -1 0 21620 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1825_
timestamp 1723858470
transform 1 0 22540 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1826_
timestamp 1723858470
transform -1 0 22724 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1827_
timestamp 1723858470
transform 1 0 17296 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1828_
timestamp 1723858470
transform -1 0 17296 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1829_
timestamp 1723858470
transform -1 0 16928 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1830_
timestamp 1723858470
transform 1 0 16836 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1831_
timestamp 1723858470
transform 1 0 13616 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _1832_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 16100 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _1833_
timestamp 1723858470
transform 1 0 16100 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1834_
timestamp 1723858470
transform 1 0 16836 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1835_
timestamp 1723858470
transform 1 0 17020 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1836_
timestamp 1723858470
transform -1 0 17388 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1837_
timestamp 1723858470
transform 1 0 17020 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1838_
timestamp 1723858470
transform -1 0 14076 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1839_
timestamp 1723858470
transform -1 0 16376 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1840_
timestamp 1723858470
transform 1 0 14904 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1841_
timestamp 1723858470
transform 1 0 21436 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1842_
timestamp 1723858470
transform 1 0 15640 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1843_
timestamp 1723858470
transform 1 0 14536 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1844_
timestamp 1723858470
transform -1 0 15180 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1845_
timestamp 1723858470
transform 1 0 14628 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1846_
timestamp 1723858470
transform 1 0 15364 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1847_
timestamp 1723858470
transform -1 0 16468 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1848_
timestamp 1723858470
transform 1 0 15364 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1849_
timestamp 1723858470
transform 1 0 16284 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1850_
timestamp 1723858470
transform 1 0 16008 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1851_
timestamp 1723858470
transform 1 0 16100 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1852_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 16560 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1853_
timestamp 1723858470
transform 1 0 9292 0 1 14688
box -38 -48 958 592
use sky130_fd_sc_hd__nand3_1  _1854_
timestamp 1723858470
transform -1 0 16008 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1855_
timestamp 1723858470
transform 1 0 17756 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1856_
timestamp 1723858470
transform -1 0 18768 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1857_
timestamp 1723858470
transform 1 0 16744 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1858_
timestamp 1723858470
transform 1 0 15916 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1859_
timestamp 1723858470
transform 1 0 17204 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1860_
timestamp 1723858470
transform 1 0 16100 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1861_
timestamp 1723858470
transform 1 0 15548 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1862_
timestamp 1723858470
transform 1 0 15548 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1863_
timestamp 1723858470
transform -1 0 13984 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1864_
timestamp 1723858470
transform 1 0 17020 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1865_
timestamp 1723858470
transform 1 0 14628 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1866_
timestamp 1723858470
transform 1 0 14076 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1867_
timestamp 1723858470
transform -1 0 14352 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1868_
timestamp 1723858470
transform -1 0 16928 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1869_
timestamp 1723858470
transform 1 0 16284 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1870_
timestamp 1723858470
transform 1 0 12420 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1871_
timestamp 1723858470
transform 1 0 13156 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _1872_
timestamp 1723858470
transform -1 0 14628 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1873_
timestamp 1723858470
transform 1 0 11776 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1874_
timestamp 1723858470
transform 1 0 12144 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1875_
timestamp 1723858470
transform 1 0 12604 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1876_
timestamp 1723858470
transform 1 0 14812 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1877_
timestamp 1723858470
transform 1 0 12696 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1878_
timestamp 1723858470
transform -1 0 14536 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1879_
timestamp 1723858470
transform -1 0 14260 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _1880_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 13800 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _1881_
timestamp 1723858470
transform 1 0 13064 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _1882_
timestamp 1723858470
transform 1 0 13432 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1883_
timestamp 1723858470
transform -1 0 15088 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1884_
timestamp 1723858470
transform -1 0 14996 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1885_
timestamp 1723858470
transform -1 0 15088 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1886_
timestamp 1723858470
transform -1 0 14628 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1887_
timestamp 1723858470
transform -1 0 12696 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1888_
timestamp 1723858470
transform -1 0 20700 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1889_
timestamp 1723858470
transform -1 0 14444 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1890_
timestamp 1723858470
transform -1 0 14720 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1891_
timestamp 1723858470
transform -1 0 15732 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1892_
timestamp 1723858470
transform -1 0 21528 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1893_
timestamp 1723858470
transform 1 0 10948 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1894_
timestamp 1723858470
transform 1 0 11224 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1895_
timestamp 1723858470
transform 1 0 6624 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1896_
timestamp 1723858470
transform -1 0 6716 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1897_
timestamp 1723858470
transform -1 0 6256 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _1898_
timestamp 1723858470
transform 1 0 5796 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1899_
timestamp 1723858470
transform 1 0 12328 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1900_
timestamp 1723858470
transform 1 0 12788 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1901_
timestamp 1723858470
transform 1 0 5796 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _1902_
timestamp 1723858470
transform 1 0 3772 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1903_
timestamp 1723858470
transform 1 0 3956 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1904_
timestamp 1723858470
transform 1 0 3956 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1905_
timestamp 1723858470
transform -1 0 5152 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _1906_
timestamp 1723858470
transform -1 0 12696 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1907_
timestamp 1723858470
transform 1 0 4232 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1908_
timestamp 1723858470
transform 1 0 7176 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1909_
timestamp 1723858470
transform -1 0 8188 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _1910_
timestamp 1723858470
transform -1 0 7636 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1911_
timestamp 1723858470
transform 1 0 7544 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1912_
timestamp 1723858470
transform 1 0 12420 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1913_
timestamp 1723858470
transform 1 0 11592 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1914_
timestamp 1723858470
transform -1 0 19596 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1915_
timestamp 1723858470
transform -1 0 11776 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1916_
timestamp 1723858470
transform -1 0 12972 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1917_
timestamp 1723858470
transform 1 0 11316 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1918_
timestamp 1723858470
transform -1 0 11592 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1919_
timestamp 1723858470
transform -1 0 11868 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1920_
timestamp 1723858470
transform 1 0 11592 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1921_
timestamp 1723858470
transform 1 0 21436 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1922_
timestamp 1723858470
transform -1 0 14168 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1923_
timestamp 1723858470
transform 1 0 11776 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1924_
timestamp 1723858470
transform 1 0 11960 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1925_
timestamp 1723858470
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1926_
timestamp 1723858470
transform -1 0 6440 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1927_
timestamp 1723858470
transform 1 0 5244 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1928_
timestamp 1723858470
transform -1 0 6256 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1929_
timestamp 1723858470
transform 1 0 6624 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _1930_
timestamp 1723858470
transform -1 0 6624 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1931_
timestamp 1723858470
transform 1 0 5980 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _1932_
timestamp 1723858470
transform 1 0 2576 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1933_
timestamp 1723858470
transform -1 0 3128 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1934_
timestamp 1723858470
transform 1 0 3496 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1935_
timestamp 1723858470
transform -1 0 4876 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1936_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3956 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1937_
timestamp 1723858470
transform 1 0 3956 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1938_
timestamp 1723858470
transform -1 0 6992 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1939_
timestamp 1723858470
transform 1 0 6440 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _1940_
timestamp 1723858470
transform -1 0 6532 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1941_
timestamp 1723858470
transform -1 0 14168 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1942_
timestamp 1723858470
transform 1 0 13248 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__o221ai_1  _1943_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 13064 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1944_
timestamp 1723858470
transform -1 0 13340 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1945_
timestamp 1723858470
transform -1 0 13708 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1946_
timestamp 1723858470
transform 1 0 9844 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1947_
timestamp 1723858470
transform 1 0 10396 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1948_
timestamp 1723858470
transform 1 0 10948 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1949_
timestamp 1723858470
transform 1 0 8832 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1950_
timestamp 1723858470
transform 1 0 5152 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1951_
timestamp 1723858470
transform -1 0 3680 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1952_
timestamp 1723858470
transform -1 0 3864 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _1953_
timestamp 1723858470
transform 1 0 3680 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1954_
timestamp 1723858470
transform 1 0 4232 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _1955_
timestamp 1723858470
transform -1 0 2392 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1956_
timestamp 1723858470
transform -1 0 1748 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1957_
timestamp 1723858470
transform -1 0 2392 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1958_
timestamp 1723858470
transform -1 0 2116 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1959_
timestamp 1723858470
transform 1 0 3404 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1960_
timestamp 1723858470
transform 1 0 2116 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1961_
timestamp 1723858470
transform 1 0 6072 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1962_
timestamp 1723858470
transform -1 0 5796 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1963_
timestamp 1723858470
transform 1 0 5152 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1964_
timestamp 1723858470
transform 1 0 5244 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _1965_
timestamp 1723858470
transform 1 0 8372 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _1966_
timestamp 1723858470
transform 1 0 8188 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1967_
timestamp 1723858470
transform 1 0 8188 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1968_
timestamp 1723858470
transform 1 0 8464 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1969_
timestamp 1723858470
transform 1 0 8188 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1970_
timestamp 1723858470
transform 1 0 7728 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1971_
timestamp 1723858470
transform -1 0 5520 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1972_
timestamp 1723858470
transform 1 0 8740 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1973_
timestamp 1723858470
transform 1 0 9292 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1974_
timestamp 1723858470
transform -1 0 6256 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1975_
timestamp 1723858470
transform 1 0 920 0 1 9248
box -38 -48 1234 592
use sky130_fd_sc_hd__o21a_1  _1976_
timestamp 1723858470
transform 1 0 6992 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1977_
timestamp 1723858470
transform -1 0 3220 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1978_
timestamp 1723858470
transform 1 0 1104 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1979_
timestamp 1723858470
transform 1 0 1472 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1980_
timestamp 1723858470
transform -1 0 2208 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1981_
timestamp 1723858470
transform -1 0 1840 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1982_
timestamp 1723858470
transform -1 0 1472 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1983_
timestamp 1723858470
transform 1 0 828 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1984_
timestamp 1723858470
transform 1 0 1748 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1985_
timestamp 1723858470
transform 1 0 3220 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1986_
timestamp 1723858470
transform -1 0 6624 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1987_
timestamp 1723858470
transform -1 0 5704 0 -1 16864
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1988_
timestamp 1723858470
transform -1 0 9384 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1989_
timestamp 1723858470
transform -1 0 9384 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1990_
timestamp 1723858470
transform 1 0 9384 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _1991_
timestamp 1723858470
transform 1 0 9568 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1992_
timestamp 1723858470
transform -1 0 9844 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1993_
timestamp 1723858470
transform 1 0 13892 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1994_
timestamp 1723858470
transform 1 0 12328 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1995_
timestamp 1723858470
transform -1 0 22448 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1996_
timestamp 1723858470
transform 1 0 21436 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1997_
timestamp 1723858470
transform 1 0 21252 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_1  _1998_
timestamp 1723858470
transform 1 0 21896 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1999_
timestamp 1723858470
transform 1 0 16376 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2000_
timestamp 1723858470
transform -1 0 17940 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2001_
timestamp 1723858470
transform 1 0 16928 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2002_
timestamp 1723858470
transform -1 0 15916 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2003_
timestamp 1723858470
transform 1 0 12880 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2004_
timestamp 1723858470
transform 1 0 14996 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2005_
timestamp 1723858470
transform -1 0 17020 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2006_
timestamp 1723858470
transform 1 0 16100 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2007_
timestamp 1723858470
transform 1 0 18400 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2008_
timestamp 1723858470
transform -1 0 17848 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2009_
timestamp 1723858470
transform 1 0 17204 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2010_
timestamp 1723858470
transform 1 0 17664 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _2011_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 17756 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2012_
timestamp 1723858470
transform -1 0 22540 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _2013_
timestamp 1723858470
transform -1 0 22632 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2014_
timestamp 1723858470
transform 1 0 22540 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2015_
timestamp 1723858470
transform -1 0 22632 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2016_
timestamp 1723858470
transform 1 0 22724 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2017_
timestamp 1723858470
transform 1 0 14076 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2018_
timestamp 1723858470
transform -1 0 14076 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2019_
timestamp 1723858470
transform -1 0 14812 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2020_
timestamp 1723858470
transform -1 0 15916 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2021_
timestamp 1723858470
transform -1 0 15640 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _2022_
timestamp 1723858470
transform 1 0 13892 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2023_
timestamp 1723858470
transform -1 0 14076 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2024_
timestamp 1723858470
transform -1 0 13984 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2025_
timestamp 1723858470
transform 1 0 13984 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2026_
timestamp 1723858470
transform -1 0 18124 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _2027_
timestamp 1723858470
transform 1 0 17020 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _2028_
timestamp 1723858470
transform 1 0 14444 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2029_
timestamp 1723858470
transform 1 0 15456 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2030_
timestamp 1723858470
transform 1 0 14904 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2031_
timestamp 1723858470
transform -1 0 15824 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2032_
timestamp 1723858470
transform 1 0 21620 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _2033_
timestamp 1723858470
transform 1 0 15180 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2034_
timestamp 1723858470
transform 1 0 16100 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _2035_
timestamp 1723858470
transform 1 0 16836 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _2036_
timestamp 1723858470
transform 1 0 18124 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2037_
timestamp 1723858470
transform -1 0 9200 0 -1 8160
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _2038_
timestamp 1723858470
transform -1 0 17848 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _2039_
timestamp 1723858470
transform -1 0 19320 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2040_
timestamp 1723858470
transform 1 0 18860 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2041_
timestamp 1723858470
transform -1 0 22908 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2042_
timestamp 1723858470
transform 1 0 22632 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2043_
timestamp 1723858470
transform -1 0 10856 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2044_
timestamp 1723858470
transform -1 0 11316 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2045_
timestamp 1723858470
transform -1 0 10856 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _2046_
timestamp 1723858470
transform 1 0 13340 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _2047_
timestamp 1723858470
transform 1 0 10948 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _2048_
timestamp 1723858470
transform -1 0 14444 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _2049_
timestamp 1723858470
transform 1 0 3404 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2050_
timestamp 1723858470
transform 1 0 4048 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2051_
timestamp 1723858470
transform -1 0 11868 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2052_
timestamp 1723858470
transform 1 0 11040 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2053_
timestamp 1723858470
transform -1 0 11592 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _2054_
timestamp 1723858470
transform 1 0 15456 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _2055_
timestamp 1723858470
transform 1 0 16008 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2056_
timestamp 1723858470
transform 1 0 16100 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _2057_
timestamp 1723858470
transform 1 0 16284 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _2058_
timestamp 1723858470
transform -1 0 16652 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2059_
timestamp 1723858470
transform -1 0 16836 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2060_
timestamp 1723858470
transform 1 0 19596 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2061_
timestamp 1723858470
transform 1 0 22172 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2062_
timestamp 1723858470
transform 1 0 2668 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2063_
timestamp 1723858470
transform -1 0 3680 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2064_
timestamp 1723858470
transform -1 0 3772 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2065_
timestamp 1723858470
transform 1 0 11592 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _2066_
timestamp 1723858470
transform 1 0 3956 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2067_
timestamp 1723858470
transform -1 0 4324 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2068_
timestamp 1723858470
transform -1 0 3864 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _2069_
timestamp 1723858470
transform 1 0 3128 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2070_
timestamp 1723858470
transform 1 0 3680 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2071_
timestamp 1723858470
transform 1 0 3680 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _2072_
timestamp 1723858470
transform 1 0 3312 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2073_
timestamp 1723858470
transform 1 0 4140 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2074_
timestamp 1723858470
transform -1 0 11224 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _2075_
timestamp 1723858470
transform 1 0 13892 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2076_
timestamp 1723858470
transform 1 0 13524 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2077_
timestamp 1723858470
transform 1 0 14628 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2078_
timestamp 1723858470
transform -1 0 14812 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _2079_
timestamp 1723858470
transform 1 0 14168 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2080_
timestamp 1723858470
transform -1 0 14996 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2081_
timestamp 1723858470
transform -1 0 15640 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2082_
timestamp 1723858470
transform 1 0 19964 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2083_
timestamp 1723858470
transform -1 0 17848 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _2084_
timestamp 1723858470
transform -1 0 20332 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2085_
timestamp 1723858470
transform 1 0 2852 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2086_
timestamp 1723858470
transform 1 0 1932 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2087_
timestamp 1723858470
transform -1 0 3404 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _2088_
timestamp 1723858470
transform -1 0 2484 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _2089_
timestamp 1723858470
transform 1 0 2484 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _2090_
timestamp 1723858470
transform 1 0 3220 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2091_
timestamp 1723858470
transform -1 0 1472 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2092_
timestamp 1723858470
transform 1 0 828 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _2093_
timestamp 1723858470
transform 1 0 1196 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _2094_
timestamp 1723858470
transform 1 0 1196 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2095_
timestamp 1723858470
transform 1 0 2944 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2096_
timestamp 1723858470
transform -1 0 7636 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _2097_
timestamp 1723858470
transform -1 0 8280 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2098_
timestamp 1723858470
transform -1 0 10396 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _2099_
timestamp 1723858470
transform 1 0 10396 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2100_
timestamp 1723858470
transform -1 0 10396 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _2101_
timestamp 1723858470
transform 1 0 9936 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2102_
timestamp 1723858470
transform 1 0 10672 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2103_
timestamp 1723858470
transform 1 0 10948 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2104_
timestamp 1723858470
transform -1 0 11040 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2105_
timestamp 1723858470
transform -1 0 20332 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2106_
timestamp 1723858470
transform 1 0 2392 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2107_
timestamp 1723858470
transform 1 0 1748 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2108_
timestamp 1723858470
transform -1 0 2576 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2109_
timestamp 1723858470
transform 1 0 2852 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2110_
timestamp 1723858470
transform 1 0 2576 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2111_
timestamp 1723858470
transform -1 0 1932 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2112_
timestamp 1723858470
transform -1 0 1932 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2113_
timestamp 1723858470
transform -1 0 2208 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2114_
timestamp 1723858470
transform -1 0 1472 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _2115_
timestamp 1723858470
transform 1 0 1012 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2116_
timestamp 1723858470
transform -1 0 4692 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2117_
timestamp 1723858470
transform -1 0 4692 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _2118_
timestamp 1723858470
transform 1 0 4784 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _2119_
timestamp 1723858470
transform -1 0 9108 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2120_
timestamp 1723858470
transform 1 0 10304 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _2121_
timestamp 1723858470
transform 1 0 10948 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2122_
timestamp 1723858470
transform 1 0 10396 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _2123_
timestamp 1723858470
transform 1 0 10396 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2124_
timestamp 1723858470
transform 1 0 11500 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2125_
timestamp 1723858470
transform 1 0 11776 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2126_
timestamp 1723858470
transform -1 0 12696 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2127_
timestamp 1723858470
transform -1 0 19964 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2128_
timestamp 1723858470
transform 1 0 2300 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _2129_
timestamp 1723858470
transform -1 0 1564 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _2130_
timestamp 1723858470
transform 1 0 1288 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2131_
timestamp 1723858470
transform 1 0 2024 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2132_
timestamp 1723858470
transform 1 0 6440 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _2133_
timestamp 1723858470
transform 1 0 6716 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _2134_
timestamp 1723858470
transform 1 0 11776 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _2135_
timestamp 1723858470
transform 1 0 12420 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2136_
timestamp 1723858470
transform 1 0 13524 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _2137_
timestamp 1723858470
transform 1 0 12972 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2138_
timestamp 1723858470
transform 1 0 13892 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2139_
timestamp 1723858470
transform 1 0 13616 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2140_
timestamp 1723858470
transform 1 0 13524 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2141_
timestamp 1723858470
transform 1 0 17756 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2142_
timestamp 1723858470
transform 1 0 19044 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _2143_
timestamp 1723858470
transform -1 0 3220 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _2144_
timestamp 1723858470
transform 1 0 2208 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2145_
timestamp 1723858470
transform 1 0 2760 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _2146_
timestamp 1723858470
transform 1 0 2392 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2147_
timestamp 1723858470
transform 1 0 2760 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2148_
timestamp 1723858470
transform 1 0 2116 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2149_
timestamp 1723858470
transform 1 0 1932 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2150_
timestamp 1723858470
transform 1 0 2576 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2151_
timestamp 1723858470
transform 1 0 3220 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _2152_
timestamp 1723858470
transform 1 0 2392 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _2153_
timestamp 1723858470
transform 1 0 3128 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2154_
timestamp 1723858470
transform -1 0 4140 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2155_
timestamp 1723858470
transform 1 0 3404 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _2156_
timestamp 1723858470
transform -1 0 6072 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2157_
timestamp 1723858470
transform -1 0 7084 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2158_
timestamp 1723858470
transform -1 0 8004 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _2159_
timestamp 1723858470
transform -1 0 8188 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _2160_
timestamp 1723858470
transform 1 0 10120 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2161_
timestamp 1723858470
transform 1 0 9200 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2162_
timestamp 1723858470
transform -1 0 9200 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _2163_
timestamp 1723858470
transform 1 0 9200 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2164_
timestamp 1723858470
transform -1 0 8464 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2165_
timestamp 1723858470
transform 1 0 9568 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _2166_
timestamp 1723858470
transform 1 0 10212 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2167_
timestamp 1723858470
transform 1 0 9200 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2168_
timestamp 1723858470
transform -1 0 10672 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2169_
timestamp 1723858470
transform 1 0 8648 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2170_
timestamp 1723858470
transform -1 0 8096 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _2171_
timestamp 1723858470
transform -1 0 19596 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2172_
timestamp 1723858470
transform -1 0 9292 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2173_
timestamp 1723858470
transform -1 0 8924 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2174_
timestamp 1723858470
transform 1 0 8924 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2175_
timestamp 1723858470
transform 1 0 20332 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2176_
timestamp 1723858470
transform 1 0 19964 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2177_
timestamp 1723858470
transform -1 0 17940 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _2178_
timestamp 1723858470
transform 1 0 21988 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _2179_
timestamp 1723858470
transform 1 0 22540 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2180_
timestamp 1723858470
transform -1 0 20608 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2181_
timestamp 1723858470
transform -1 0 13984 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _2182_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 21436 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2183_
timestamp 1723858470
transform -1 0 10120 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _2184_
timestamp 1723858470
transform -1 0 9384 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _2185_
timestamp 1723858470
transform 1 0 3312 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2186_
timestamp 1723858470
transform -1 0 12880 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _2187_
timestamp 1723858470
transform 1 0 8372 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _2188_
timestamp 1723858470
transform 1 0 4232 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _2189_
timestamp 1723858470
transform 1 0 3864 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _2190_
timestamp 1723858470
transform 1 0 4232 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _2191_
timestamp 1723858470
transform 1 0 8004 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2192_
timestamp 1723858470
transform 1 0 8556 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _2193_
timestamp 1723858470
transform -1 0 10396 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2194_
timestamp 1723858470
transform 1 0 8740 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _2195_
timestamp 1723858470
transform -1 0 6256 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _2196_
timestamp 1723858470
transform 1 0 9936 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _2197_
timestamp 1723858470
transform -1 0 10856 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _2198_
timestamp 1723858470
transform -1 0 21528 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _2199_
timestamp 1723858470
transform -1 0 11040 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2200_
timestamp 1723858470
transform 1 0 11132 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2201_
timestamp 1723858470
transform -1 0 11960 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2202_
timestamp 1723858470
transform -1 0 9844 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2203_
timestamp 1723858470
transform -1 0 9660 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2204_
timestamp 1723858470
transform -1 0 9936 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _2205_
timestamp 1723858470
transform -1 0 7820 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2206_
timestamp 1723858470
transform 1 0 8740 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _2207_
timestamp 1723858470
transform 1 0 8372 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _2208_
timestamp 1723858470
transform -1 0 9292 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _2209_
timestamp 1723858470
transform -1 0 6440 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2210_
timestamp 1723858470
transform -1 0 6716 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2211_
timestamp 1723858470
transform -1 0 5980 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _2212_
timestamp 1723858470
transform -1 0 8648 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2213_
timestamp 1723858470
transform -1 0 6900 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2214_
timestamp 1723858470
transform 1 0 5796 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _2215_
timestamp 1723858470
transform -1 0 5704 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _2216_
timestamp 1723858470
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _2217_
timestamp 1723858470
transform 1 0 5888 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2218_
timestamp 1723858470
transform 1 0 1840 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _2219_
timestamp 1723858470
transform 1 0 8832 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2220_
timestamp 1723858470
transform -1 0 2116 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2221_
timestamp 1723858470
transform 1 0 1564 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2222_
timestamp 1723858470
transform -1 0 3128 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2223_
timestamp 1723858470
transform 1 0 2392 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2224_
timestamp 1723858470
transform -1 0 3128 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2225_
timestamp 1723858470
transform -1 0 3128 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2226_
timestamp 1723858470
transform 1 0 2852 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2227_
timestamp 1723858470
transform -1 0 3128 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2228_
timestamp 1723858470
transform 1 0 2392 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2229_
timestamp 1723858470
transform 1 0 3128 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2230_
timestamp 1723858470
transform -1 0 12236 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _2231_
timestamp 1723858470
transform -1 0 12144 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _2232_
timestamp 1723858470
transform -1 0 8280 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2233_
timestamp 1723858470
transform 1 0 5428 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _2234_
timestamp 1723858470
transform -1 0 11960 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2235_
timestamp 1723858470
transform -1 0 8832 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _2236_
timestamp 1723858470
transform -1 0 7176 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2237_
timestamp 1723858470
transform 1 0 5796 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_2  _2238_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 6532 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _2239_
timestamp 1723858470
transform 1 0 16836 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2240_
timestamp 1723858470
transform 1 0 16376 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _2241_
timestamp 1723858470
transform 1 0 17296 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _2242_
timestamp 1723858470
transform -1 0 21160 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2243_
timestamp 1723858470
transform 1 0 17572 0 1 19040
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _2244_
timestamp 1723858470
transform 1 0 16652 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2245_
timestamp 1723858470
transform 1 0 18676 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _2246_
timestamp 1723858470
transform 1 0 17572 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _2247_
timestamp 1723858470
transform -1 0 18492 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2248_
timestamp 1723858470
transform -1 0 17664 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2249_
timestamp 1723858470
transform 1 0 18676 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _2250_
timestamp 1723858470
transform 1 0 17664 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _2251_
timestamp 1723858470
transform 1 0 19136 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2252_
timestamp 1723858470
transform -1 0 18216 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _2253_
timestamp 1723858470
transform -1 0 15456 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2254_
timestamp 1723858470
transform -1 0 17204 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _2255_
timestamp 1723858470
transform 1 0 14904 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _2256_
timestamp 1723858470
transform -1 0 15824 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2257_
timestamp 1723858470
transform -1 0 14352 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2258_
timestamp 1723858470
transform -1 0 14812 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _2259_
timestamp 1723858470
transform 1 0 13984 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _2260_
timestamp 1723858470
transform 1 0 15456 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2261_
timestamp 1723858470
transform -1 0 13984 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _2262_
timestamp 1723858470
transform -1 0 12420 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2263_
timestamp 1723858470
transform -1 0 13340 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _2264_
timestamp 1723858470
transform 1 0 12512 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _2265_
timestamp 1723858470
transform -1 0 13800 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2266_
timestamp 1723858470
transform -1 0 11868 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2267_
timestamp 1723858470
transform 1 0 11960 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2268_
timestamp 1723858470
transform 1 0 11868 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2269_
timestamp 1723858470
transform -1 0 12696 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2270_
timestamp 1723858470
transform 1 0 10948 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2271_
timestamp 1723858470
transform 1 0 11592 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _2272_
timestamp 1723858470
transform -1 0 11592 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _2273_
timestamp 1723858470
transform -1 0 10488 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2274_
timestamp 1723858470
transform -1 0 1380 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _2275_
timestamp 1723858470
transform -1 0 11684 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2276_
timestamp 1723858470
transform -1 0 2392 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _2277_
timestamp 1723858470
transform 1 0 1380 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _2278_
timestamp 1723858470
transform 1 0 2392 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _2279_
timestamp 1723858470
transform 1 0 1656 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2280_
timestamp 1723858470
transform 1 0 2024 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2281_
timestamp 1723858470
transform -1 0 1564 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2282_
timestamp 1723858470
transform -1 0 1380 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2283_
timestamp 1723858470
transform -1 0 1288 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2284_
timestamp 1723858470
transform -1 0 1380 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _2285_
timestamp 1723858470
transform 1 0 1380 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _2286_
timestamp 1723858470
transform 1 0 828 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _2287_
timestamp 1723858470
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2288_
timestamp 1723858470
transform 1 0 920 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2289_
timestamp 1723858470
transform 1 0 828 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _2290_
timestamp 1723858470
transform 1 0 1472 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _2291_
timestamp 1723858470
transform 1 0 1840 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2292_
timestamp 1723858470
transform -1 0 1840 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2293_
timestamp 1723858470
transform 1 0 1656 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2294_
timestamp 1723858470
transform 1 0 1196 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2295_
timestamp 1723858470
transform 1 0 3404 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2296_
timestamp 1723858470
transform 1 0 20332 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2297_
timestamp 1723858470
transform -1 0 14904 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _2298_
timestamp 1723858470
transform -1 0 23092 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2299_
timestamp 1723858470
transform -1 0 21436 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _2300_
timestamp 1723858470
transform 1 0 19320 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _2301_
timestamp 1723858470
transform 1 0 20148 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _2302_
timestamp 1723858470
transform 1 0 20792 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _2303_
timestamp 1723858470
transform -1 0 19320 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2304_
timestamp 1723858470
transform 1 0 17572 0 -1 21216
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _2305_
timestamp 1723858470
transform 1 0 15732 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2306_
timestamp 1723858470
transform -1 0 15916 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2307_
timestamp 1723858470
transform -1 0 20792 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2308_
timestamp 1723858470
transform 1 0 16468 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2309_
timestamp 1723858470
transform 1 0 16560 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _2310_
timestamp 1723858470
transform 1 0 15088 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2311_
timestamp 1723858470
transform -1 0 20884 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2312_
timestamp 1723858470
transform 1 0 17020 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2313_
timestamp 1723858470
transform -1 0 14628 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2314_
timestamp 1723858470
transform -1 0 21160 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2315_
timestamp 1723858470
transform -1 0 15548 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2316_
timestamp 1723858470
transform -1 0 15640 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _2317_
timestamp 1723858470
transform 1 0 15732 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2318_
timestamp 1723858470
transform -1 0 20976 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _2319_
timestamp 1723858470
transform 1 0 15732 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2320_
timestamp 1723858470
transform 1 0 19504 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2321_
timestamp 1723858470
transform -1 0 13432 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2322_
timestamp 1723858470
transform -1 0 20240 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2323_
timestamp 1723858470
transform -1 0 19596 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2324_
timestamp 1723858470
transform 1 0 22816 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2325_
timestamp 1723858470
transform -1 0 21160 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2326_
timestamp 1723858470
transform 1 0 18676 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2327_
timestamp 1723858470
transform -1 0 16376 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2328_
timestamp 1723858470
transform -1 0 20516 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2329_
timestamp 1723858470
transform -1 0 19872 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2330_
timestamp 1723858470
transform 1 0 20884 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2331_
timestamp 1723858470
transform 1 0 7268 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _2332_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 9016 0 -1 16864
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _2333_
timestamp 1723858470
transform -1 0 8648 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _2334_
timestamp 1723858470
transform 1 0 6992 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _2335_
timestamp 1723858470
transform -1 0 8740 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _2336_
timestamp 1723858470
transform -1 0 8924 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _2337_
timestamp 1723858470
transform 1 0 6716 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2338_
timestamp 1723858470
transform 1 0 7084 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2339_
timestamp 1723858470
transform 1 0 7728 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2340_
timestamp 1723858470
transform 1 0 8924 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2341_
timestamp 1723858470
transform 1 0 7728 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2342_
timestamp 1723858470
transform 1 0 8740 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _2343_
timestamp 1723858470
transform 1 0 7360 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _2344_
timestamp 1723858470
transform 1 0 6440 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2345_
timestamp 1723858470
transform -1 0 7728 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2346_
timestamp 1723858470
transform 1 0 7176 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _2347_
timestamp 1723858470
transform -1 0 10672 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2348_
timestamp 1723858470
transform -1 0 11960 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2349_
timestamp 1723858470
transform -1 0 11500 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _2350_
timestamp 1723858470
transform 1 0 11040 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _2351_
timestamp 1723858470
transform 1 0 13524 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2352_
timestamp 1723858470
transform -1 0 8648 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _2353_
timestamp 1723858470
transform -1 0 8832 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _2354_
timestamp 1723858470
transform 1 0 9292 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2355_
timestamp 1723858470
transform 1 0 10580 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2356_
timestamp 1723858470
transform -1 0 11684 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2357_
timestamp 1723858470
transform -1 0 16376 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _2358_
timestamp 1723858470
transform -1 0 3496 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _2359_
timestamp 1723858470
transform -1 0 11132 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _2360_
timestamp 1723858470
transform 1 0 9752 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2361_
timestamp 1723858470
transform -1 0 10856 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2362_
timestamp 1723858470
transform 1 0 10028 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2363_
timestamp 1723858470
transform 1 0 9936 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2364_
timestamp 1723858470
transform -1 0 11224 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _2365_
timestamp 1723858470
transform -1 0 8648 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2366_
timestamp 1723858470
transform -1 0 9384 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _2367_
timestamp 1723858470
transform 1 0 9476 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _2368_
timestamp 1723858470
transform -1 0 10028 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2369_
timestamp 1723858470
transform 1 0 10028 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _2370_
timestamp 1723858470
transform 1 0 6164 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _2371_
timestamp 1723858470
transform 1 0 8004 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _2372_
timestamp 1723858470
transform 1 0 18676 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _2373_
timestamp 1723858470
transform 1 0 9292 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _2374_
timestamp 1723858470
transform 1 0 8648 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _2375_
timestamp 1723858470
transform -1 0 9292 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2376_
timestamp 1723858470
transform -1 0 3404 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _2377_
timestamp 1723858470
transform -1 0 4140 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2378_
timestamp 1723858470
transform -1 0 3036 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2379_
timestamp 1723858470
transform -1 0 3680 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2380_
timestamp 1723858470
transform -1 0 3128 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2381_
timestamp 1723858470
transform -1 0 1932 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2382_
timestamp 1723858470
transform -1 0 3036 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2383_
timestamp 1723858470
transform 1 0 1564 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2384_
timestamp 1723858470
transform 1 0 2116 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2385_
timestamp 1723858470
transform -1 0 2760 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2386_
timestamp 1723858470
transform 1 0 3772 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2387_
timestamp 1723858470
transform 1 0 2208 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _2388_
timestamp 1723858470
transform 1 0 2484 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _2389_
timestamp 1723858470
transform -1 0 2944 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2390_
timestamp 1723858470
transform -1 0 2576 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2391_
timestamp 1723858470
transform 1 0 2484 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2392_
timestamp 1723858470
transform 1 0 2576 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2393_
timestamp 1723858470
transform 1 0 3496 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2394_
timestamp 1723858470
transform -1 0 6992 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _2395_
timestamp 1723858470
transform 1 0 5060 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_2  _2396_
timestamp 1723858470
transform 1 0 5428 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _2397_
timestamp 1723858470
transform -1 0 8004 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _2398_
timestamp 1723858470
transform 1 0 6532 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2399_
timestamp 1723858470
transform 1 0 7176 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2400_
timestamp 1723858470
transform -1 0 7360 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2401_
timestamp 1723858470
transform 1 0 9016 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _2402_
timestamp 1723858470
transform -1 0 9016 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2403_
timestamp 1723858470
transform 1 0 7912 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _2404_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 6624 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _2405_
timestamp 1723858470
transform -1 0 7912 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2406_
timestamp 1723858470
transform 1 0 6716 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2407_
timestamp 1723858470
transform -1 0 6716 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2408_
timestamp 1723858470
transform 1 0 22448 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2409_
timestamp 1723858470
transform 1 0 22816 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2410_
timestamp 1723858470
transform -1 0 22540 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2411_
timestamp 1723858470
transform 1 0 22264 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2412_
timestamp 1723858470
transform -1 0 21160 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2413_
timestamp 1723858470
transform -1 0 21712 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2414_
timestamp 1723858470
transform -1 0 21252 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2415_
timestamp 1723858470
transform -1 0 21528 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2416_
timestamp 1723858470
transform -1 0 20332 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2417_
timestamp 1723858470
transform 1 0 21252 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _2418_
timestamp 1723858470
transform 1 0 9016 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2419_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 21620 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2420_
timestamp 1723858470
transform -1 0 23092 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2421_
timestamp 1723858470
transform -1 0 22724 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2422_
timestamp 1723858470
transform -1 0 22816 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2423_
timestamp 1723858470
transform -1 0 23000 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2424_
timestamp 1723858470
transform 1 0 10948 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2425_
timestamp 1723858470
transform 1 0 11960 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2426_
timestamp 1723858470
transform 1 0 9384 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2427_
timestamp 1723858470
transform 1 0 9016 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2428_
timestamp 1723858470
transform 1 0 5796 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2429_
timestamp 1723858470
transform 1 0 828 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2430_
timestamp 1723858470
transform 1 0 920 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2431_
timestamp 1723858470
transform 1 0 2760 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2432_
timestamp 1723858470
transform 1 0 3220 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2433_
timestamp 1723858470
transform 1 0 920 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2434_
timestamp 1723858470
transform 1 0 18676 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2435_
timestamp 1723858470
transform 1 0 18768 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2436_
timestamp 1723858470
transform 1 0 16100 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2437_
timestamp 1723858470
transform 1 0 14628 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2438_
timestamp 1723858470
transform 1 0 13708 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2439_
timestamp 1723858470
transform 1 0 12236 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2440_
timestamp 1723858470
transform -1 0 10856 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2441_
timestamp 1723858470
transform 1 0 2024 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2442_
timestamp 1723858470
transform 1 0 1012 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2443_
timestamp 1723858470
transform 1 0 828 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2444_
timestamp 1723858470
transform 1 0 1288 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2445_
timestamp 1723858470
transform -1 0 2392 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2446_
timestamp 1723858470
transform 1 0 16744 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2447_
timestamp 1723858470
transform 1 0 16100 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2448_
timestamp 1723858470
transform 1 0 15548 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2449_
timestamp 1723858470
transform -1 0 16008 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2450_
timestamp 1723858470
transform 1 0 18676 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2451_
timestamp 1723858470
transform -1 0 18768 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2452_
timestamp 1723858470
transform 1 0 16560 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2453_
timestamp 1723858470
transform -1 0 18584 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2454_
timestamp 1723858470
transform 1 0 6808 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2455_
timestamp 1723858470
transform -1 0 13616 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2456_
timestamp 1723858470
transform 1 0 11776 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2457_
timestamp 1723858470
transform 1 0 11960 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2458_
timestamp 1723858470
transform 1 0 10028 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2459_
timestamp 1723858470
transform -1 0 10028 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2460_
timestamp 1723858470
transform 1 0 3220 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2461_
timestamp 1723858470
transform -1 0 2300 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2462_
timestamp 1723858470
transform 1 0 3220 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2463_
timestamp 1723858470
transform 1 0 2944 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2464_
timestamp 1723858470
transform 1 0 3128 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2465_
timestamp 1723858470
transform 1 0 6440 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2466_
timestamp 1723858470
transform -1 0 23092 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2467_
timestamp 1723858470
transform 1 0 21252 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2468_
timestamp 1723858470
transform 1 0 21620 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2469_
timestamp 1723858470
transform 1 0 21620 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2470_
timestamp 1723858470
transform 1 0 21620 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2471_
timestamp 1723858470
transform 1 0 21620 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2472_
timestamp 1723858470
transform -1 0 23092 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2473_
timestamp 1723858470
transform 1 0 21344 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2474_
timestamp 1723858470
transform 1 0 19412 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2475_
timestamp 1723858470
transform -1 0 6808 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _2476_
timestamp 1723858470
transform 1 0 1656 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2477_
timestamp 1723858470
transform 1 0 828 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2478_
timestamp 1723858470
transform -1 0 7728 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2479_
timestamp 1723858470
transform -1 0 7452 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2480_
timestamp 1723858470
transform -1 0 18952 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2481_
timestamp 1723858470
transform -1 0 18124 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 1564 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1723858470
transform 1 0 12512 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 13432 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_clk
timestamp 1723858470
transform -1 0 5704 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_clk
timestamp 1723858470
transform -1 0 5060 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_clk
timestamp 1723858470
transform 1 0 4876 0 1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_clk
timestamp 1723858470
transform 1 0 9016 0 -1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_clk
timestamp 1723858470
transform 1 0 16836 0 -1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_clk
timestamp 1723858470
transform 1 0 19412 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_clk
timestamp 1723858470
transform -1 0 16744 0 1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_clk
timestamp 1723858470
transform 1 0 18676 0 -1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 828 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_57
timestamp 1723858470
transform 1 0 5796 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_62
timestamp 1723858470
transform 1 0 6256 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_82 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 8096 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_113
timestamp 1723858470
transform 1 0 10948 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_118
timestamp 1723858470
transform 1 0 11408 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 1723858470
transform 1 0 13340 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_169 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 16100 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_176 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 16744 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_184
timestamp 1723858470
transform 1 0 17480 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_195
timestamp 1723858470
transform 1 0 18492 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_223
timestamp 1723858470
transform 1 0 21068 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_11
timestamp 1723858470
transform 1 0 1564 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_15
timestamp 1723858470
transform 1 0 1932 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_23
timestamp 1723858470
transform 1 0 2668 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_49
timestamp 1723858470
transform 1 0 5060 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_64
timestamp 1723858470
transform 1 0 6440 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_90
timestamp 1723858470
transform 1 0 8832 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_110
timestamp 1723858470
transform 1 0 10672 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_113
timestamp 1723858470
transform 1 0 10948 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_122
timestamp 1723858470
transform 1 0 11776 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_146
timestamp 1723858470
transform 1 0 13984 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_162
timestamp 1723858470
transform 1 0 15456 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1723858470
transform 1 0 15916 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_169
timestamp 1723858470
transform 1 0 16100 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_177
timestamp 1723858470
transform 1 0 16836 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_183
timestamp 1723858470
transform 1 0 17388 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_189
timestamp 1723858470
transform 1 0 17940 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_193
timestamp 1723858470
transform 1 0 18308 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_204
timestamp 1723858470
transform 1 0 19320 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1723858470
transform 1 0 21068 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_243
timestamp 1723858470
transform 1 0 22908 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_6
timestamp 1723858470
transform 1 0 1104 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_14 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 1840 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_24
timestamp 1723858470
transform 1 0 2760 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_29
timestamp 1723858470
transform 1 0 3220 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_39
timestamp 1723858470
transform 1 0 4140 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_44
timestamp 1723858470
transform 1 0 4600 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_48
timestamp 1723858470
transform 1 0 4968 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_52
timestamp 1723858470
transform 1 0 5336 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_59
timestamp 1723858470
transform 1 0 5980 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_66 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 6624 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_72
timestamp 1723858470
transform 1 0 7176 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_76
timestamp 1723858470
transform 1 0 7544 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_80
timestamp 1723858470
transform 1 0 7912 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_85
timestamp 1723858470
transform 1 0 8372 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_108
timestamp 1723858470
transform 1 0 10488 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_126
timestamp 1723858470
transform 1 0 12144 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_132
timestamp 1723858470
transform 1 0 12696 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_137
timestamp 1723858470
transform 1 0 13156 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_141
timestamp 1723858470
transform 1 0 13524 0 1 1632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_147 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 14076 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_159
timestamp 1723858470
transform 1 0 15180 0 1 1632
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_167
timestamp 1723858470
transform 1 0 15916 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_179
timestamp 1723858470
transform 1 0 17020 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_191
timestamp 1723858470
transform 1 0 18124 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1723858470
transform 1 0 18492 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_200
timestamp 1723858470
transform 1 0 18952 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_218
timestamp 1723858470
transform 1 0 20608 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_231
timestamp 1723858470
transform 1 0 21804 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_244
timestamp 1723858470
transform 1 0 23000 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1723858470
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_15
timestamp 1723858470
transform 1 0 1932 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_23
timestamp 1723858470
transform 1 0 2668 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_47
timestamp 1723858470
transform 1 0 4876 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_57
timestamp 1723858470
transform 1 0 5796 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_77
timestamp 1723858470
transform 1 0 7636 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_87
timestamp 1723858470
transform 1 0 8556 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_93
timestamp 1723858470
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_110
timestamp 1723858470
transform 1 0 10672 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_116
timestamp 1723858470
transform 1 0 11224 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_148
timestamp 1723858470
transform 1 0 14168 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_152
timestamp 1723858470
transform 1 0 14536 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_164
timestamp 1723858470
transform 1 0 15640 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_177
timestamp 1723858470
transform 1 0 16836 0 -1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_183
timestamp 1723858470
transform 1 0 17388 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_203
timestamp 1723858470
transform 1 0 19228 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_211
timestamp 1723858470
transform 1 0 19964 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_215
timestamp 1723858470
transform 1 0 20332 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_222
timestamp 1723858470
transform 1 0 20976 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_233
timestamp 1723858470
transform 1 0 21988 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_243
timestamp 1723858470
transform 1 0 22908 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_3
timestamp 1723858470
transform 1 0 828 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_20
timestamp 1723858470
transform 1 0 2392 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_36
timestamp 1723858470
transform 1 0 3864 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_55
timestamp 1723858470
transform 1 0 5612 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_62
timestamp 1723858470
transform 1 0 6256 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_76
timestamp 1723858470
transform 1 0 7544 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_85
timestamp 1723858470
transform 1 0 8372 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_100
timestamp 1723858470
transform 1 0 9752 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_105
timestamp 1723858470
transform 1 0 10212 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_113
timestamp 1723858470
transform 1 0 10948 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_121
timestamp 1723858470
transform 1 0 11684 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_126
timestamp 1723858470
transform 1 0 12144 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_134
timestamp 1723858470
transform 1 0 12880 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_148
timestamp 1723858470
transform 1 0 14168 0 1 2720
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_159
timestamp 1723858470
transform 1 0 15180 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_174
timestamp 1723858470
transform 1 0 16560 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_178
timestamp 1723858470
transform 1 0 16928 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_186
timestamp 1723858470
transform 1 0 17664 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_191
timestamp 1723858470
transform 1 0 18124 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1723858470
transform 1 0 18492 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_197
timestamp 1723858470
transform 1 0 18676 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_201
timestamp 1723858470
transform 1 0 19044 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_205
timestamp 1723858470
transform 1 0 19412 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_212
timestamp 1723858470
transform 1 0 20056 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_3
timestamp 1723858470
transform 1 0 828 0 -1 3808
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_13
timestamp 1723858470
transform 1 0 1748 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_25
timestamp 1723858470
transform 1 0 2852 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_33
timestamp 1723858470
transform 1 0 3588 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_41
timestamp 1723858470
transform 1 0 4324 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_46
timestamp 1723858470
transform 1 0 4784 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_54
timestamp 1723858470
transform 1 0 5520 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_57
timestamp 1723858470
transform 1 0 5796 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_65
timestamp 1723858470
transform 1 0 6532 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_77
timestamp 1723858470
transform 1 0 7636 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_120
timestamp 1723858470
transform 1 0 11592 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_135
timestamp 1723858470
transform 1 0 12972 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_141
timestamp 1723858470
transform 1 0 13524 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_149
timestamp 1723858470
transform 1 0 14260 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_158
timestamp 1723858470
transform 1 0 15088 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_166
timestamp 1723858470
transform 1 0 15824 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_176
timestamp 1723858470
transform 1 0 16744 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_180
timestamp 1723858470
transform 1 0 17112 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_184
timestamp 1723858470
transform 1 0 17480 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_189
timestamp 1723858470
transform 1 0 17940 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_193
timestamp 1723858470
transform 1 0 18308 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_211
timestamp 1723858470
transform 1 0 19964 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_225
timestamp 1723858470
transform 1 0 21252 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_238
timestamp 1723858470
transform 1 0 22448 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_243
timestamp 1723858470
transform 1 0 22908 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_3
timestamp 1723858470
transform 1 0 828 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_14
timestamp 1723858470
transform 1 0 1840 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_29
timestamp 1723858470
transform 1 0 3220 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_33
timestamp 1723858470
transform 1 0 3588 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_44
timestamp 1723858470
transform 1 0 4600 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_64
timestamp 1723858470
transform 1 0 6440 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_90
timestamp 1723858470
transform 1 0 8832 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_94
timestamp 1723858470
transform 1 0 9200 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_111
timestamp 1723858470
transform 1 0 10764 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_116
timestamp 1723858470
transform 1 0 11224 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_136
timestamp 1723858470
transform 1 0 13064 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_141
timestamp 1723858470
transform 1 0 13524 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_148
timestamp 1723858470
transform 1 0 14168 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_167
timestamp 1723858470
transform 1 0 15916 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_175
timestamp 1723858470
transform 1 0 16652 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_187
timestamp 1723858470
transform 1 0 17756 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1723858470
transform 1 0 18492 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_197
timestamp 1723858470
transform 1 0 18676 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_201
timestamp 1723858470
transform 1 0 19044 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_205
timestamp 1723858470
transform 1 0 19412 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_212
timestamp 1723858470
transform 1 0 20056 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_222
timestamp 1723858470
transform 1 0 20976 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_232
timestamp 1723858470
transform 1 0 21896 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_240
timestamp 1723858470
transform 1 0 22632 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_244
timestamp 1723858470
transform 1 0 23000 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_10
timestamp 1723858470
transform 1 0 1472 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_37
timestamp 1723858470
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_42
timestamp 1723858470
transform 1 0 4416 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_79
timestamp 1723858470
transform 1 0 7820 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_108
timestamp 1723858470
transform 1 0 10488 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_113
timestamp 1723858470
transform 1 0 10948 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_119
timestamp 1723858470
transform 1 0 11500 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_133
timestamp 1723858470
transform 1 0 12788 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_159
timestamp 1723858470
transform 1 0 15180 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1723858470
transform 1 0 15916 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_176
timestamp 1723858470
transform 1 0 16744 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_189
timestamp 1723858470
transform 1 0 17940 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_203
timestamp 1723858470
transform 1 0 19228 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_207
timestamp 1723858470
transform 1 0 19596 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_211
timestamp 1723858470
transform 1 0 19964 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_235
timestamp 1723858470
transform 1 0 22172 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_239
timestamp 1723858470
transform 1 0 22540 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_3
timestamp 1723858470
transform 1 0 828 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_13
timestamp 1723858470
transform 1 0 1748 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_20
timestamp 1723858470
transform 1 0 2392 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_26
timestamp 1723858470
transform 1 0 2944 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_29
timestamp 1723858470
transform 1 0 3220 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_54
timestamp 1723858470
transform 1 0 5520 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_75
timestamp 1723858470
transform 1 0 7452 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_85
timestamp 1723858470
transform 1 0 8372 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_96
timestamp 1723858470
transform 1 0 9384 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_135
timestamp 1723858470
transform 1 0 12972 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1723858470
transform 1 0 13340 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_156
timestamp 1723858470
transform 1 0 14904 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_160
timestamp 1723858470
transform 1 0 15272 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_170
timestamp 1723858470
transform 1 0 16192 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_177
timestamp 1723858470
transform 1 0 16836 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_188
timestamp 1723858470
transform 1 0 17848 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_225
timestamp 1723858470
transform 1 0 21252 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_234
timestamp 1723858470
transform 1 0 22080 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_242
timestamp 1723858470
transform 1 0 22816 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_16
timestamp 1723858470
transform 1 0 2024 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_24
timestamp 1723858470
transform 1 0 2760 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_38
timestamp 1723858470
transform 1 0 4048 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_45
timestamp 1723858470
transform 1 0 4692 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1723858470
transform 1 0 5612 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_60
timestamp 1723858470
transform 1 0 6072 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_73
timestamp 1723858470
transform 1 0 7268 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_101
timestamp 1723858470
transform 1 0 9844 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_113
timestamp 1723858470
transform 1 0 10948 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_129
timestamp 1723858470
transform 1 0 12420 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_142
timestamp 1723858470
transform 1 0 13616 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_154
timestamp 1723858470
transform 1 0 14720 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_164
timestamp 1723858470
transform 1 0 15640 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_169
timestamp 1723858470
transform 1 0 16100 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_182
timestamp 1723858470
transform 1 0 17296 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_191
timestamp 1723858470
transform 1 0 18124 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_200
timestamp 1723858470
transform 1 0 18952 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_222
timestamp 1723858470
transform 1 0 20976 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_225
timestamp 1723858470
transform 1 0 21252 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_242
timestamp 1723858470
transform 1 0 22816 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_3
timestamp 1723858470
transform 1 0 828 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_11
timestamp 1723858470
transform 1 0 1564 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_20
timestamp 1723858470
transform 1 0 2392 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_24
timestamp 1723858470
transform 1 0 2760 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_29
timestamp 1723858470
transform 1 0 3220 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_47
timestamp 1723858470
transform 1 0 4876 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_63
timestamp 1723858470
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1723858470
transform 1 0 7636 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1723858470
transform 1 0 8188 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_93
timestamp 1723858470
transform 1 0 9108 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_99
timestamp 1723858470
transform 1 0 9660 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_111
timestamp 1723858470
transform 1 0 10764 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_115
timestamp 1723858470
transform 1 0 11132 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_119
timestamp 1723858470
transform 1 0 11500 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_128
timestamp 1723858470
transform 1 0 12328 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_141
timestamp 1723858470
transform 1 0 13524 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_154
timestamp 1723858470
transform 1 0 14720 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_174
timestamp 1723858470
transform 1 0 16560 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_185
timestamp 1723858470
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_206
timestamp 1723858470
transform 1 0 19504 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_215
timestamp 1723858470
transform 1 0 20332 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_228
timestamp 1723858470
transform 1 0 21528 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_240
timestamp 1723858470
transform 1 0 22632 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_244
timestamp 1723858470
transform 1 0 23000 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_3
timestamp 1723858470
transform 1 0 828 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_18
timestamp 1723858470
transform 1 0 2208 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_29
timestamp 1723858470
transform 1 0 3220 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_37
timestamp 1723858470
transform 1 0 3956 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_45
timestamp 1723858470
transform 1 0 4692 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_96
timestamp 1723858470
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_127
timestamp 1723858470
transform 1 0 12236 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_146
timestamp 1723858470
transform 1 0 13984 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_164
timestamp 1723858470
transform 1 0 15640 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_178
timestamp 1723858470
transform 1 0 16928 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_187
timestamp 1723858470
transform 1 0 17756 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_191
timestamp 1723858470
transform 1 0 18124 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_196
timestamp 1723858470
transform 1 0 18584 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_202
timestamp 1723858470
transform 1 0 19136 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_221
timestamp 1723858470
transform 1 0 20884 0 -1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_232
timestamp 1723858470
transform 1 0 21896 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_244
timestamp 1723858470
transform 1 0 23000 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_3
timestamp 1723858470
transform 1 0 828 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_11
timestamp 1723858470
transform 1 0 1564 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_29
timestamp 1723858470
transform 1 0 3220 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_40
timestamp 1723858470
transform 1 0 4232 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_45
timestamp 1723858470
transform 1 0 4692 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_57
timestamp 1723858470
transform 1 0 5796 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_66
timestamp 1723858470
transform 1 0 6624 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_80
timestamp 1723858470
transform 1 0 7912 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_97
timestamp 1723858470
transform 1 0 9476 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_108
timestamp 1723858470
transform 1 0 10488 0 1 7072
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_120
timestamp 1723858470
transform 1 0 11592 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_132
timestamp 1723858470
transform 1 0 12696 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_155
timestamp 1723858470
transform 1 0 14812 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_161
timestamp 1723858470
transform 1 0 15364 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_165
timestamp 1723858470
transform 1 0 15732 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_173
timestamp 1723858470
transform 1 0 16468 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_180
timestamp 1723858470
transform 1 0 17112 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1723858470
transform 1 0 18492 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_197
timestamp 1723858470
transform 1 0 18676 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_203
timestamp 1723858470
transform 1 0 19228 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_221
timestamp 1723858470
transform 1 0 20884 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_238
timestamp 1723858470
transform 1 0 22448 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_244
timestamp 1723858470
transform 1 0 23000 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_18
timestamp 1723858470
transform 1 0 2208 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_38
timestamp 1723858470
transform 1 0 4048 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_49
timestamp 1723858470
transform 1 0 5060 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1723858470
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_57
timestamp 1723858470
transform 1 0 5796 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_83
timestamp 1723858470
transform 1 0 8188 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_98
timestamp 1723858470
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1723858470
transform 1 0 10764 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_122
timestamp 1723858470
transform 1 0 11776 0 -1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_129
timestamp 1723858470
transform 1 0 12420 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_141
timestamp 1723858470
transform 1 0 13524 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_157
timestamp 1723858470
transform 1 0 14996 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_161
timestamp 1723858470
transform 1 0 15364 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1723858470
transform 1 0 16100 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_181
timestamp 1723858470
transform 1 0 17204 0 -1 8160
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_210
timestamp 1723858470
transform 1 0 19872 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_222
timestamp 1723858470
transform 1 0 20976 0 -1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_230
timestamp 1723858470
transform 1 0 21712 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_242
timestamp 1723858470
transform 1 0 22816 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_3
timestamp 1723858470
transform 1 0 828 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_7
timestamp 1723858470
transform 1 0 1196 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_15
timestamp 1723858470
transform 1 0 1932 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_23
timestamp 1723858470
transform 1 0 2668 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1723858470
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_29
timestamp 1723858470
transform 1 0 3220 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_39
timestamp 1723858470
transform 1 0 4140 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_47
timestamp 1723858470
transform 1 0 4876 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_57
timestamp 1723858470
transform 1 0 5796 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_72
timestamp 1723858470
transform 1 0 7176 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_111
timestamp 1723858470
transform 1 0 10764 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_126
timestamp 1723858470
transform 1 0 12144 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_138
timestamp 1723858470
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_148
timestamp 1723858470
transform 1 0 14168 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_160
timestamp 1723858470
transform 1 0 15272 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_193
timestamp 1723858470
transform 1 0 18308 0 1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_197
timestamp 1723858470
transform 1 0 18676 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_215
timestamp 1723858470
transform 1 0 20332 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_219
timestamp 1723858470
transform 1 0 20700 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_223
timestamp 1723858470
transform 1 0 21068 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_230
timestamp 1723858470
transform 1 0 21712 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_3
timestamp 1723858470
transform 1 0 828 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_9
timestamp 1723858470
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_14
timestamp 1723858470
transform 1 0 1840 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_35
timestamp 1723858470
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_43
timestamp 1723858470
transform 1 0 4508 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1723858470
transform 1 0 5612 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_63
timestamp 1723858470
transform 1 0 6348 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_69
timestamp 1723858470
transform 1 0 6900 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_76
timestamp 1723858470
transform 1 0 7544 0 -1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_94
timestamp 1723858470
transform 1 0 9200 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_106
timestamp 1723858470
transform 1 0 10304 0 -1 9248
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_118
timestamp 1723858470
transform 1 0 11408 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_130
timestamp 1723858470
transform 1 0 12512 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_142
timestamp 1723858470
transform 1 0 13616 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1723858470
transform 1 0 15916 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_174
timestamp 1723858470
transform 1 0 16560 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_186
timestamp 1723858470
transform 1 0 17664 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_206
timestamp 1723858470
transform 1 0 19504 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_215
timestamp 1723858470
transform 1 0 20332 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 1723858470
transform 1 0 21068 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_228
timestamp 1723858470
transform 1 0 21528 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_232
timestamp 1723858470
transform 1 0 21896 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_244
timestamp 1723858470
transform 1 0 23000 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_3
timestamp 1723858470
transform 1 0 828 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1723858470
transform 1 0 3036 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_50
timestamp 1723858470
transform 1 0 5152 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_64
timestamp 1723858470
transform 1 0 6440 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1723858470
transform 1 0 8188 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_88
timestamp 1723858470
transform 1 0 8648 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1723858470
transform 1 0 13340 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_141
timestamp 1723858470
transform 1 0 13524 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_150
timestamp 1723858470
transform 1 0 14352 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_162
timestamp 1723858470
transform 1 0 15456 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_170
timestamp 1723858470
transform 1 0 16192 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_178
timestamp 1723858470
transform 1 0 16928 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_189
timestamp 1723858470
transform 1 0 17940 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1723858470
transform 1 0 18492 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_197
timestamp 1723858470
transform 1 0 18676 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_224
timestamp 1723858470
transform 1 0 21160 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_244
timestamp 1723858470
transform 1 0 23000 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_27
timestamp 1723858470
transform 1 0 3036 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_34
timestamp 1723858470
transform 1 0 3680 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_45
timestamp 1723858470
transform 1 0 4692 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_53
timestamp 1723858470
transform 1 0 5428 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_70
timestamp 1723858470
transform 1 0 6992 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_75
timestamp 1723858470
transform 1 0 7452 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_97
timestamp 1723858470
transform 1 0 9476 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_107
timestamp 1723858470
transform 1 0 10396 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1723858470
transform 1 0 10764 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_113
timestamp 1723858470
transform 1 0 10948 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_121
timestamp 1723858470
transform 1 0 11684 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_128
timestamp 1723858470
transform 1 0 12328 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_132
timestamp 1723858470
transform 1 0 12696 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_149
timestamp 1723858470
transform 1 0 14260 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_158
timestamp 1723858470
transform 1 0 15088 0 -1 10336
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_172
timestamp 1723858470
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_184
timestamp 1723858470
transform 1 0 17480 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_189
timestamp 1723858470
transform 1 0 17940 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_194
timestamp 1723858470
transform 1 0 18400 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_210
timestamp 1723858470
transform 1 0 19872 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_222
timestamp 1723858470
transform 1 0 20976 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_232
timestamp 1723858470
transform 1 0 21896 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_3
timestamp 1723858470
transform 1 0 828 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_11
timestamp 1723858470
transform 1 0 1564 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_15
timestamp 1723858470
transform 1 0 1932 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_26
timestamp 1723858470
transform 1 0 2944 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_29
timestamp 1723858470
transform 1 0 3220 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_37
timestamp 1723858470
transform 1 0 3956 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_46
timestamp 1723858470
transform 1 0 4784 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_50
timestamp 1723858470
transform 1 0 5152 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_62
timestamp 1723858470
transform 1 0 6256 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_66
timestamp 1723858470
transform 1 0 6624 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_75
timestamp 1723858470
transform 1 0 7452 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1723858470
transform 1 0 8188 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_85
timestamp 1723858470
transform 1 0 8372 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_96
timestamp 1723858470
transform 1 0 9384 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_100
timestamp 1723858470
transform 1 0 9752 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1723858470
transform 1 0 13340 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_141
timestamp 1723858470
transform 1 0 13524 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_145
timestamp 1723858470
transform 1 0 13892 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_150
timestamp 1723858470
transform 1 0 14352 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_154
timestamp 1723858470
transform 1 0 14720 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_162
timestamp 1723858470
transform 1 0 15456 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_180
timestamp 1723858470
transform 1 0 17112 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_191
timestamp 1723858470
transform 1 0 18124 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_221
timestamp 1723858470
transform 1 0 20884 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_228
timestamp 1723858470
transform 1 0 21528 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_3
timestamp 1723858470
transform 1 0 828 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_21
timestamp 1723858470
transform 1 0 2484 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_44
timestamp 1723858470
transform 1 0 4600 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_50
timestamp 1723858470
transform 1 0 5152 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_64
timestamp 1723858470
transform 1 0 6440 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_82
timestamp 1723858470
transform 1 0 8096 0 -1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_91
timestamp 1723858470
transform 1 0 8924 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_103
timestamp 1723858470
transform 1 0 10028 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_107
timestamp 1723858470
transform 1 0 10396 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1723858470
transform 1 0 10764 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_113
timestamp 1723858470
transform 1 0 10948 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_123
timestamp 1723858470
transform 1 0 11868 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_127
timestamp 1723858470
transform 1 0 12236 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_152
timestamp 1723858470
transform 1 0 14536 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1723858470
transform 1 0 15916 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_172
timestamp 1723858470
transform 1 0 16376 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_206
timestamp 1723858470
transform 1 0 19504 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_3
timestamp 1723858470
transform 1 0 828 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_21
timestamp 1723858470
transform 1 0 2484 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_47
timestamp 1723858470
transform 1 0 4876 0 1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_54
timestamp 1723858470
transform 1 0 5520 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_66
timestamp 1723858470
transform 1 0 6624 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_78
timestamp 1723858470
transform 1 0 7728 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_88
timestamp 1723858470
transform 1 0 8648 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_97
timestamp 1723858470
transform 1 0 9476 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_127
timestamp 1723858470
transform 1 0 12236 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1723858470
transform 1 0 13340 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_141
timestamp 1723858470
transform 1 0 13524 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_152
timestamp 1723858470
transform 1 0 14536 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_166
timestamp 1723858470
transform 1 0 15824 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_193
timestamp 1723858470
transform 1 0 18308 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_203
timestamp 1723858470
transform 1 0 19228 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_208
timestamp 1723858470
transform 1 0 19688 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_215
timestamp 1723858470
transform 1 0 20332 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_222
timestamp 1723858470
transform 1 0 20976 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_239
timestamp 1723858470
transform 1 0 22540 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_3
timestamp 1723858470
transform 1 0 828 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_64
timestamp 1723858470
transform 1 0 6440 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_81
timestamp 1723858470
transform 1 0 8004 0 -1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_94
timestamp 1723858470
transform 1 0 9200 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_106
timestamp 1723858470
transform 1 0 10304 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_113
timestamp 1723858470
transform 1 0 10948 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_136
timestamp 1723858470
transform 1 0 13064 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_144
timestamp 1723858470
transform 1 0 13800 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 1723858470
transform 1 0 15916 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_181
timestamp 1723858470
transform 1 0 17204 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_199
timestamp 1723858470
transform 1 0 18860 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_208
timestamp 1723858470
transform 1 0 19688 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_228
timestamp 1723858470
transform 1 0 21528 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_3
timestamp 1723858470
transform 1 0 828 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_9
timestamp 1723858470
transform 1 0 1380 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_13
timestamp 1723858470
transform 1 0 1748 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_23
timestamp 1723858470
transform 1 0 2668 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1723858470
transform 1 0 3036 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_29
timestamp 1723858470
transform 1 0 3220 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_40
timestamp 1723858470
transform 1 0 4232 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_68
timestamp 1723858470
transform 1 0 6808 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_79
timestamp 1723858470
transform 1 0 7820 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1723858470
transform 1 0 8188 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_85
timestamp 1723858470
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_90
timestamp 1723858470
transform 1 0 8832 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_96
timestamp 1723858470
transform 1 0 9384 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_107
timestamp 1723858470
transform 1 0 10396 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_129
timestamp 1723858470
transform 1 0 12420 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_133
timestamp 1723858470
transform 1 0 12788 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_137
timestamp 1723858470
transform 1 0 13156 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_141
timestamp 1723858470
transform 1 0 13524 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_145
timestamp 1723858470
transform 1 0 13892 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_162
timestamp 1723858470
transform 1 0 15456 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_174
timestamp 1723858470
transform 1 0 16560 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_186
timestamp 1723858470
transform 1 0 17664 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_194
timestamp 1723858470
transform 1 0 18400 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_207
timestamp 1723858470
transform 1 0 19596 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_213
timestamp 1723858470
transform 1 0 20148 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_225
timestamp 1723858470
transform 1 0 21252 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_242
timestamp 1723858470
transform 1 0 22816 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_17
timestamp 1723858470
transform 1 0 2116 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_29
timestamp 1723858470
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_45
timestamp 1723858470
transform 1 0 4692 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_53
timestamp 1723858470
transform 1 0 5428 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_78
timestamp 1723858470
transform 1 0 7728 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_89
timestamp 1723858470
transform 1 0 8740 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_93
timestamp 1723858470
transform 1 0 9108 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_125
timestamp 1723858470
transform 1 0 12052 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_150
timestamp 1723858470
transform 1 0 14352 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_161
timestamp 1723858470
transform 1 0 15364 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1723858470
transform 1 0 15916 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_194
timestamp 1723858470
transform 1 0 18400 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_202
timestamp 1723858470
transform 1 0 19136 0 -1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_208
timestamp 1723858470
transform 1 0 19688 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_220
timestamp 1723858470
transform 1 0 20792 0 -1 13600
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_225
timestamp 1723858470
transform 1 0 21252 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_237
timestamp 1723858470
transform 1 0 22356 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_29
timestamp 1723858470
transform 1 0 3220 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_33
timestamp 1723858470
transform 1 0 3588 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_39
timestamp 1723858470
transform 1 0 4140 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_51
timestamp 1723858470
transform 1 0 5244 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_60
timestamp 1723858470
transform 1 0 6072 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_103
timestamp 1723858470
transform 1 0 10028 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_124
timestamp 1723858470
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_147
timestamp 1723858470
transform 1 0 14076 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_163
timestamp 1723858470
transform 1 0 15548 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_167
timestamp 1723858470
transform 1 0 15916 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_180
timestamp 1723858470
transform 1 0 17112 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_224
timestamp 1723858470
transform 1 0 21160 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_241
timestamp 1723858470
transform 1 0 22724 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_3
timestamp 1723858470
transform 1 0 828 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_34
timestamp 1723858470
transform 1 0 3680 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_67
timestamp 1723858470
transform 1 0 6716 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_73
timestamp 1723858470
transform 1 0 7268 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_81
timestamp 1723858470
transform 1 0 8004 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_95
timestamp 1723858470
transform 1 0 9292 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_107
timestamp 1723858470
transform 1 0 10396 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1723858470
transform 1 0 10764 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_113
timestamp 1723858470
transform 1 0 10948 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_132
timestamp 1723858470
transform 1 0 12696 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_163
timestamp 1723858470
transform 1 0 15548 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1723858470
transform 1 0 15916 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 1723858470
transform 1 0 16100 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_181
timestamp 1723858470
transform 1 0 17204 0 -1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_189
timestamp 1723858470
transform 1 0 17940 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_217
timestamp 1723858470
transform 1 0 20516 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 1723858470
transform 1 0 21068 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_225
timestamp 1723858470
transform 1 0 21252 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_237
timestamp 1723858470
transform 1 0 22356 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_3
timestamp 1723858470
transform 1 0 828 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1723858470
transform 1 0 3036 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_29
timestamp 1723858470
transform 1 0 3220 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_80
timestamp 1723858470
transform 1 0 7912 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_94
timestamp 1723858470
transform 1 0 9200 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_108
timestamp 1723858470
transform 1 0 10488 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1723858470
transform 1 0 13340 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_149
timestamp 1723858470
transform 1 0 14260 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_163
timestamp 1723858470
transform 1 0 15548 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_185
timestamp 1723858470
transform 1 0 17572 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_193
timestamp 1723858470
transform 1 0 18308 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_219
timestamp 1723858470
transform 1 0 20700 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_225
timestamp 1723858470
transform 1 0 21252 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_233
timestamp 1723858470
transform 1 0 21988 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_241
timestamp 1723858470
transform 1 0 22724 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_3
timestamp 1723858470
transform 1 0 828 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_15
timestamp 1723858470
transform 1 0 1932 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_19
timestamp 1723858470
transform 1 0 2300 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_28
timestamp 1723858470
transform 1 0 3128 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_78
timestamp 1723858470
transform 1 0 7728 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_90
timestamp 1723858470
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1723858470
transform 1 0 10764 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_116
timestamp 1723858470
transform 1 0 11224 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_124
timestamp 1723858470
transform 1 0 11960 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_135
timestamp 1723858470
transform 1 0 12972 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_147
timestamp 1723858470
transform 1 0 14076 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_154
timestamp 1723858470
transform 1 0 14720 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1723858470
transform 1 0 15916 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_169
timestamp 1723858470
transform 1 0 16100 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_202
timestamp 1723858470
transform 1 0 19136 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_219
timestamp 1723858470
transform 1 0 20700 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_225
timestamp 1723858470
transform 1 0 21252 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_19
timestamp 1723858470
transform 1 0 2300 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_79
timestamp 1723858470
transform 1 0 7820 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_88
timestamp 1723858470
transform 1 0 8648 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_120
timestamp 1723858470
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1723858470
transform 1 0 13340 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_160
timestamp 1723858470
transform 1 0 15272 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_168
timestamp 1723858470
transform 1 0 16008 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_176
timestamp 1723858470
transform 1 0 16744 0 1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_182
timestamp 1723858470
transform 1 0 17296 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_194
timestamp 1723858470
transform 1 0 18400 0 1 15776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_197
timestamp 1723858470
transform 1 0 18676 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_215
timestamp 1723858470
transform 1 0 20332 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_223
timestamp 1723858470
transform 1 0 21068 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_235
timestamp 1723858470
transform 1 0 22172 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_3
timestamp 1723858470
transform 1 0 828 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_44
timestamp 1723858470
transform 1 0 4600 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_81
timestamp 1723858470
transform 1 0 8004 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_108
timestamp 1723858470
transform 1 0 10488 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_143
timestamp 1723858470
transform 1 0 13708 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_151
timestamp 1723858470
transform 1 0 14444 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_173
timestamp 1723858470
transform 1 0 16468 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_190
timestamp 1723858470
transform 1 0 18032 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_207
timestamp 1723858470
transform 1 0 19596 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_228
timestamp 1723858470
transform 1 0 21528 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_3
timestamp 1723858470
transform 1 0 828 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_9
timestamp 1723858470
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_19
timestamp 1723858470
transform 1 0 2300 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_56
timestamp 1723858470
transform 1 0 5704 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_69
timestamp 1723858470
transform 1 0 6900 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_79
timestamp 1723858470
transform 1 0 7820 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1723858470
transform 1 0 8188 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_95
timestamp 1723858470
transform 1 0 9292 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_101
timestamp 1723858470
transform 1 0 9844 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_108
timestamp 1723858470
transform 1 0 10488 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_112
timestamp 1723858470
transform 1 0 10856 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_141
timestamp 1723858470
transform 1 0 13524 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_170
timestamp 1723858470
transform 1 0 16192 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_174
timestamp 1723858470
transform 1 0 16560 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_180
timestamp 1723858470
transform 1 0 17112 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 1723858470
transform 1 0 18492 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_200
timestamp 1723858470
transform 1 0 18952 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_3
timestamp 1723858470
transform 1 0 828 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_48
timestamp 1723858470
transform 1 0 4968 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_155
timestamp 1723858470
transform 1 0 14812 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 1723858470
transform 1 0 15916 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_179
timestamp 1723858470
transform 1 0 17020 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_192
timestamp 1723858470
transform 1 0 18216 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_214
timestamp 1723858470
transform 1 0 20240 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_228
timestamp 1723858470
transform 1 0 21528 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_3
timestamp 1723858470
transform 1 0 828 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_11
timestamp 1723858470
transform 1 0 1564 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_17
timestamp 1723858470
transform 1 0 2116 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_29
timestamp 1723858470
transform 1 0 3220 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_46
timestamp 1723858470
transform 1 0 4784 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_53
timestamp 1723858470
transform 1 0 5428 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_62
timestamp 1723858470
transform 1 0 6256 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_94
timestamp 1723858470
transform 1 0 9200 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_102
timestamp 1723858470
transform 1 0 9936 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_108
timestamp 1723858470
transform 1 0 10488 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_112
timestamp 1723858470
transform 1 0 10856 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_118
timestamp 1723858470
transform 1 0 11408 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_146
timestamp 1723858470
transform 1 0 13984 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_151
timestamp 1723858470
transform 1 0 14444 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_159
timestamp 1723858470
transform 1 0 15180 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_167
timestamp 1723858470
transform 1 0 15916 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_3
timestamp 1723858470
transform 1 0 828 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_22
timestamp 1723858470
transform 1 0 2576 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1723858470
transform 1 0 5612 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_63
timestamp 1723858470
transform 1 0 6348 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_132
timestamp 1723858470
transform 1 0 12696 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_142
timestamp 1723858470
transform 1 0 13616 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_155
timestamp 1723858470
transform 1 0 14812 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_166
timestamp 1723858470
transform 1 0 15824 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_169
timestamp 1723858470
transform 1 0 16100 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_180
timestamp 1723858470
transform 1 0 17112 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_195
timestamp 1723858470
transform 1 0 18492 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_222
timestamp 1723858470
transform 1 0 20976 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_228
timestamp 1723858470
transform 1 0 21528 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_16
timestamp 1723858470
transform 1 0 2024 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_38
timestamp 1723858470
transform 1 0 4048 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_51
timestamp 1723858470
transform 1 0 5244 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_85
timestamp 1723858470
transform 1 0 8372 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_100
timestamp 1723858470
transform 1 0 9752 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_110
timestamp 1723858470
transform 1 0 10672 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_128
timestamp 1723858470
transform 1 0 12328 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_137
timestamp 1723858470
transform 1 0 13156 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_144
timestamp 1723858470
transform 1 0 13800 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_195
timestamp 1723858470
transform 1 0 18492 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_228
timestamp 1723858470
transform 1 0 21528 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_244
timestamp 1723858470
transform 1 0 23000 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_3
timestamp 1723858470
transform 1 0 828 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_27
timestamp 1723858470
transform 1 0 3036 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_52
timestamp 1723858470
transform 1 0 5336 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_75
timestamp 1723858470
transform 1 0 7452 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_81
timestamp 1723858470
transform 1 0 8004 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_88
timestamp 1723858470
transform 1 0 8648 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_211
timestamp 1723858470
transform 1 0 19964 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_228
timestamp 1723858470
transform 1 0 21528 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_3
timestamp 1723858470
transform 1 0 828 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_17
timestamp 1723858470
transform 1 0 2116 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_24
timestamp 1723858470
transform 1 0 2760 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_45
timestamp 1723858470
transform 1 0 4692 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_70
timestamp 1723858470
transform 1 0 6992 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_85
timestamp 1723858470
transform 1 0 8372 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_90
timestamp 1723858470
transform 1 0 8832 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_110
timestamp 1723858470
transform 1 0 10672 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_121
timestamp 1723858470
transform 1 0 11684 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_138
timestamp 1723858470
transform 1 0 13248 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_144
timestamp 1723858470
transform 1 0 13800 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_156
timestamp 1723858470
transform 1 0 14904 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_163
timestamp 1723858470
transform 1 0 15548 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_211
timestamp 1723858470
transform 1 0 19964 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_243
timestamp 1723858470
transform 1 0 22908 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_3
timestamp 1723858470
transform 1 0 828 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_27
timestamp 1723858470
transform 1 0 3036 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_31
timestamp 1723858470
transform 1 0 3404 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_83
timestamp 1723858470
transform 1 0 8188 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_95
timestamp 1723858470
transform 1 0 9292 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_104
timestamp 1723858470
transform 1 0 10120 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_152
timestamp 1723858470
transform 1 0 14536 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_195
timestamp 1723858470
transform 1 0 18492 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_19
timestamp 1723858470
transform 1 0 2300 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_39
timestamp 1723858470
transform 1 0 4140 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_51
timestamp 1723858470
transform 1 0 5244 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_64
timestamp 1723858470
transform 1 0 6440 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_78
timestamp 1723858470
transform 1 0 7728 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_98
timestamp 1723858470
transform 1 0 9568 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_106
timestamp 1723858470
transform 1 0 10304 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_115
timestamp 1723858470
transform 1 0 11132 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_124
timestamp 1723858470
transform 1 0 11960 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_134
timestamp 1723858470
transform 1 0 12880 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_141
timestamp 1723858470
transform 1 0 13524 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_224
timestamp 1723858470
transform 1 0 21160 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_3
timestamp 1723858470
transform 1 0 828 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_11
timestamp 1723858470
transform 1 0 1564 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_23
timestamp 1723858470
transform 1 0 2668 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_31
timestamp 1723858470
transform 1 0 3404 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_50
timestamp 1723858470
transform 1 0 5152 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 1723858470
transform 1 0 5612 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_64
timestamp 1723858470
transform 1 0 6440 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_113
timestamp 1723858470
transform 1 0 10948 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_119
timestamp 1723858470
transform 1 0 11500 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_127
timestamp 1723858470
transform 1 0 12236 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_132
timestamp 1723858470
transform 1 0 12696 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_167
timestamp 1723858470
transform 1 0 15916 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_172
timestamp 1723858470
transform 1 0 16376 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_3
timestamp 1723858470
transform 1 0 828 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_9
timestamp 1723858470
transform 1 0 1380 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1723858470
transform 1 0 3036 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_29
timestamp 1723858470
transform 1 0 3220 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_138
timestamp 1723858470
transform 1 0 13248 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_152
timestamp 1723858470
transform 1 0 14536 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_226
timestamp 1723858470
transform 1 0 21344 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_244
timestamp 1723858470
transform 1 0 23000 0 1 22304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 1723858470
transform 1 0 828 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_15
timestamp 1723858470
transform 1 0 1932 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_21
timestamp 1723858470
transform 1 0 2484 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_27
timestamp 1723858470
transform 1 0 3036 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_49
timestamp 1723858470
transform 1 0 5060 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 1723858470
transform 1 0 5612 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_60
timestamp 1723858470
transform 1 0 6072 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_85
timestamp 1723858470
transform 1 0 8372 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_103
timestamp 1723858470
transform 1 0 10028 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_169
timestamp 1723858470
transform 1 0 16100 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_190
timestamp 1723858470
transform 1 0 18032 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_213
timestamp 1723858470
transform 1 0 20148 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 8280 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1723858470
transform -1 0 18584 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1723858470
transform 1 0 13800 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1723858470
transform -1 0 8464 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1723858470
transform -1 0 23092 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1723858470
transform -1 0 23000 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1723858470
transform -1 0 23092 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1723858470
transform -1 0 21620 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1723858470
transform 1 0 20240 0 -1 23392
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1723858470
transform 1 0 18216 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1723858470
transform -1 0 21344 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1723858470
transform 1 0 18216 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1723858470
transform -1 0 16560 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 9660 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1723858470
transform 1 0 11592 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1723858470
transform -1 0 5704 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1723858470
transform -1 0 4968 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1723858470
transform -1 0 4232 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1723858470
transform -1 0 3128 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1723858470
transform 1 0 2760 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 1723858470
transform 1 0 2300 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 1723858470
transform -1 0 1656 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 1723858470
transform 1 0 828 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 1723858470
transform -1 0 5336 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1723858470
transform -1 0 4600 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1723858470
transform -1 0 3864 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1723858470
transform -1 0 2760 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1723858470
transform -1 0 2392 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1723858470
transform -1 0 2024 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1723858470
transform -1 0 1288 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1723858470
transform -1 0 1564 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1723858470
transform 1 0 10120 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1723858470
transform 1 0 12880 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1723858470
transform -1 0 15732 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1723858470
transform 1 0 14628 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1723858470
transform -1 0 13892 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1723858470
transform 1 0 12604 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1723858470
transform 1 0 11868 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1723858470
transform 1 0 10120 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1723858470
transform 1 0 9384 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1723858470
transform 1 0 8648 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1723858470
transform -1 0 15364 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1723858470
transform -1 0 14260 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1723858470
transform -1 0 13340 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1723858470
transform -1 0 12604 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1723858470
transform -1 0 10856 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1723858470
transform 1 0 9752 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 1723858470
transform 1 0 9016 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 1723858470
transform 1 0 9292 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1723858470
transform 1 0 7912 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1723858470
transform 1 0 9292 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1723858470
transform -1 0 10856 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1723858470
transform -1 0 13616 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1723858470
transform -1 0 22724 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1723858470
transform 1 0 22724 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1723858470
transform 1 0 22632 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1723858470
transform 1 0 22356 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1723858470
transform 1 0 21620 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1723858470
transform 1 0 20700 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1723858470
transform 1 0 19412 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1723858470
transform 1 0 18676 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1723858470
transform -1 0 21160 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1723858470
transform -1 0 22264 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1723858470
transform 1 0 22724 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1723858470
transform 1 0 21988 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1723858470
transform 1 0 21252 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1723858470
transform 1 0 20332 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1723858470
transform 1 0 19044 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1723858470
transform 1 0 18124 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1723858470
transform -1 0 9292 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1723858470
transform 1 0 11224 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_42
timestamp 1723858470
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1723858470
transform -1 0 23368 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_43
timestamp 1723858470
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1723858470
transform -1 0 23368 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_44
timestamp 1723858470
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1723858470
transform -1 0 23368 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_45
timestamp 1723858470
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1723858470
transform -1 0 23368 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_46
timestamp 1723858470
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1723858470
transform -1 0 23368 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_47
timestamp 1723858470
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1723858470
transform -1 0 23368 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_48
timestamp 1723858470
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1723858470
transform -1 0 23368 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_49
timestamp 1723858470
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1723858470
transform -1 0 23368 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_50
timestamp 1723858470
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1723858470
transform -1 0 23368 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_51
timestamp 1723858470
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1723858470
transform -1 0 23368 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_52
timestamp 1723858470
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1723858470
transform -1 0 23368 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_53
timestamp 1723858470
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1723858470
transform -1 0 23368 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_54
timestamp 1723858470
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1723858470
transform -1 0 23368 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_55
timestamp 1723858470
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1723858470
transform -1 0 23368 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_56
timestamp 1723858470
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1723858470
transform -1 0 23368 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_57
timestamp 1723858470
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1723858470
transform -1 0 23368 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_58
timestamp 1723858470
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1723858470
transform -1 0 23368 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_59
timestamp 1723858470
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1723858470
transform -1 0 23368 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_60
timestamp 1723858470
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1723858470
transform -1 0 23368 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_61
timestamp 1723858470
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1723858470
transform -1 0 23368 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_62
timestamp 1723858470
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1723858470
transform -1 0 23368 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_63
timestamp 1723858470
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1723858470
transform -1 0 23368 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_64
timestamp 1723858470
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1723858470
transform -1 0 23368 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_65
timestamp 1723858470
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1723858470
transform -1 0 23368 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_66
timestamp 1723858470
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1723858470
transform -1 0 23368 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_67
timestamp 1723858470
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1723858470
transform -1 0 23368 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_68
timestamp 1723858470
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1723858470
transform -1 0 23368 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_69
timestamp 1723858470
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1723858470
transform -1 0 23368 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_70
timestamp 1723858470
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1723858470
transform -1 0 23368 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_71
timestamp 1723858470
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1723858470
transform -1 0 23368 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_72
timestamp 1723858470
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1723858470
transform -1 0 23368 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_73
timestamp 1723858470
transform 1 0 552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1723858470
transform -1 0 23368 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_74
timestamp 1723858470
transform 1 0 552 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1723858470
transform -1 0 23368 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_75
timestamp 1723858470
transform 1 0 552 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1723858470
transform -1 0 23368 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_76
timestamp 1723858470
transform 1 0 552 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1723858470
transform -1 0 23368 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_77
timestamp 1723858470
transform 1 0 552 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1723858470
transform -1 0 23368 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_78
timestamp 1723858470
transform 1 0 552 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1723858470
transform -1 0 23368 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_79
timestamp 1723858470
transform 1 0 552 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1723858470
transform -1 0 23368 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_80
timestamp 1723858470
transform 1 0 552 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1723858470
transform -1 0 23368 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_81
timestamp 1723858470
transform 1 0 552 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 1723858470
transform -1 0 23368 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_82
timestamp 1723858470
transform 1 0 552 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 1723858470
transform -1 0 23368 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_83
timestamp 1723858470
transform 1 0 552 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 1723858470
transform -1 0 23368 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_84 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_85
timestamp 1723858470
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_86
timestamp 1723858470
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_87
timestamp 1723858470
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_88
timestamp 1723858470
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_89
timestamp 1723858470
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_90
timestamp 1723858470
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_91
timestamp 1723858470
transform 1 0 21160 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_92
timestamp 1723858470
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_93
timestamp 1723858470
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_94
timestamp 1723858470
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_95
timestamp 1723858470
transform 1 0 21160 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_96
timestamp 1723858470
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_97
timestamp 1723858470
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_98
timestamp 1723858470
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_99
timestamp 1723858470
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_100
timestamp 1723858470
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_101
timestamp 1723858470
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_102
timestamp 1723858470
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_103
timestamp 1723858470
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_104
timestamp 1723858470
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_105
timestamp 1723858470
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_106
timestamp 1723858470
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_107
timestamp 1723858470
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_108
timestamp 1723858470
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_109
timestamp 1723858470
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_110
timestamp 1723858470
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_111
timestamp 1723858470
transform 1 0 21160 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_112
timestamp 1723858470
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_113
timestamp 1723858470
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_114
timestamp 1723858470
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_115
timestamp 1723858470
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_116
timestamp 1723858470
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_117
timestamp 1723858470
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_118
timestamp 1723858470
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_119
timestamp 1723858470
transform 1 0 21160 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_120
timestamp 1723858470
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_121
timestamp 1723858470
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_122
timestamp 1723858470
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_123
timestamp 1723858470
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_124
timestamp 1723858470
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_125
timestamp 1723858470
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_126
timestamp 1723858470
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_127
timestamp 1723858470
transform 1 0 21160 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_128
timestamp 1723858470
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_129
timestamp 1723858470
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_130
timestamp 1723858470
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_131
timestamp 1723858470
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_132
timestamp 1723858470
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_133
timestamp 1723858470
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_134
timestamp 1723858470
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_135
timestamp 1723858470
transform 1 0 21160 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_136
timestamp 1723858470
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_137
timestamp 1723858470
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_138
timestamp 1723858470
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_139
timestamp 1723858470
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_140
timestamp 1723858470
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_141
timestamp 1723858470
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_142
timestamp 1723858470
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_143
timestamp 1723858470
transform 1 0 21160 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_144
timestamp 1723858470
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_145
timestamp 1723858470
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_146
timestamp 1723858470
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_147
timestamp 1723858470
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_148
timestamp 1723858470
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_149
timestamp 1723858470
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_150
timestamp 1723858470
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_151
timestamp 1723858470
transform 1 0 21160 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_152
timestamp 1723858470
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_153
timestamp 1723858470
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_154
timestamp 1723858470
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_155
timestamp 1723858470
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_156
timestamp 1723858470
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_157
timestamp 1723858470
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_158
timestamp 1723858470
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_159
timestamp 1723858470
transform 1 0 21160 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_160
timestamp 1723858470
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_161
timestamp 1723858470
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_162
timestamp 1723858470
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_163
timestamp 1723858470
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_164
timestamp 1723858470
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_165
timestamp 1723858470
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_166
timestamp 1723858470
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_167
timestamp 1723858470
transform 1 0 21160 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_168
timestamp 1723858470
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_169
timestamp 1723858470
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_170
timestamp 1723858470
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_171
timestamp 1723858470
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_172
timestamp 1723858470
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_173
timestamp 1723858470
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_174
timestamp 1723858470
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_175
timestamp 1723858470
transform 1 0 21160 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_176
timestamp 1723858470
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_177
timestamp 1723858470
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_178
timestamp 1723858470
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_179
timestamp 1723858470
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_180
timestamp 1723858470
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_181
timestamp 1723858470
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_182
timestamp 1723858470
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_183
timestamp 1723858470
transform 1 0 21160 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_184
timestamp 1723858470
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_185
timestamp 1723858470
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_186
timestamp 1723858470
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_187
timestamp 1723858470
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_188
timestamp 1723858470
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_189
timestamp 1723858470
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_190
timestamp 1723858470
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_191
timestamp 1723858470
transform 1 0 21160 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_192
timestamp 1723858470
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_193
timestamp 1723858470
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_194
timestamp 1723858470
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_195
timestamp 1723858470
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_196
timestamp 1723858470
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_197
timestamp 1723858470
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_198
timestamp 1723858470
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_199
timestamp 1723858470
transform 1 0 21160 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_200
timestamp 1723858470
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_201
timestamp 1723858470
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_202
timestamp 1723858470
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_203
timestamp 1723858470
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_204
timestamp 1723858470
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_205
timestamp 1723858470
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_206
timestamp 1723858470
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_207
timestamp 1723858470
transform 1 0 21160 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_208
timestamp 1723858470
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_209
timestamp 1723858470
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_210
timestamp 1723858470
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_211
timestamp 1723858470
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_212
timestamp 1723858470
transform 1 0 5704 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_213
timestamp 1723858470
transform 1 0 10856 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_214
timestamp 1723858470
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_215
timestamp 1723858470
transform 1 0 21160 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_216
timestamp 1723858470
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_217
timestamp 1723858470
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_218
timestamp 1723858470
transform 1 0 13432 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_219
timestamp 1723858470
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_220
timestamp 1723858470
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_221
timestamp 1723858470
transform 1 0 10856 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_222
timestamp 1723858470
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_223
timestamp 1723858470
transform 1 0 21160 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_224
timestamp 1723858470
transform 1 0 3128 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_225
timestamp 1723858470
transform 1 0 8280 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_226
timestamp 1723858470
transform 1 0 13432 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_227
timestamp 1723858470
transform 1 0 18584 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_228
timestamp 1723858470
transform 1 0 5704 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_229
timestamp 1723858470
transform 1 0 10856 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_230
timestamp 1723858470
transform 1 0 16008 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_231
timestamp 1723858470
transform 1 0 21160 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_232
timestamp 1723858470
transform 1 0 3128 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_233
timestamp 1723858470
transform 1 0 8280 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_234
timestamp 1723858470
transform 1 0 13432 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_235
timestamp 1723858470
transform 1 0 18584 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_236
timestamp 1723858470
transform 1 0 5704 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_237
timestamp 1723858470
transform 1 0 10856 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_238
timestamp 1723858470
transform 1 0 16008 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_239
timestamp 1723858470
transform 1 0 21160 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_240
timestamp 1723858470
transform 1 0 3128 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_241
timestamp 1723858470
transform 1 0 8280 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_242
timestamp 1723858470
transform 1 0 13432 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_243
timestamp 1723858470
transform 1 0 18584 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_244
timestamp 1723858470
transform 1 0 5704 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_245
timestamp 1723858470
transform 1 0 10856 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_246
timestamp 1723858470
transform 1 0 16008 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_247
timestamp 1723858470
transform 1 0 21160 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_248
timestamp 1723858470
transform 1 0 3128 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_249
timestamp 1723858470
transform 1 0 8280 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_250
timestamp 1723858470
transform 1 0 13432 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_251
timestamp 1723858470
transform 1 0 18584 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_252
timestamp 1723858470
transform 1 0 3128 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_253
timestamp 1723858470
transform 1 0 5704 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_254
timestamp 1723858470
transform 1 0 8280 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_255
timestamp 1723858470
transform 1 0 10856 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_256
timestamp 1723858470
transform 1 0 13432 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_257
timestamp 1723858470
transform 1 0 16008 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_258
timestamp 1723858470
transform 1 0 18584 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_259
timestamp 1723858470
transform 1 0 21160 0 -1 23392
box -38 -48 130 592
<< labels >>
rlabel metal1 s 11960 23392 11960 23392 4 VGND
rlabel metal1 s 11960 22848 11960 22848 4 VPWR
rlabel metal1 s 21666 19414 21666 19414 4 _0000_
rlabel metal1 s 22908 16218 22908 16218 4 _0001_
rlabel metal2 s 21390 20196 21390 20196 4 _0002_
rlabel metal1 s 21298 18938 21298 18938 4 _0003_
rlabel metal1 s 21114 21462 21114 21462 4 _0004_
rlabel metal1 s 20792 22134 20792 22134 4 _0005_
rlabel metal1 s 21436 21590 21436 21590 4 _0006_
rlabel metal1 s 21252 22678 21252 22678 4 _0007_
rlabel metal1 s 21160 21114 21160 21114 4 _0008_
rlabel metal1 s 23000 18054 23000 18054 4 _0009_
rlabel metal2 s 22310 20978 22310 20978 4 _0010_
rlabel metal2 s 23000 20876 23000 20876 4 _0011_
rlabel metal1 s 10948 17306 10948 17306 4 _0012_
rlabel metal1 s 12082 18122 12082 18122 4 _0013_
rlabel metal2 s 9701 17714 9701 17714 4 _0014_
rlabel metal2 s 9333 16626 9333 16626 4 _0015_
rlabel metal1 s 6016 16626 6016 16626 4 _0016_
rlabel metal2 s 1145 16014 1145 16014 4 _0017_
rlabel metal1 s 1426 17306 1426 17306 4 _0018_
rlabel metal2 s 3077 17714 3077 17714 4 _0019_
rlabel metal1 s 3440 16014 3440 16014 4 _0020_
rlabel metal1 s 2203 16694 2203 16694 4 _0021_
rlabel metal1 s 18722 18938 18722 18938 4 _0022_
rlabel metal1 s 19131 17782 19131 17782 4 _0023_
rlabel metal2 s 15778 19074 15778 19074 4 _0024_
rlabel metal2 s 14945 19210 14945 19210 4 _0025_
rlabel metal1 s 13800 19482 13800 19482 4 _0026_
rlabel metal1 s 12604 18938 12604 18938 4 _0027_
rlabel metal1 s 10488 18394 10488 18394 4 _0028_
rlabel metal1 s 2387 12342 2387 12342 4 _0029_
rlabel metal2 s 1242 10880 1242 10880 4 _0030_
rlabel metal2 s 1150 9622 1150 9622 4 _0031_
rlabel metal1 s 1743 13838 1743 13838 4 _0032_
rlabel metal2 s 3450 14722 3450 14722 4 _0033_
rlabel metal1 s 17046 21420 17046 21420 4 _0034_
rlabel metal1 s 16514 20570 16514 20570 4 _0035_
rlabel metal1 s 15210 22474 15210 22474 4 _0036_
rlabel metal1 s 15640 22202 15640 22202 4 _0037_
rlabel metal1 s 14720 21590 14720 21590 4 _0038_
rlabel metal2 s 18630 21556 18630 21556 4 _0039_
rlabel metal1 s 16284 22202 16284 22202 4 _0040_
rlabel metal1 s 18461 20298 18461 20298 4 _0041_
rlabel metal1 s 7171 19210 7171 19210 4 _0042_
rlabel metal1 s 13432 20570 13432 20570 4 _0043_
rlabel metal2 s 12093 20298 12093 20298 4 _0044_
rlabel metal1 s 12180 23154 12180 23154 4 _0045_
rlabel metal1 s 10442 20570 10442 20570 4 _0046_
rlabel metal2 s 9246 22950 9246 22950 4 _0047_
rlabel metal1 s 3128 22202 3128 22202 4 _0048_
rlabel metal2 s 1982 21454 1982 21454 4 _0049_
rlabel metal2 s 2622 20808 2622 20808 4 _0050_
rlabel metal1 s 3164 18802 3164 18802 4 _0051_
rlabel metal1 s 3496 19482 3496 19482 4 _0052_
rlabel metal1 s 6716 22746 6716 22746 4 _0053_
rlabel metal2 s 22862 17952 22862 17952 4 _0054_
rlabel metal2 s 21569 22066 21569 22066 4 _0055_
rlabel metal2 s 22218 11390 22218 11390 4 _0056_
rlabel metal1 s 22167 16626 22167 16626 4 _0057_
rlabel metal1 s 22264 16150 22264 16150 4 _0058_
rlabel metal2 s 22218 16932 22218 16932 4 _0059_
rlabel metal1 s 21712 11866 21712 11866 4 _0060_
rlabel metal1 s 21558 12682 21558 12682 4 _0061_
rlabel metal1 s 19867 18190 19867 18190 4 _0062_
rlabel metal1 s 9154 19176 9154 19176 4 _0063_
rlabel metal1 s 18446 6800 18446 6800 4 _0064_
rlabel metal2 s 22126 4250 22126 4250 4 _0065_
rlabel metal1 s 22908 2482 22908 2482 4 _0066_
rlabel metal1 s 22540 2074 22540 2074 4 _0067_
rlabel metal1 s 14076 17306 14076 17306 4 _0068_
rlabel metal1 s 14260 17850 14260 17850 4 _0069_
rlabel metal1 s 14122 17680 14122 17680 4 _0070_
rlabel metal1 s 15732 17306 15732 17306 4 _0071_
rlabel metal1 s 14030 17612 14030 17612 4 _0072_
rlabel metal1 s 15686 12240 15686 12240 4 _0073_
rlabel metal2 s 14398 14212 14398 14212 4 _0074_
rlabel metal1 s 13800 14926 13800 14926 4 _0075_
rlabel metal1 s 14444 14450 14444 14450 4 _0076_
rlabel metal1 s 17618 15470 17618 15470 4 _0077_
rlabel metal1 s 14766 14348 14766 14348 4 _0078_
rlabel metal1 s 14950 14246 14950 14246 4 _0079_
rlabel metal2 s 15502 11900 15502 11900 4 _0080_
rlabel metal2 s 15594 11679 15594 11679 4 _0081_
rlabel metal1 s 15686 11526 15686 11526 4 _0082_
rlabel metal1 s 15318 9010 15318 9010 4 _0083_
rlabel metal1 s 14214 8976 14214 8976 4 _0084_
rlabel metal2 s 16882 8602 16882 8602 4 _0085_
rlabel metal2 s 17618 6732 17618 6732 4 _0086_
rlabel metal1 s 18676 4794 18676 4794 4 _0087_
rlabel metal1 s 16790 5236 16790 5236 4 _0088_
rlabel metal2 s 19090 5270 19090 5270 4 _0089_
rlabel metal1 s 19228 4998 19228 4998 4 _0090_
rlabel metal2 s 20930 748 20930 748 4 _0091_
rlabel metal3 s 10626 16643 10626 16643 4 _0092_
rlabel metal1 s 10856 16218 10856 16218 4 _0093_
rlabel metal1 s 12098 16660 12098 16660 4 _0094_
rlabel metal2 s 12006 17102 12006 17102 4 _0095_
rlabel metal1 s 11592 11186 11592 11186 4 _0096_
rlabel metal2 s 12742 14025 12742 14025 4 _0097_
rlabel metal1 s 4094 13294 4094 13294 4 _0098_
rlabel metal1 s 5014 13226 5014 13226 4 _0099_
rlabel metal1 s 11408 11322 11408 11322 4 _0100_
rlabel metal2 s 11086 11356 11086 11356 4 _0101_
rlabel metal2 s 15594 6919 15594 6919 4 _0102_
rlabel metal2 s 16054 8602 16054 8602 4 _0103_
rlabel metal2 s 16790 7548 16790 7548 4 _0104_
rlabel metal3 s 16330 4131 16330 4131 4 _0105_
rlabel metal2 s 16422 4199 16422 4199 4 _0106_
rlabel metal1 s 16514 2516 16514 2516 4 _0107_
rlabel metal1 s 18400 2074 18400 2074 4 _0108_
rlabel metal2 s 3450 11968 3450 11968 4 _0109_
rlabel metal1 s 3588 12614 3588 12614 4 _0110_
rlabel metal1 s 4094 11662 4094 11662 4 _0111_
rlabel metal3 s 11477 15300 11477 15300 4 _0112_
rlabel metal2 s 4324 10574 4324 10574 4 _0113_
rlabel metal1 s 3082 11220 3082 11220 4 _0114_
rlabel metal1 s 3312 10982 3312 10982 4 _0115_
rlabel metal2 s 3634 10404 3634 10404 4 _0116_
rlabel metal2 s 3910 13226 3910 13226 4 _0117_
rlabel metal1 s 3542 12682 3542 12682 4 _0118_
rlabel metal1 s 4278 10676 4278 10676 4 _0119_
rlabel metal2 s 10902 10506 10902 10506 4 _0120_
rlabel metal1 s 13938 10744 13938 10744 4 _0121_
rlabel metal2 s 13846 8636 13846 8636 4 _0122_
rlabel metal1 s 14582 7344 14582 7344 4 _0123_
rlabel metal1 s 14398 6664 14398 6664 4 _0124_
rlabel metal2 s 14214 7004 14214 7004 4 _0125_
rlabel metal1 s 14628 2482 14628 2482 4 _0126_
rlabel metal1 s 15594 2448 15594 2448 4 _0127_
rlabel metal2 s 20102 2227 20102 2227 4 _0128_
rlabel metal1 s 8096 782 8096 782 4 _0129_
rlabel metal1 s 3036 4794 3036 4794 4 _0130_
rlabel metal1 s 2484 4658 2484 4658 4 _0131_
rlabel metal1 s 2438 4012 2438 4012 4 _0132_
rlabel metal1 s 2300 4114 2300 4114 4 _0133_
rlabel metal2 s 3174 3740 3174 3740 4 _0134_
rlabel metal1 s 1610 4658 1610 4658 4 _0135_
rlabel metal2 s 1334 4828 1334 4828 4 _0136_
rlabel metal2 s 1150 4012 1150 4012 4 _0137_
rlabel metal2 s 1702 3910 1702 3910 4 _0138_
rlabel metal2 s 3082 3842 3082 3842 4 _0139_
rlabel metal1 s 7130 3638 7130 3638 4 _0140_
rlabel metal1 s 7774 3706 7774 3706 4 _0141_
rlabel metal1 s 8602 5270 8602 5270 4 _0142_
rlabel metal1 s 10212 9486 10212 9486 4 _0143_
rlabel metal1 s 9936 5202 9936 5202 4 _0144_
rlabel metal1 s 10166 5338 10166 5338 4 _0145_
rlabel metal1 s 11132 3570 11132 3570 4 _0146_
rlabel metal2 s 10810 3332 10810 3332 4 _0147_
rlabel metal1 s 10534 1870 10534 1870 4 _0148_
rlabel metal1 s 19872 918 19872 918 4 _0149_
rlabel metal2 s 2714 5814 2714 5814 4 _0150_
rlabel metal2 s 2530 7718 2530 7718 4 _0151_
rlabel metal2 s 2806 6715 2806 6715 4 _0152_
rlabel metal2 s 2806 7990 2806 7990 4 _0153_
rlabel metal1 s 4278 6800 4278 6800 4 _0154_
rlabel metal1 s 1610 6970 1610 6970 4 _0155_
rlabel metal1 s 1150 7208 1150 7208 4 _0156_
rlabel metal1 s 1242 6800 1242 6800 4 _0157_
rlabel metal2 s 1150 5780 1150 5780 4 _0158_
rlabel metal1 s 2162 6664 2162 6664 4 _0159_
rlabel metal2 s 4830 7004 4830 7004 4 _0160_
rlabel metal1 s 4784 6630 4784 6630 4 _0161_
rlabel metal1 s 6302 6902 6302 6902 4 _0162_
rlabel metal1 s 10304 5542 10304 5542 4 _0163_
rlabel metal1 s 10856 7922 10856 7922 4 _0164_
rlabel metal1 s 11040 5202 11040 5202 4 _0165_
rlabel metal2 s 10442 5542 10442 5542 4 _0166_
rlabel metal1 s 12098 4012 12098 4012 4 _0167_
rlabel metal1 s 11822 4114 11822 4114 4 _0168_
rlabel metal1 s 12328 2482 12328 2482 4 _0169_
rlabel metal2 s 20102 646 20102 646 4 _0170_
rlabel metal1 s 2300 8058 2300 8058 4 _0171_
rlabel metal1 s 2392 13294 2392 13294 4 _0172_
rlabel metal1 s 2162 8500 2162 8500 4 _0173_
rlabel metal1 s 2691 8534 2691 8534 4 _0174_
rlabel metal1 s 6808 7854 6808 7854 4 _0175_
rlabel metal1 s 13018 4488 13018 4488 4 _0176_
rlabel metal1 s 12328 6834 12328 6834 4 _0177_
rlabel metal2 s 14122 5916 14122 5916 4 _0178_
rlabel metal2 s 13018 4828 13018 4828 4 _0179_
rlabel metal1 s 13616 3502 13616 3502 4 _0180_
rlabel metal2 s 13846 3740 13846 3740 4 _0181_
rlabel metal1 s 13754 3366 13754 3366 4 _0182_
rlabel metal1 s 15962 2006 15962 2006 4 _0183_
rlabel metal2 s 1058 14110 1058 14110 4 _0184_
rlabel metal1 s 2990 13430 2990 13430 4 _0185_
rlabel metal2 s 2990 14246 2990 14246 4 _0186_
rlabel metal2 s 2898 14688 2898 14688 4 _0187_
rlabel metal1 s 3220 14246 3220 14246 4 _0188_
rlabel metal1 s 3128 14314 3128 14314 4 _0189_
rlabel metal1 s 2484 9010 2484 9010 4 _0190_
rlabel metal2 s 2990 9452 2990 9452 4 _0191_
rlabel metal2 s 3082 9180 3082 9180 4 _0192_
rlabel metal1 s 2599 8874 2599 8874 4 _0193_
rlabel metal2 s 3542 8704 3542 8704 4 _0194_
rlabel metal1 s 3727 8466 3727 8466 4 _0195_
rlabel metal3 s 8142 5661 8142 5661 4 _0196_
rlabel metal1 s 2898 16082 2898 16082 4 _0197_
rlabel metal1 s 7130 15878 7130 15878 4 _0198_
rlabel metal2 s 7912 7922 7912 7922 4 _0199_
rlabel metal2 s 8234 6732 8234 6732 4 _0200_
rlabel metal1 s 9522 8296 9522 8296 4 _0201_
rlabel metal2 s 9430 6732 9430 6732 4 _0202_
rlabel metal1 s 9706 5780 9706 5780 4 _0203_
rlabel metal1 s 7958 5610 7958 5610 4 _0204_
rlabel metal3 s 10534 3587 10534 3587 4 _0205_
rlabel metal1 s 10304 3570 10304 3570 4 _0206_
rlabel metal1 s 9890 3434 9890 3434 4 _0207_
rlabel metal1 s 10534 1258 10534 1258 4 _0208_
rlabel metal3 s 19366 1717 19366 1717 4 _0209_
rlabel metal1 s 22632 18190 22632 18190 4 _0210_
rlabel metal1 s 18262 19720 18262 19720 4 _0211_
rlabel metal2 s 9982 19040 9982 19040 4 _0212_
rlabel metal1 s 16146 19924 16146 19924 4 _0213_
rlabel metal1 s 8188 19346 8188 19346 4 _0214_
rlabel metal2 s 12466 17340 12466 17340 4 _0215_
rlabel metal1 s 8832 19482 8832 19482 4 _0216_
rlabel metal1 s 4784 17714 4784 17714 4 _0217_
rlabel metal2 s 3910 17204 3910 17204 4 _0218_
rlabel metal1 s 7084 18666 7084 18666 4 _0219_
rlabel metal1 s 8464 18394 8464 18394 4 _0220_
rlabel metal1 s 13570 19346 13570 19346 4 _0221_
rlabel metal2 s 9798 20128 9798 20128 4 _0222_
rlabel metal1 s 8924 18802 8924 18802 4 _0223_
rlabel metal1 s 10258 17204 10258 17204 4 _0224_
rlabel metal1 s 10626 17136 10626 17136 4 _0225_
rlabel metal2 s 20470 19890 20470 19890 4 _0226_
rlabel metal1 s 10534 20978 10534 20978 4 _0227_
rlabel metal1 s 11638 17306 11638 17306 4 _0228_
rlabel metal2 s 9614 17714 9614 17714 4 _0229_
rlabel metal2 s 9798 17646 9798 17646 4 _0230_
rlabel metal1 s 6210 17714 6210 17714 4 _0231_
rlabel metal2 s 8786 16592 8786 16592 4 _0232_
rlabel metal1 s 9016 17102 9016 17102 4 _0233_
rlabel metal1 s 5980 17850 5980 17850 4 _0234_
rlabel metal2 s 6394 17986 6394 17986 4 _0235_
rlabel metal1 s 8464 16558 8464 16558 4 _0236_
rlabel metal1 s 5762 17578 5762 17578 4 _0237_
rlabel metal1 s 5428 17510 5428 17510 4 _0238_
rlabel metal1 s 1334 17136 1334 17136 4 _0239_
rlabel metal1 s 6440 17238 6440 17238 4 _0240_
rlabel metal1 s 2392 17306 2392 17306 4 _0241_
rlabel metal2 s 10442 20298 10442 20298 4 _0242_
rlabel metal1 s 1656 17102 1656 17102 4 _0243_
rlabel metal1 s 2760 17306 2760 17306 4 _0244_
rlabel metal2 s 2714 17986 2714 17986 4 _0245_
rlabel metal1 s 2599 15606 2599 15606 4 _0246_
rlabel metal1 s 2576 16626 2576 16626 4 _0247_
rlabel metal1 s 2990 15470 2990 15470 4 _0248_
rlabel metal1 s 12098 20944 12098 20944 4 _0249_
rlabel metal1 s 10695 20774 10695 20774 4 _0250_
rlabel metal2 s 6210 20162 6210 20162 4 _0251_
rlabel metal1 s 6946 19788 6946 19788 4 _0252_
rlabel metal2 s 9798 20740 9798 20740 4 _0253_
rlabel metal1 s 8556 20230 8556 20230 4 _0254_
rlabel metal1 s 6486 20026 6486 20026 4 _0255_
rlabel metal2 s 5842 20502 5842 20502 4 _0256_
rlabel metal3 s 14628 20264 14628 20264 4 _0257_
rlabel metal1 s 16803 20026 16803 20026 4 _0258_
rlabel metal2 s 17618 19244 17618 19244 4 _0259_
rlabel metal1 s 17664 18938 17664 18938 4 _0260_
rlabel metal1 s 17618 19244 17618 19244 4 _0261_
rlabel metal2 s 1242 15793 1242 15793 4 _0262_
rlabel metal1 s 16514 19890 16514 19890 4 _0263_
rlabel metal2 s 17986 19584 17986 19584 4 _0264_
rlabel metal1 s 18216 18802 18216 18802 4 _0265_
rlabel metal1 s 17480 18258 17480 18258 4 _0266_
rlabel metal1 s 18308 18122 18308 18122 4 _0267_
rlabel metal1 s 19044 18190 19044 18190 4 _0268_
rlabel metal1 s 15180 18666 15180 18666 4 _0269_
rlabel metal1 s 12880 19482 12880 19482 4 _0270_
rlabel metal1 s 16054 18394 16054 18394 4 _0271_
rlabel metal1 s 15548 18802 15548 18802 4 _0272_
rlabel metal1 s 13984 18938 13984 18938 4 _0273_
rlabel metal2 s 14398 19040 14398 19040 4 _0274_
rlabel metal1 s 14720 19482 14720 19482 4 _0275_
rlabel metal1 s 11822 18258 11822 18258 4 _0276_
rlabel metal2 s 11822 19618 11822 19618 4 _0277_
rlabel metal2 s 12926 19040 12926 19040 4 _0278_
rlabel metal1 s 13570 19210 13570 19210 4 _0279_
rlabel metal1 s 11776 19482 11776 19482 4 _0280_
rlabel metal2 s 12106 19210 12106 19210 4 _0281_
rlabel metal2 s 12466 18972 12466 18972 4 _0282_
rlabel metal1 s 11454 18054 11454 18054 4 _0283_
rlabel metal1 s 11408 18870 11408 18870 4 _0284_
rlabel metal1 s 10350 18190 10350 18190 4 _0285_
rlabel metal2 s 1058 12733 1058 12733 4 _0286_
rlabel metal2 s 2024 15708 2024 15708 4 _0287_
rlabel metal1 s 1886 12410 1886 12410 4 _0288_
rlabel metal1 s 2346 12750 2346 12750 4 _0289_
rlabel metal1 s 2116 11662 2116 11662 4 _0290_
rlabel metal1 s 1794 11866 1794 11866 4 _0291_
rlabel metal1 s 1242 10710 1242 10710 4 _0292_
rlabel metal1 s 1012 10574 1012 10574 4 _0293_
rlabel metal1 s 1012 13838 1012 13838 4 _0294_
rlabel metal1 s 1196 13430 1196 13430 4 _0295_
rlabel metal1 s 1610 13158 1610 13158 4 _0296_
rlabel metal2 s 1794 15028 1794 15028 4 _0297_
rlabel metal1 s 1610 13498 1610 13498 4 _0298_
rlabel metal2 s 2070 13974 2070 13974 4 _0299_
rlabel metal1 s 1656 14586 1656 14586 4 _0300_
rlabel metal1 s 1626 15606 1626 15606 4 _0301_
rlabel metal1 s 2185 15334 2185 15334 4 _0302_
rlabel metal2 s 21022 19822 21022 19822 4 _0303_
rlabel metal1 s 15824 19890 15824 19890 4 _0304_
rlabel metal1 s 22402 18292 22402 18292 4 _0305_
rlabel metal3 s 16238 20451 16238 20451 4 _0306_
rlabel metal1 s 20838 19448 20838 19448 4 _0307_
rlabel metal2 s 20746 19856 20746 19856 4 _0308_
rlabel metal2 s 19090 19516 19090 19516 4 _0309_
rlabel metal2 s 17618 20468 17618 20468 4 _0310_
rlabel metal2 s 17894 20740 17894 20740 4 _0311_
rlabel metal1 s 15732 20570 15732 20570 4 _0312_
rlabel metal1 s 19182 20570 19182 20570 4 _0313_
rlabel metal1 s 16790 20400 16790 20400 4 _0314_
rlabel metal1 s 16330 21930 16330 21930 4 _0315_
rlabel metal2 s 20286 22338 20286 22338 4 _0316_
rlabel metal1 s 16698 20298 16698 20298 4 _0317_
rlabel metal1 s 20010 21624 20010 21624 4 _0318_
rlabel metal1 s 15456 22406 15456 22406 4 _0319_
rlabel metal1 s 20286 21522 20286 21522 4 _0320_
rlabel metal1 s 20194 22406 20194 22406 4 _0321_
rlabel metal2 s 19044 21998 19044 21998 4 _0322_
rlabel metal3 s 16284 21964 16284 21964 4 _0323_
rlabel metal1 s 19366 21930 19366 21930 4 _0324_
rlabel metal2 s 20838 21760 20838 21760 4 _0325_
rlabel metal1 s 20516 21114 20516 21114 4 _0326_
rlabel metal1 s 16376 22542 16376 22542 4 _0327_
rlabel metal1 s 19458 21386 19458 21386 4 _0328_
rlabel metal1 s 19826 21352 19826 21352 4 _0329_
rlabel metal1 s 8694 17544 8694 17544 4 _0330_
rlabel metal1 s 8326 16762 8326 16762 4 _0331_
rlabel metal2 s 8418 16150 8418 16150 4 _0332_
rlabel metal2 s 7958 17476 7958 17476 4 _0333_
rlabel metal1 s 7958 18258 7958 18258 4 _0334_
rlabel metal2 s 8050 17850 8050 17850 4 _0335_
rlabel metal1 s 7084 17782 7084 17782 4 _0336_
rlabel metal1 s 7452 18258 7452 18258 4 _0337_
rlabel metal1 s 7544 18394 7544 18394 4 _0338_
rlabel metal2 s 8970 17884 8970 17884 4 _0339_
rlabel metal2 s 9062 18496 9062 18496 4 _0340_
rlabel metal2 s 8786 17986 8786 17986 4 _0341_
rlabel metal2 s 7406 17765 7406 17765 4 _0342_
rlabel metal2 s 6486 18564 6486 18564 4 _0343_
rlabel metal1 s 7498 18938 7498 18938 4 _0344_
rlabel metal1 s 9660 20910 9660 20910 4 _0345_
rlabel metal1 s 11316 20366 11316 20366 4 _0346_
rlabel metal2 s 11454 20128 11454 20128 4 _0347_
rlabel metal1 s 13754 20332 13754 20332 4 _0348_
rlabel metal2 s 8510 19278 8510 19278 4 _0349_
rlabel metal2 s 9338 20196 9338 20196 4 _0350_
rlabel metal1 s 10718 21454 10718 21454 4 _0351_
rlabel metal1 s 11178 21012 11178 21012 4 _0352_
rlabel metal2 s 16330 19533 16330 19533 4 _0353_
rlabel metal2 s 2162 21216 2162 21216 4 _0354_
rlabel metal1 s 7774 22066 7774 22066 4 _0355_
rlabel metal1 s 9936 21318 9936 21318 4 _0356_
rlabel metal1 s 10304 21862 10304 21862 4 _0357_
rlabel metal1 s 10120 21658 10120 21658 4 _0358_
rlabel metal1 s 10672 22202 10672 22202 4 _0359_
rlabel metal1 s 10166 20910 10166 20910 4 _0360_
rlabel metal1 s 10212 20366 10212 20366 4 _0361_
rlabel metal1 s 9568 20366 9568 20366 4 _0362_
rlabel metal1 s 10074 20400 10074 20400 4 _0363_
rlabel metal1 s 9798 21930 9798 21930 4 _0364_
rlabel metal1 s 8648 21930 8648 21930 4 _0365_
rlabel metal2 s 18906 21165 18906 21165 4 _0366_
rlabel metal1 s 9200 22202 9200 22202 4 _0367_
rlabel metal1 s 9154 22542 9154 22542 4 _0368_
rlabel metal1 s 2990 21930 2990 21930 4 _0369_
rlabel metal1 s 3358 21522 3358 21522 4 _0370_
rlabel metal1 s 1610 21046 1610 21046 4 _0371_
rlabel metal2 s 1886 21862 1886 21862 4 _0372_
rlabel metal1 s 2484 20774 2484 20774 4 _0373_
rlabel metal2 s 2254 19193 2254 19193 4 _0374_
rlabel metal2 s 2530 21284 2530 21284 4 _0375_
rlabel metal2 s 2530 20162 2530 20162 4 _0376_
rlabel metal1 s 2668 19142 2668 19142 4 _0377_
rlabel metal1 s 2714 18870 2714 18870 4 _0378_
rlabel metal1 s 2484 19686 2484 19686 4 _0379_
rlabel metal2 s 2714 20128 2714 20128 4 _0380_
rlabel metal1 s 3634 19278 3634 19278 4 _0381_
rlabel metal2 s 6670 21012 6670 21012 4 _0382_
rlabel metal2 s 5658 21284 5658 21284 4 _0383_
rlabel metal1 s 8602 20978 8602 20978 4 _0384_
rlabel metal1 s 7682 21930 7682 21930 4 _0385_
rlabel metal1 s 7038 21114 7038 21114 4 _0386_
rlabel metal1 s 7176 21454 7176 21454 4 _0387_
rlabel metal1 s 7268 22202 7268 22202 4 _0388_
rlabel metal1 s 8819 21046 8819 21046 4 _0389_
rlabel metal1 s 7958 20842 7958 20842 4 _0390_
rlabel metal1 s 7774 20910 7774 20910 4 _0391_
rlabel metal1 s 7176 20978 7176 20978 4 _0392_
rlabel metal1 s 7636 22610 7636 22610 4 _0393_
rlabel metal1 s 6624 22542 6624 22542 4 _0394_
rlabel metal2 s 23046 17884 23046 17884 4 _0395_
rlabel metal1 s 22402 10778 22402 10778 4 _0396_
rlabel metal2 s 21482 11866 21482 11866 4 _0397_
rlabel metal1 s 21252 12614 21252 12614 4 _0398_
rlabel metal1 s 21482 18734 21482 18734 4 _0399_
rlabel metal1 s 5106 19142 5106 19142 4 _0400_
rlabel metal1 s 5382 18836 5382 18836 4 _0401_
rlabel metal1 s 4968 8534 4968 8534 4 _0402_
rlabel metal2 s 2714 13634 2714 13634 4 _0403_
rlabel metal2 s 5658 16932 5658 16932 4 _0404_
rlabel metal2 s 2530 15436 2530 15436 4 _0405_
rlabel metal2 s 6578 16218 6578 16218 4 _0406_
rlabel metal2 s 1702 5066 1702 5066 4 _0407_
rlabel metal1 s 3496 7922 3496 7922 4 _0408_
rlabel metal1 s 12236 15606 12236 15606 4 _0409_
rlabel metal1 s 8832 14926 8832 14926 4 _0410_
rlabel metal1 s 8372 13430 8372 13430 4 _0411_
rlabel metal1 s 8464 14450 8464 14450 4 _0412_
rlabel metal1 s 3634 15436 3634 15436 4 _0413_
rlabel metal1 s 4922 12614 4922 12614 4 _0414_
rlabel metal1 s 7038 15130 7038 15130 4 _0415_
rlabel metal1 s 1426 5168 1426 5168 4 _0416_
rlabel metal1 s 782 4658 782 4658 4 _0417_
rlabel metal1 s 6440 14042 6440 14042 4 _0418_
rlabel metal1 s 4002 14892 4002 14892 4 _0419_
rlabel metal1 s 4600 15130 4600 15130 4 _0420_
rlabel metal1 s 6670 16048 6670 16048 4 _0421_
rlabel metal1 s 5842 16218 5842 16218 4 _0422_
rlabel metal1 s 4692 20842 4692 20842 4 _0423_
rlabel metal1 s 4830 20978 4830 20978 4 _0424_
rlabel metal2 s 5290 21284 5290 21284 4 _0425_
rlabel metal2 s 1886 20774 1886 20774 4 _0426_
rlabel metal1 s 2070 20876 2070 20876 4 _0427_
rlabel metal1 s 2530 22202 2530 22202 4 _0428_
rlabel metal1 s 4738 21318 4738 21318 4 _0429_
rlabel metal2 s 5934 20740 5934 20740 4 _0430_
rlabel metal2 s 3450 21862 3450 21862 4 _0431_
rlabel metal1 s 4554 21012 4554 21012 4 _0432_
rlabel metal2 s 6210 21455 6210 21455 4 _0433_
rlabel metal1 s 13524 22542 13524 22542 4 _0434_
rlabel metal1 s 8004 21454 8004 21454 4 _0435_
rlabel metal1 s 5290 19754 5290 19754 4 _0436_
rlabel metal1 s 4968 19890 4968 19890 4 _0437_
rlabel metal1 s 4738 20026 4738 20026 4 _0438_
rlabel metal2 s 22494 9724 22494 9724 4 _0439_
rlabel metal1 s 20654 9146 20654 9146 4 _0440_
rlabel metal2 s 21528 15300 21528 15300 4 _0441_
rlabel metal1 s 21482 18190 21482 18190 4 _0442_
rlabel metal2 s 19366 16762 19366 16762 4 _0443_
rlabel metal2 s 17342 19295 17342 19295 4 _0444_
rlabel metal1 s 14674 21488 14674 21488 4 _0445_
rlabel metal1 s 22908 15946 22908 15946 4 _0446_
rlabel metal1 s 20746 17646 20746 17646 4 _0447_
rlabel metal1 s 21344 17714 21344 17714 4 _0448_
rlabel metal2 s 21942 18122 21942 18122 4 _0449_
rlabel metal1 s 21666 20366 21666 20366 4 _0450_
rlabel metal1 s 23092 16014 23092 16014 4 _0451_
rlabel metal1 s 7360 20910 7360 20910 4 _0452_
rlabel metal1 s 20700 11186 20700 11186 4 _0453_
rlabel metal1 s 20056 6222 20056 6222 4 _0454_
rlabel metal1 s 20700 10574 20700 10574 4 _0455_
rlabel metal1 s 19872 19890 19872 19890 4 _0456_
rlabel metal1 s 20562 11220 20562 11220 4 _0457_
rlabel metal1 s 20838 9520 20838 9520 4 _0458_
rlabel metal1 s 19366 5780 19366 5780 4 _0459_
rlabel metal2 s 21206 5338 21206 5338 4 _0460_
rlabel metal1 s 20930 5032 20930 5032 4 _0461_
rlabel metal1 s 17802 5100 17802 5100 4 _0462_
rlabel metal2 s 20746 1972 20746 1972 4 _0463_
rlabel metal1 s 20700 1870 20700 1870 4 _0464_
rlabel metal2 s 21574 1632 21574 1632 4 _0465_
rlabel metal2 s 4278 17374 4278 17374 4 _0466_
rlabel metal1 s 3450 16592 3450 16592 4 _0467_
rlabel metal1 s 7682 17612 7682 17612 4 _0468_
rlabel metal1 s 5888 17102 5888 17102 4 _0469_
rlabel metal1 s 13754 7242 13754 7242 4 _0470_
rlabel metal2 s 8234 16898 8234 16898 4 _0471_
rlabel metal3 s 8579 13668 8579 13668 4 _0472_
rlabel metal1 s 12098 2924 12098 2924 4 _0473_
rlabel metal1 s 20930 2482 20930 2482 4 _0474_
rlabel metal4 s 19021 19380 19021 19380 4 _0475_
rlabel metal1 s 21390 2992 21390 2992 4 _0476_
rlabel metal1 s 20286 6256 20286 6256 4 _0477_
rlabel metal1 s 20010 6426 20010 6426 4 _0478_
rlabel metal1 s 16790 5746 16790 5746 4 _0479_
rlabel metal1 s 14812 20570 14812 20570 4 _0480_
rlabel metal2 s 15318 20570 15318 20570 4 _0481_
rlabel metal2 s 19550 14586 19550 14586 4 _0482_
rlabel metal2 s 19366 15045 19366 15045 4 _0483_
rlabel metal2 s 21390 14654 21390 14654 4 _0484_
rlabel metal1 s 19504 13838 19504 13838 4 _0485_
rlabel metal1 s 19550 9962 19550 9962 4 _0486_
rlabel metal2 s 9614 6273 9614 6273 4 _0487_
rlabel metal1 s 22586 10472 22586 10472 4 _0488_
rlabel metal1 s 22402 9520 22402 9520 4 _0489_
rlabel metal2 s 19826 7106 19826 7106 4 _0490_
rlabel metal1 s 20378 6800 20378 6800 4 _0491_
rlabel metal1 s 19366 7344 19366 7344 4 _0492_
rlabel metal1 s 13156 16422 13156 16422 4 _0493_
rlabel metal1 s 11224 14586 11224 14586 4 _0494_
rlabel metal1 s 15916 17102 15916 17102 4 _0495_
rlabel metal1 s 13064 16626 13064 16626 4 _0496_
rlabel metal2 s 12926 17102 12926 17102 4 _0497_
rlabel metal1 s 13386 15504 13386 15504 4 _0498_
rlabel metal2 s 13846 15266 13846 15266 4 _0499_
rlabel metal2 s 12834 14620 12834 14620 4 _0500_
rlabel metal1 s 19458 7412 19458 7412 4 _0501_
rlabel metal1 s 20516 8398 20516 8398 4 _0502_
rlabel metal1 s 20056 7378 20056 7378 4 _0503_
rlabel metal2 s 19366 10336 19366 10336 4 _0504_
rlabel metal2 s 20194 6970 20194 6970 4 _0505_
rlabel metal1 s 20792 6426 20792 6426 4 _0506_
rlabel metal1 s 20102 13362 20102 13362 4 _0507_
rlabel metal1 s 19642 13872 19642 13872 4 _0508_
rlabel metal2 s 20470 14620 20470 14620 4 _0509_
rlabel metal2 s 20378 14620 20378 14620 4 _0510_
rlabel metal2 s 19872 9010 19872 9010 4 _0511_
rlabel metal1 s 21528 11186 21528 11186 4 _0512_
rlabel metal1 s 20194 10574 20194 10574 4 _0513_
rlabel metal1 s 18492 13294 18492 13294 4 _0514_
rlabel metal1 s 9844 9418 9844 9418 4 _0515_
rlabel metal2 s 17894 9248 17894 9248 4 _0516_
rlabel metal2 s 19964 8908 19964 8908 4 _0517_
rlabel metal2 s 14306 9741 14306 9741 4 _0518_
rlabel metal2 s 9430 9996 9430 9996 4 _0519_
rlabel metal2 s 8418 7361 8418 7361 4 _0520_
rlabel metal1 s 21298 6188 21298 6188 4 _0521_
rlabel metal2 s 19918 9707 19918 9707 4 _0522_
rlabel metal2 s 12098 14501 12098 14501 4 _0523_
rlabel metal1 s 13294 10064 13294 10064 4 _0524_
rlabel metal1 s 13984 6222 13984 6222 4 _0525_
rlabel metal1 s 19182 6324 19182 6324 4 _0526_
rlabel metal2 s 14214 6273 14214 6273 4 _0527_
rlabel metal2 s 19090 5984 19090 5984 4 _0528_
rlabel metal1 s 21206 6256 21206 6256 4 _0529_
rlabel metal2 s 21298 4522 21298 4522 4 _0530_
rlabel metal1 s 21298 4522 21298 4522 4 _0531_
rlabel metal1 s 22034 4658 22034 4658 4 _0532_
rlabel metal1 s 21390 2550 21390 2550 4 _0533_
rlabel metal1 s 22310 2448 22310 2448 4 _0534_
rlabel metal2 s 8694 13600 8694 13600 4 _0535_
rlabel metal1 s 9798 14484 9798 14484 4 _0536_
rlabel metal1 s 11638 13804 11638 13804 4 _0537_
rlabel metal2 s 11822 13940 11822 13940 4 _0538_
rlabel metal1 s 9614 13396 9614 13396 4 _0539_
rlabel metal2 s 1794 22746 1794 22746 4 _0540_
rlabel metal1 s 1748 22202 1748 22202 4 _0541_
rlabel metal1 s 1794 22610 1794 22610 4 _0542_
rlabel metal1 s 5520 23086 5520 23086 4 _0543_
rlabel metal2 s 5750 22950 5750 22950 4 _0544_
rlabel metal1 s 5750 22134 5750 22134 4 _0545_
rlabel metal1 s 9890 22032 9890 22032 4 _0546_
rlabel metal1 s 12742 22508 12742 22508 4 _0547_
rlabel metal1 s 10534 19278 10534 19278 4 _0548_
rlabel metal1 s 14490 20910 14490 20910 4 _0549_
rlabel metal1 s 14398 20570 14398 20570 4 _0550_
rlabel metal2 s 14214 21862 14214 21862 4 _0551_
rlabel metal1 s 14306 22134 14306 22134 4 _0552_
rlabel metal1 s 13984 22474 13984 22474 4 _0553_
rlabel metal1 s 12558 21454 12558 21454 4 _0554_
rlabel metal1 s 12627 22610 12627 22610 4 _0555_
rlabel metal1 s 4830 21930 4830 21930 4 _0556_
rlabel metal1 s 4094 22066 4094 22066 4 _0557_
rlabel metal1 s 4554 22406 4554 22406 4 _0558_
rlabel metal1 s 4370 21998 4370 21998 4 _0559_
rlabel metal1 s 4462 22066 4462 22066 4 _0560_
rlabel metal1 s 2714 22644 2714 22644 4 _0561_
rlabel metal1 s 1840 22406 1840 22406 4 _0562_
rlabel metal2 s 2070 20060 2070 20060 4 _0563_
rlabel metal1 s 1518 19890 1518 19890 4 _0564_
rlabel metal2 s 1886 19482 1886 19482 4 _0565_
rlabel metal1 s 736 19346 736 19346 4 _0566_
rlabel metal1 s 1978 8976 1978 8976 4 _0567_
rlabel metal2 s 9614 9486 9614 9486 4 _0568_
rlabel metal1 s 10174 13838 10174 13838 4 _0569_
rlabel metal3 s 3174 7939 3174 7939 4 _0570_
rlabel metal1 s 2484 1938 2484 1938 4 _0571_
rlabel metal1 s 9752 11322 9752 11322 4 _0572_
rlabel metal1 s 13892 13702 13892 13702 4 _0573_
rlabel metal1 s 9430 13328 9430 13328 4 _0574_
rlabel metal1 s 11178 12784 11178 12784 4 _0575_
rlabel metal1 s 4830 22542 4830 22542 4 _0576_
rlabel metal1 s 5106 4046 5106 4046 4 _0577_
rlabel metal1 s 2162 4624 2162 4624 4 _0578_
rlabel metal1 s 7314 6256 7314 6256 4 _0579_
rlabel metal3 s 6647 20740 6647 20740 4 _0580_
rlabel metal2 s 6210 10370 6210 10370 4 _0581_
rlabel metal1 s 6992 12818 6992 12818 4 _0582_
rlabel metal2 s 11370 17034 11370 17034 4 _0583_
rlabel metal1 s 9384 12954 9384 12954 4 _0584_
rlabel metal1 s 9798 13498 9798 13498 4 _0585_
rlabel metal1 s 12282 21522 12282 21522 4 _0586_
rlabel metal2 s 12834 13345 12834 13345 4 _0587_
rlabel metal1 s 8786 12716 8786 12716 4 _0588_
rlabel metal1 s 11914 11764 11914 11764 4 _0589_
rlabel metal1 s 11500 13362 11500 13362 4 _0590_
rlabel metal1 s 14398 22406 14398 22406 4 _0591_
rlabel metal2 s 15042 18700 15042 18700 4 _0592_
rlabel metal2 s 15502 14620 15502 14620 4 _0593_
rlabel metal1 s 15732 13294 15732 13294 4 _0594_
rlabel metal2 s 11270 13668 11270 13668 4 _0595_
rlabel metal1 s 17066 15980 17066 15980 4 _0596_
rlabel metal2 s 17894 15708 17894 15708 4 _0597_
rlabel metal1 s 21574 15980 21574 15980 4 _0598_
rlabel metal1 s 20194 15538 20194 15538 4 _0599_
rlabel metal2 s 10994 13124 10994 13124 4 _0600_
rlabel metal1 s 9246 15980 9246 15980 4 _0601_
rlabel metal1 s 9154 18224 9154 18224 4 _0602_
rlabel metal1 s 10994 13464 10994 13464 4 _0603_
rlabel metal1 s 16054 12410 16054 12410 4 _0604_
rlabel metal2 s 1978 19380 1978 19380 4 _0605_
rlabel metal1 s 4416 18734 4416 18734 4 _0606_
rlabel metal2 s 8786 15249 8786 15249 4 _0607_
rlabel metal1 s 6532 19890 6532 19890 4 _0608_
rlabel metal2 s 2438 15181 2438 15181 4 _0609_
rlabel metal1 s 9200 15130 9200 15130 4 _0610_
rlabel metal2 s 9430 14892 9430 14892 4 _0611_
rlabel metal2 s 10258 2125 10258 2125 4 _0612_
rlabel metal3 s 20746 2448 20746 2448 4 _0613_
rlabel metal1 s 17802 2856 17802 2856 4 _0614_
rlabel metal1 s 21758 2550 21758 2550 4 _0615_
rlabel metal2 s 21390 2074 21390 2074 4 _0616_
rlabel metal1 s 20654 5338 20654 5338 4 _0617_
rlabel metal1 s 19067 3366 19067 3366 4 _0618_
rlabel metal2 s 20378 4794 20378 4794 4 _0619_
rlabel metal1 s 18906 3570 18906 3570 4 _0620_
rlabel metal2 s 21758 2618 21758 2618 4 _0621_
rlabel metal1 s 18032 12410 18032 12410 4 _0622_
rlabel metal1 s 22494 10132 22494 10132 4 _0623_
rlabel metal1 s 17802 9078 17802 9078 4 _0624_
rlabel metal1 s 18354 8398 18354 8398 4 _0625_
rlabel metal2 s 21942 7786 21942 7786 4 _0626_
rlabel metal2 s 21114 15980 21114 15980 4 _0627_
rlabel metal1 s 21344 16762 21344 16762 4 _0628_
rlabel metal1 s 19228 9010 19228 9010 4 _0629_
rlabel metal1 s 8234 13770 8234 13770 4 _0630_
rlabel metal2 s 8786 14178 8786 14178 4 _0631_
rlabel metal4 s 12972 13192 12972 13192 4 _0632_
rlabel metal1 s 19596 7922 19596 7922 4 _0633_
rlabel metal1 s 18400 6290 18400 6290 4 _0634_
rlabel metal3 s 20631 18020 20631 18020 4 _0635_
rlabel metal1 s 18492 5610 18492 5610 4 _0636_
rlabel metal1 s 20378 16014 20378 16014 4 _0637_
rlabel metal2 s 20102 16218 20102 16218 4 _0638_
rlabel metal1 s 20424 15334 20424 15334 4 _0639_
rlabel metal2 s 20286 14620 20286 14620 4 _0640_
rlabel metal1 s 20056 12274 20056 12274 4 _0641_
rlabel metal1 s 19366 12308 19366 12308 4 _0642_
rlabel metal1 s 18814 11084 18814 11084 4 _0643_
rlabel metal1 s 14214 7242 14214 7242 4 _0644_
rlabel metal2 s 20102 12308 20102 12308 4 _0645_
rlabel metal2 s 18584 9146 18584 9146 4 _0646_
rlabel metal1 s 17710 6154 17710 6154 4 _0647_
rlabel metal1 s 17618 6086 17618 6086 4 _0648_
rlabel metal2 s 18538 5814 18538 5814 4 _0649_
rlabel metal1 s 19642 11016 19642 11016 4 _0650_
rlabel metal2 s 12006 10557 12006 10557 4 _0651_
rlabel metal1 s 8004 14450 8004 14450 4 _0652_
rlabel metal1 s 15778 9622 15778 9622 4 _0653_
rlabel metal1 s 19550 11118 19550 11118 4 _0654_
rlabel metal1 s 7820 8942 7820 8942 4 _0655_
rlabel metal3 s 16698 9469 16698 9469 4 _0656_
rlabel metal1 s 18216 10098 18216 10098 4 _0657_
rlabel metal1 s 6624 7922 6624 7922 4 _0658_
rlabel metal1 s 21942 15572 21942 15572 4 _0659_
rlabel metal1 s 22126 14416 22126 14416 4 _0660_
rlabel metal2 s 22494 14042 22494 14042 4 _0661_
rlabel metal2 s 21390 16626 21390 16626 4 _0662_
rlabel metal2 s 22034 14943 22034 14943 4 _0663_
rlabel metal2 s 21666 14042 21666 14042 4 _0664_
rlabel metal1 s 22218 13906 22218 13906 4 _0665_
rlabel metal1 s 19642 13226 19642 13226 4 _0666_
rlabel metal1 s 18400 10438 18400 10438 4 _0667_
rlabel metal1 s 18492 5746 18492 5746 4 _0668_
rlabel metal1 s 18814 4658 18814 4658 4 _0669_
rlabel metal1 s 19734 5338 19734 5338 4 _0670_
rlabel metal1 s 19182 4590 19182 4590 4 _0671_
rlabel metal1 s 18722 4590 18722 4590 4 _0672_
rlabel metal2 s 18814 3468 18814 3468 4 _0673_
rlabel metal1 s 13754 2992 13754 2992 4 _0674_
rlabel metal1 s 17940 2550 17940 2550 4 _0675_
rlabel metal2 s 18630 1836 18630 1836 4 _0676_
rlabel metal2 s 18998 782 18998 782 4 _0677_
rlabel metal2 s 20838 714 20838 714 4 _0678_
rlabel metal1 s 17342 2958 17342 2958 4 _0679_
rlabel metal1 s 16330 2550 16330 2550 4 _0680_
rlabel metal2 s 12926 2176 12926 2176 4 _0681_
rlabel metal1 s 15732 2550 15732 2550 4 _0682_
rlabel metal1 s 16192 2278 16192 2278 4 _0683_
rlabel metal1 s 19274 12240 19274 12240 4 _0684_
rlabel metal1 s 14306 16626 14306 16626 4 _0685_
rlabel metal1 s 17158 13362 17158 13362 4 _0686_
rlabel metal2 s 17526 14892 17526 14892 4 _0687_
rlabel metal1 s 17388 13294 17388 13294 4 _0688_
rlabel metal2 s 18906 12954 18906 12954 4 _0689_
rlabel metal2 s 18814 12716 18814 12716 4 _0690_
rlabel metal2 s 19274 11917 19274 11917 4 _0691_
rlabel metal1 s 18446 11594 18446 11594 4 _0692_
rlabel metal2 s 19550 12223 19550 12223 4 _0693_
rlabel metal1 s 18538 11662 18538 11662 4 _0694_
rlabel metal2 s 15686 15691 15686 15691 4 _0695_
rlabel metal1 s 18860 15402 18860 15402 4 _0696_
rlabel metal2 s 17434 15538 17434 15538 4 _0697_
rlabel metal1 s 18814 15504 18814 15504 4 _0698_
rlabel metal1 s 18814 14994 18814 14994 4 _0699_
rlabel metal1 s 19320 13906 19320 13906 4 _0700_
rlabel metal1 s 18584 12410 18584 12410 4 _0701_
rlabel metal1 s 18860 17102 18860 17102 4 _0702_
rlabel metal1 s 18722 17068 18722 17068 4 _0703_
rlabel metal1 s 18722 16660 18722 16660 4 _0704_
rlabel metal1 s 19366 16694 19366 16694 4 _0705_
rlabel metal1 s 17986 12240 17986 12240 4 _0706_
rlabel metal1 s 18446 11730 18446 11730 4 _0707_
rlabel metal2 s 18814 11968 18814 11968 4 _0708_
rlabel metal2 s 17434 5185 17434 5185 4 _0709_
rlabel metal1 s 16882 11696 16882 11696 4 _0710_
rlabel metal1 s 18584 11798 18584 11798 4 _0711_
rlabel metal2 s 13386 10336 13386 10336 4 _0712_
rlabel metal2 s 15318 7276 15318 7276 4 _0713_
rlabel metal2 s 18078 8670 18078 8670 4 _0714_
rlabel metal1 s 18078 7922 18078 7922 4 _0715_
rlabel metal1 s 17158 18122 17158 18122 4 _0716_
rlabel metal2 s 4922 15538 4922 15538 4 _0717_
rlabel metal2 s 15916 9996 15916 9996 4 _0718_
rlabel metal1 s 18952 7922 18952 7922 4 _0719_
rlabel metal1 s 19274 6256 19274 6256 4 _0720_
rlabel metal1 s 17986 5780 17986 5780 4 _0721_
rlabel metal2 s 17342 4318 17342 4318 4 _0722_
rlabel metal2 s 17434 3230 17434 3230 4 _0723_
rlabel metal1 s 16744 782 16744 782 4 _0724_
rlabel metal1 s 16652 986 16652 986 4 _0725_
rlabel metal1 s 21482 3434 21482 3434 4 _0726_
rlabel metal1 s 20884 3570 20884 3570 4 _0727_
rlabel metal1 s 19918 1972 19918 1972 4 _0728_
rlabel metal2 s 15226 1479 15226 1479 4 _0729_
rlabel metal1 s 17434 4522 17434 4522 4 _0730_
rlabel metal1 s 9062 9486 9062 9486 4 _0731_
rlabel metal1 s 15410 12852 15410 12852 4 _0732_
rlabel metal1 s 12742 15606 12742 15606 4 _0733_
rlabel metal2 s 13018 14416 13018 14416 4 _0734_
rlabel metal1 s 12880 14926 12880 14926 4 _0735_
rlabel metal1 s 12972 14042 12972 14042 4 _0736_
rlabel metal2 s 14214 12954 14214 12954 4 _0737_
rlabel metal1 s 15134 12682 15134 12682 4 _0738_
rlabel metal1 s 15134 12784 15134 12784 4 _0739_
rlabel metal1 s 15180 12886 15180 12886 4 _0740_
rlabel metal1 s 14904 10642 14904 10642 4 _0741_
rlabel metal1 s 15732 17714 15732 17714 4 _0742_
rlabel metal1 s 14720 15402 14720 15402 4 _0743_
rlabel metal2 s 13938 14348 13938 14348 4 _0744_
rlabel metal1 s 15088 13838 15088 13838 4 _0745_
rlabel metal2 s 8418 13464 8418 13464 4 _0746_
rlabel metal1 s 15226 13872 15226 13872 4 _0747_
rlabel metal1 s 14996 13702 14996 13702 4 _0748_
rlabel metal1 s 14858 13838 14858 13838 4 _0749_
rlabel metal1 s 14904 13158 14904 13158 4 _0750_
rlabel metal1 s 15594 15504 15594 15504 4 _0751_
rlabel metal2 s 13846 15810 13846 15810 4 _0752_
rlabel metal1 s 13570 16048 13570 16048 4 _0753_
rlabel metal1 s 14858 15980 14858 15980 4 _0754_
rlabel metal1 s 17020 16082 17020 16082 4 _0755_
rlabel metal1 s 14950 15878 14950 15878 4 _0756_
rlabel metal1 s 15318 11322 15318 11322 4 _0757_
rlabel metal1 s 17342 11118 17342 11118 4 _0758_
rlabel metal1 s 15364 11186 15364 11186 4 _0759_
rlabel metal1 s 15548 11186 15548 11186 4 _0760_
rlabel metal2 s 16698 12750 16698 12750 4 _0761_
rlabel metal1 s 15824 11254 15824 11254 4 _0762_
rlabel metal2 s 15318 10812 15318 10812 4 _0763_
rlabel metal1 s 15042 10778 15042 10778 4 _0764_
rlabel metal1 s 8970 5814 8970 5814 4 _0765_
rlabel metal1 s 13340 8398 13340 8398 4 _0766_
rlabel metal1 s 14214 18156 14214 18156 4 _0767_
rlabel metal3 s 14398 18037 14398 18037 4 _0768_
rlabel metal1 s 15088 8806 15088 8806 4 _0769_
rlabel metal1 s 3680 5134 3680 5134 4 _0770_
rlabel metal1 s 3542 1326 3542 1326 4 _0771_
rlabel metal1 s 14030 10574 14030 10574 4 _0772_
rlabel metal1 s 14582 7850 14582 7850 4 _0773_
rlabel metal1 s 15318 6256 15318 6256 4 _0774_
rlabel metal1 s 15410 6188 15410 6188 4 _0775_
rlabel metal1 s 14996 6426 14996 6426 4 _0776_
rlabel metal2 s 15318 5406 15318 5406 4 _0777_
rlabel metal2 s 15226 4828 15226 4828 4 _0778_
rlabel metal1 s 15548 4046 15548 4046 4 _0779_
rlabel metal1 s 15088 3910 15088 3910 4 _0780_
rlabel metal1 s 14904 2550 14904 2550 4 _0781_
rlabel metal2 s 15410 2414 15410 2414 4 _0782_
rlabel metal1 s 14808 1530 14808 1530 4 _0783_
rlabel metal1 s 14536 1462 14536 1462 4 _0784_
rlabel metal1 s 14490 6222 14490 6222 4 _0785_
rlabel metal2 s 13892 4046 13892 4046 4 _0786_
rlabel metal1 s 11960 5746 11960 5746 4 _0787_
rlabel metal1 s 13340 12954 13340 12954 4 _0788_
rlabel metal1 s 6486 10778 6486 10778 4 _0789_
rlabel metal1 s 6946 14246 6946 14246 4 _0790_
rlabel metal1 s 7314 12240 7314 12240 4 _0791_
rlabel metal2 s 7130 11594 7130 11594 4 _0792_
rlabel metal2 s 8694 10812 8694 10812 4 _0793_
rlabel metal1 s 9522 13838 9522 13838 4 _0794_
rlabel metal1 s 10074 10676 10074 10676 4 _0795_
rlabel metal1 s 10120 10098 10120 10098 4 _0796_
rlabel metal2 s 9982 10268 9982 10268 4 _0797_
rlabel metal1 s 13018 13736 13018 13736 4 _0798_
rlabel metal2 s 13846 14042 13846 14042 4 _0799_
rlabel metal1 s 12926 13362 12926 13362 4 _0800_
rlabel metal2 s 8602 11628 8602 11628 4 _0801_
rlabel metal1 s 8648 12750 8648 12750 4 _0802_
rlabel metal2 s 8878 12444 8878 12444 4 _0803_
rlabel metal1 s 8970 11764 8970 11764 4 _0804_
rlabel metal1 s 9568 11662 9568 11662 4 _0805_
rlabel metal1 s 10304 15538 10304 15538 4 _0806_
rlabel metal1 s 10304 15402 10304 15402 4 _0807_
rlabel metal1 s 9614 16048 9614 16048 4 _0808_
rlabel metal1 s 9522 16116 9522 16116 4 _0809_
rlabel metal2 s 9936 15878 9936 15878 4 _0810_
rlabel metal1 s 10212 11526 10212 11526 4 _0811_
rlabel metal2 s 7682 11356 7682 11356 4 _0812_
rlabel metal1 s 10488 11662 10488 11662 4 _0813_
rlabel metal1 s 12788 11050 12788 11050 4 _0814_
rlabel metal1 s 14306 7310 14306 7310 4 _0815_
rlabel metal1 s 12558 10982 12558 10982 4 _0816_
rlabel metal1 s 9890 10132 9890 10132 4 _0817_
rlabel metal1 s 11178 9962 11178 9962 4 _0818_
rlabel metal2 s 13294 14620 13294 14620 4 _0819_
rlabel metal1 s 12834 18802 12834 18802 4 _0820_
rlabel metal2 s 10764 9486 10764 9486 4 _0821_
rlabel metal3 s 1426 9469 1426 9469 4 _0822_
rlabel metal1 s 6440 12614 6440 12614 4 _0823_
rlabel metal1 s 12558 9554 12558 9554 4 _0824_
rlabel metal1 s 13248 5678 13248 5678 4 _0825_
rlabel metal1 s 12374 5610 12374 5610 4 _0826_
rlabel metal1 s 20332 5678 20332 5678 4 _0827_
rlabel metal1 s 12788 5338 12788 5338 4 _0828_
rlabel metal2 s 11638 4284 11638 4284 4 _0829_
rlabel metal2 s 20378 3485 20378 3485 4 _0830_
rlabel metal2 s 11178 2550 11178 2550 4 _0831_
rlabel metal2 s 11546 2720 11546 2720 4 _0832_
rlabel metal1 s 11408 1870 11408 1870 4 _0833_
rlabel metal2 s 11362 1190 11362 1190 4 _0834_
rlabel metal1 s 20148 782 20148 782 4 _0835_
rlabel metal1 s 15548 6630 15548 6630 4 _0836_
rlabel metal2 s 13018 7888 13018 7888 4 _0837_
rlabel metal1 s 15916 7718 15916 7718 4 _0838_
rlabel metal1 s 5934 10166 5934 10166 4 _0839_
rlabel metal2 s 11822 13294 11822 13294 4 _0840_
rlabel metal1 s 5980 14790 5980 14790 4 _0841_
rlabel metal2 s 11546 7820 11546 7820 4 _0842_
rlabel metal1 s 11730 5134 11730 5134 4 _0843_
rlabel metal1 s 15180 4998 15180 4998 4 _0844_
rlabel metal2 s 9246 4964 9246 4964 4 _0845_
rlabel metal1 s 8970 10098 8970 10098 4 _0846_
rlabel metal2 s 8234 10268 8234 10268 4 _0847_
rlabel metal1 s 5520 4046 5520 4046 4 _0848_
rlabel metal1 s 3312 6222 3312 6222 4 _0849_
rlabel metal1 s 5152 4794 5152 4794 4 _0850_
rlabel metal2 s 5382 4794 5382 4794 4 _0851_
rlabel metal1 s 6072 5066 6072 5066 4 _0852_
rlabel metal1 s 6716 5678 6716 5678 4 _0853_
rlabel metal1 s 7360 10030 7360 10030 4 _0854_
rlabel metal2 s 8602 9690 8602 9690 4 _0855_
rlabel metal1 s 8050 4216 8050 4216 4 _0856_
rlabel metal1 s 8648 9690 8648 9690 4 _0857_
rlabel metal2 s 3634 13600 3634 13600 4 _0858_
rlabel metal1 s 4968 10234 4968 10234 4 _0859_
rlabel metal1 s 5428 10778 5428 10778 4 _0860_
rlabel metal1 s 4738 5134 4738 5134 4 _0861_
rlabel metal1 s 5658 11220 5658 11220 4 _0862_
rlabel metal1 s 6026 11152 6026 11152 4 _0863_
rlabel metal2 s 6118 11390 6118 11390 4 _0864_
rlabel metal1 s 6808 11186 6808 11186 4 _0865_
rlabel metal1 s 4646 12308 4646 12308 4 _0866_
rlabel metal1 s 5152 12274 5152 12274 4 _0867_
rlabel metal1 s 6026 12308 6026 12308 4 _0868_
rlabel metal2 s 5980 12206 5980 12206 4 _0869_
rlabel metal1 s 6578 11254 6578 11254 4 _0870_
rlabel metal1 s 7360 10778 7360 10778 4 _0871_
rlabel metal1 s 7866 11220 7866 11220 4 _0872_
rlabel metal1 s 7682 12886 7682 12886 4 _0873_
rlabel metal1 s 7527 9486 7527 9486 4 _0874_
rlabel metal1 s 8694 10132 8694 10132 4 _0875_
rlabel metal2 s 11362 5185 11362 5185 4 _0876_
rlabel metal1 s 11684 4658 11684 4658 4 _0877_
rlabel metal2 s 12374 4012 12374 4012 4 _0878_
rlabel metal1 s 15686 3944 15686 3944 4 _0879_
rlabel metal1 s 12374 3366 12374 3366 4 _0880_
rlabel metal1 s 13064 3570 13064 3570 4 _0881_
rlabel metal1 s 12880 3706 12880 3706 4 _0882_
rlabel metal1 s 12006 3400 12006 3400 4 _0883_
rlabel metal1 s 12793 1462 12793 1462 4 _0884_
rlabel metal1 s 12383 1394 12383 1394 4 _0885_
rlabel metal3 s 19734 1411 19734 1411 4 _0886_
rlabel metal2 s 17802 1921 17802 1921 4 _0887_
rlabel metal1 s 9430 1326 9430 1326 4 _0888_
rlabel metal1 s 10948 1734 10948 1734 4 _0889_
rlabel metal1 s 9154 3638 9154 3638 4 _0890_
rlabel metal1 s 15134 4624 15134 4624 4 _0891_
rlabel metal2 s 14950 4352 14950 4352 4 _0892_
rlabel metal1 s 6946 3910 6946 3910 4 _0893_
rlabel metal2 s 3450 2176 3450 2176 4 _0894_
rlabel metal2 s 4278 5066 4278 5066 4 _0895_
rlabel metal1 s 4232 5338 4232 5338 4 _0896_
rlabel metal2 s 4186 5270 4186 5270 4 _0897_
rlabel metal1 s 5842 4046 5842 4046 4 _0898_
rlabel metal1 s 5842 4114 5842 4114 4 _0899_
rlabel metal1 s 6624 4046 6624 4046 4 _0900_
rlabel metal1 s 7820 3910 7820 3910 4 _0901_
rlabel metal2 s 7038 4641 7038 4641 4 _0902_
rlabel metal1 s 7820 4250 7820 4250 4 _0903_
rlabel metal3 s 6762 1411 6762 1411 4 _0904_
rlabel metal1 s 4738 11322 4738 11322 4 _0905_
rlabel metal1 s 3910 1972 3910 1972 4 _0906_
rlabel metal2 s 5750 1632 5750 1632 4 _0907_
rlabel metal2 s 5934 1258 5934 1258 4 _0908_
rlabel metal2 s 6210 986 6210 986 4 _0909_
rlabel metal2 s 6854 1156 6854 1156 4 _0910_
rlabel metal1 s 7222 1870 7222 1870 4 _0911_
rlabel metal1 s 4416 3570 4416 3570 4 _0912_
rlabel metal1 s 4968 3570 4968 3570 4 _0913_
rlabel metal2 s 4646 3196 4646 3196 4 _0914_
rlabel metal3 s 5014 3043 5014 3043 4 _0915_
rlabel metal1 s 6992 2482 6992 2482 4 _0916_
rlabel metal1 s 7360 2074 7360 2074 4 _0917_
rlabel metal1 s 7544 2618 7544 2618 4 _0918_
rlabel metal2 s 7820 7378 7820 7378 4 _0919_
rlabel metal1 s 6791 6834 6791 6834 4 _0920_
rlabel metal1 s 7130 3162 7130 3162 4 _0921_
rlabel metal2 s 8418 4386 8418 4386 4 _0922_
rlabel metal1 s 9522 5678 9522 5678 4 _0923_
rlabel metal1 s 13938 5134 13938 5134 4 _0924_
rlabel metal1 s 12972 4250 12972 4250 4 _0925_
rlabel metal1 s 6716 5610 6716 5610 4 _0926_
rlabel metal1 s 11040 18122 11040 18122 4 _0927_
rlabel metal1 s 11408 6766 11408 6766 4 _0928_
rlabel metal1 s 8924 6630 8924 6630 4 _0929_
rlabel metal3 s 5773 13804 5773 13804 4 _0930_
rlabel metal2 s 9614 6630 9614 6630 4 _0931_
rlabel metal2 s 10258 5610 10258 5610 4 _0932_
rlabel metal1 s 8418 4080 8418 4080 4 _0933_
rlabel metal1 s 9430 3060 9430 3060 4 _0934_
rlabel metal1 s 8510 3536 8510 3536 4 _0935_
rlabel metal2 s 9338 3230 9338 3230 4 _0936_
rlabel metal3 s 14122 3587 14122 3587 4 _0937_
rlabel metal1 s 8648 2550 8648 2550 4 _0938_
rlabel metal1 s 13938 2958 13938 2958 4 _0939_
rlabel metal2 s 13524 2482 13524 2482 4 _0940_
rlabel metal1 s 7728 1394 7728 1394 4 _0941_
rlabel metal1 s 8234 1938 8234 1938 4 _0942_
rlabel metal1 s 8234 1734 8234 1734 4 _0943_
rlabel metal1 s 6670 4658 6670 4658 4 _0944_
rlabel metal1 s 4600 4794 4600 4794 4 _0945_
rlabel metal1 s 10258 7888 10258 7888 4 _0946_
rlabel metal1 s 4784 7854 4784 7854 4 _0947_
rlabel metal2 s 5106 6732 5106 6732 4 _0948_
rlabel metal1 s 5750 5134 5750 5134 4 _0949_
rlabel metal1 s 7130 5168 7130 5168 4 _0950_
rlabel metal1 s 6900 4794 6900 4794 4 _0951_
rlabel metal2 s 17618 10625 17618 10625 4 _0952_
rlabel metal2 s 4462 6902 4462 6902 4 _0953_
rlabel metal2 s 6026 1190 6026 1190 4 _0954_
rlabel metal1 s 2162 1870 2162 1870 4 _0955_
rlabel metal2 s 2714 1598 2714 1598 4 _0956_
rlabel metal1 s 4140 1394 4140 1394 4 _0957_
rlabel metal1 s 3818 1326 3818 1326 4 _0958_
rlabel metal1 s 4370 1292 4370 1292 4 _0959_
rlabel metal1 s 5014 1292 5014 1292 4 _0960_
rlabel metal2 s 6394 3400 6394 3400 4 _0961_
rlabel metal1 s 7130 7820 7130 7820 4 _0962_
rlabel metal1 s 6486 5678 6486 5678 4 _0963_
rlabel metal2 s 6946 5338 6946 5338 4 _0964_
rlabel metal3 s 16330 6205 16330 6205 4 _0965_
rlabel metal1 s 8004 5202 8004 5202 4 _0966_
rlabel metal1 s 13248 5882 13248 5882 4 _0967_
rlabel metal2 s 9246 7616 9246 7616 4 _0968_
rlabel metal1 s 5980 15674 5980 15674 4 _0969_
rlabel metal1 s 6854 15470 6854 15470 4 _0970_
rlabel metal1 s 6624 15334 6624 15334 4 _0971_
rlabel metal1 s 9568 7378 9568 7378 4 _0972_
rlabel metal2 s 9154 6188 9154 6188 4 _0973_
rlabel metal1 s 8556 5338 8556 5338 4 _0974_
rlabel metal1 s 9062 3638 9062 3638 4 _0975_
rlabel metal2 s 8970 3774 8970 3774 4 _0976_
rlabel metal1 s 9292 3570 9292 3570 4 _0977_
rlabel metal2 s 8786 2924 8786 2924 4 _0978_
rlabel metal1 s 10028 2550 10028 2550 4 _0979_
rlabel metal1 s 9890 2482 9890 2482 4 _0980_
rlabel metal2 s 9154 1666 9154 1666 4 _0981_
rlabel metal1 s 9200 1326 9200 1326 4 _0982_
rlabel metal2 s 8510 1190 8510 1190 4 _0983_
rlabel metal1 s 17066 1428 17066 1428 4 _0984_
rlabel metal1 s 20240 7378 20240 7378 4 _0985_
rlabel metal1 s 21666 9452 21666 9452 4 _0986_
rlabel metal1 s 21022 8364 21022 8364 4 _0987_
rlabel metal1 s 20792 8262 20792 8262 4 _0988_
rlabel metal1 s 21068 6766 21068 6766 4 _0989_
rlabel metal2 s 21482 6188 21482 6188 4 _0990_
rlabel metal2 s 19366 14433 19366 14433 4 _0991_
rlabel metal1 s 14674 10642 14674 10642 4 _0992_
rlabel metal2 s 14490 9741 14490 9741 4 _0993_
rlabel metal3 s 16146 10115 16146 10115 4 _0994_
rlabel metal1 s 18078 10132 18078 10132 4 _0995_
rlabel metal1 s 18722 10030 18722 10030 4 _0996_
rlabel metal2 s 21574 6052 21574 6052 4 _0997_
rlabel metal1 s 21942 5338 21942 5338 4 _0998_
rlabel metal1 s 21390 4692 21390 4692 4 _0999_
rlabel metal1 s 21758 4454 21758 4454 4 _1000_
rlabel metal2 s 21942 1802 21942 1802 4 _1001_
rlabel metal2 s 15778 1564 15778 1564 4 _1002_
rlabel metal2 s 18906 17595 18906 17595 4 _1003_
rlabel metal1 s 17388 7378 17388 7378 4 _1004_
rlabel metal2 s 16882 6494 16882 6494 4 _1005_
rlabel metal2 s 16238 4726 16238 4726 4 _1006_
rlabel metal1 s 16790 18258 16790 18258 4 _1007_
rlabel metal2 s 16974 13362 16974 13362 4 _1008_
rlabel metal1 s 16606 16694 16606 16694 4 _1009_
rlabel metal1 s 21896 15402 21896 15402 4 _1010_
rlabel metal1 s 22770 15572 22770 15572 4 _1011_
rlabel metal2 s 21850 15708 21850 15708 4 _1012_
rlabel metal2 s 22586 15164 22586 15164 4 _1013_
rlabel metal1 s 17618 12750 17618 12750 4 _1014_
rlabel metal1 s 17342 12410 17342 12410 4 _1015_
rlabel metal1 s 17204 12614 17204 12614 4 _1016_
rlabel metal2 s 16882 12070 16882 12070 4 _1017_
rlabel metal1 s 16698 12240 16698 12240 4 _1018_
rlabel metal3 s 13662 7293 13662 7293 4 _1019_
rlabel metal2 s 16146 6783 16146 6783 4 _1020_
rlabel metal1 s 17020 4590 17020 4590 4 _1021_
rlabel metal2 s 17250 5100 17250 5100 4 _1022_
rlabel metal2 s 17066 3468 17066 3468 4 _1023_
rlabel metal2 s 17158 1836 17158 1836 4 _1024_
rlabel metal1 s 11316 11662 11316 11662 4 _1025_
rlabel metal1 s 15870 14994 15870 14994 4 _1026_
rlabel metal1 s 18584 15130 18584 15130 4 _1027_
rlabel metal2 s 16238 14314 16238 14314 4 _1028_
rlabel metal1 s 15042 16694 15042 16694 4 _1029_
rlabel metal1 s 17204 15538 17204 15538 4 _1030_
rlabel metal1 s 15410 17068 15410 17068 4 _1031_
rlabel metal2 s 15594 16796 15594 16796 4 _1032_
rlabel metal1 s 15686 16626 15686 16626 4 _1033_
rlabel metal1 s 16008 13838 16008 13838 4 _1034_
rlabel metal1 s 16284 13906 16284 13906 4 _1035_
rlabel metal1 s 16238 10608 16238 10608 4 _1036_
rlabel metal1 s 16054 10234 16054 10234 4 _1037_
rlabel metal2 s 16280 10404 16280 10404 4 _1038_
rlabel metal1 s 9614 14892 9614 14892 4 _1039_
rlabel metal1 s 16054 6290 16054 6290 4 _1040_
rlabel metal2 s 18722 8279 18722 8279 4 _1041_
rlabel metal1 s 17434 6324 17434 6324 4 _1042_
rlabel metal1 s 16422 6324 16422 6324 4 _1043_
rlabel metal1 s 16146 3570 16146 3570 4 _1044_
rlabel metal1 s 16606 3536 16606 3536 4 _1045_
rlabel metal1 s 16008 3366 16008 3366 4 _1046_
rlabel metal2 s 15689 1530 15689 1530 4 _1047_
rlabel metal1 s 16008 7854 16008 7854 4 _1048_
rlabel metal1 s 14812 4590 14812 4590 4 _1049_
rlabel metal1 s 13846 4488 13846 4488 4 _1050_
rlabel metal1 s 14122 10778 14122 10778 4 _1051_
rlabel metal1 s 16698 14994 16698 14994 4 _1052_
rlabel metal1 s 13938 12274 13938 12274 4 _1053_
rlabel metal1 s 13156 12206 13156 12206 4 _1054_
rlabel metal2 s 13846 11866 13846 11866 4 _1055_
rlabel metal2 s 14398 16864 14398 16864 4 _1056_
rlabel metal1 s 12834 16660 12834 16660 4 _1057_
rlabel metal1 s 12604 16626 12604 16626 4 _1058_
rlabel metal1 s 12696 16082 12696 16082 4 _1059_
rlabel metal2 s 13018 16286 13018 16286 4 _1060_
rlabel metal1 s 13754 11696 13754 11696 4 _1061_
rlabel metal2 s 14490 11356 14490 11356 4 _1062_
rlabel metal1 s 14306 11186 14306 11186 4 _1063_
rlabel metal1 s 13662 11152 13662 11152 4 _1064_
rlabel metal1 s 13340 4658 13340 4658 4 _1065_
rlabel metal1 s 14352 4114 14352 4114 4 _1066_
rlabel metal1 s 14720 3706 14720 3706 4 _1067_
rlabel metal1 s 14858 1462 14858 1462 4 _1068_
rlabel metal1 s 14766 986 14766 986 4 _1069_
rlabel metal2 s 20470 2057 20470 2057 4 _1070_
rlabel metal2 s 14674 6528 14674 6528 4 _1071_
rlabel metal1 s 14628 6358 14628 6358 4 _1072_
rlabel metal1 s 11454 9520 11454 9520 4 _1073_
rlabel metal1 s 21206 8806 21206 8806 4 _1074_
rlabel metal2 s 11362 9316 11362 9316 4 _1075_
rlabel metal1 s 11914 6086 11914 6086 4 _1076_
rlabel metal1 s 7130 9350 7130 9350 4 _1077_
rlabel metal1 s 5520 9486 5520 9486 4 _1078_
rlabel metal2 s 5658 9690 5658 9690 4 _1079_
rlabel metal2 s 6302 9316 6302 9316 4 _1080_
rlabel metal1 s 12880 13158 12880 13158 4 _1081_
rlabel metal2 s 12834 11305 12834 11305 4 _1082_
rlabel metal1 s 7360 10098 7360 10098 4 _1083_
rlabel metal1 s 3910 12682 3910 12682 4 _1084_
rlabel metal1 s 4508 9418 4508 9418 4 _1085_
rlabel metal1 s 4324 9146 4324 9146 4 _1086_
rlabel metal1 s 4462 9520 4462 9520 4 _1087_
rlabel metal1 s 4646 9010 4646 9010 4 _1088_
rlabel metal1 s 7176 10098 7176 10098 4 _1089_
rlabel metal1 s 7084 9554 7084 9554 4 _1090_
rlabel metal1 s 7590 9622 7590 9622 4 _1091_
rlabel metal1 s 11776 6290 11776 6290 4 _1092_
rlabel metal4 s 12581 11492 12581 11492 4 _1093_
rlabel metal2 s 12466 6783 12466 6783 4 _1094_
rlabel metal2 s 11546 5916 11546 5916 4 _1095_
rlabel metal1 s 19366 5032 19366 5032 4 _1096_
rlabel metal1 s 11638 2516 11638 2516 4 _1097_
rlabel metal1 s 13064 2278 13064 2278 4 _1098_
rlabel metal2 s 11546 2074 11546 2074 4 _1099_
rlabel metal1 s 11592 918 11592 918 4 _1100_
rlabel metal1 s 21390 8262 21390 8262 4 _1101_
rlabel metal1 s 13800 8534 13800 8534 4 _1102_
rlabel metal2 s 12650 9384 12650 9384 4 _1103_
rlabel metal2 s 12466 8228 12466 8228 4 _1104_
rlabel metal1 s 13018 6970 13018 6970 4 _1105_
rlabel metal2 s 6302 7344 6302 7344 4 _1106_
rlabel metal2 s 5566 3808 5566 3808 4 _1107_
rlabel metal2 s 5842 2448 5842 2448 4 _1108_
rlabel metal1 s 6302 1870 6302 1870 4 _1109_
rlabel metal1 s 6164 1938 6164 1938 4 _1110_
rlabel metal1 s 6716 6086 6716 6086 4 _1111_
rlabel metal1 s 3220 12750 3220 12750 4 _1112_
rlabel metal1 s 3634 6256 3634 6256 4 _1113_
rlabel metal1 s 4830 6256 4830 6256 4 _1114_
rlabel metal1 s 4186 6188 4186 6188 4 _1115_
rlabel metal2 s 4094 6307 4094 6307 4 _1116_
rlabel metal1 s 6946 6188 6946 6188 4 _1117_
rlabel metal1 s 6394 6766 6394 6766 4 _1118_
rlabel metal1 s 6210 6426 6210 6426 4 _1119_
rlabel metal3 s 13938 6749 13938 6749 4 _1120_
rlabel metal1 s 13984 6834 13984 6834 4 _1121_
rlabel metal2 s 12834 5338 12834 5338 4 _1122_
rlabel metal2 s 13018 2652 13018 2652 4 _1123_
rlabel metal1 s 13524 1258 13524 1258 4 _1124_
rlabel metal1 s 10902 6834 10902 6834 4 _1125_
rlabel metal1 s 9522 4556 9522 4556 4 _1126_
rlabel metal1 s 8602 4488 8602 4488 4 _1127_
rlabel metal1 s 4462 2550 4462 2550 4 _1128_
rlabel metal1 s 3542 2278 3542 2278 4 _1129_
rlabel metal1 s 3726 2516 3726 2516 4 _1130_
rlabel metal1 s 4278 2414 4278 2414 4 _1131_
rlabel metal1 s 4968 2618 4968 2618 4 _1132_
rlabel metal1 s 1564 5134 1564 5134 4 _1133_
rlabel metal1 s 1748 5746 1748 5746 4 _1134_
rlabel metal1 s 2024 5338 2024 5338 4 _1135_
rlabel metal2 s 1978 5916 1978 5916 4 _1136_
rlabel metal2 s 2438 5882 2438 5882 4 _1137_
rlabel metal1 s 2714 5848 2714 5848 4 _1138_
rlabel metal1 s 5980 6290 5980 6290 4 _1139_
rlabel metal1 s 5704 6426 5704 6426 4 _1140_
rlabel metal2 s 5474 6426 5474 6426 4 _1141_
rlabel metal1 s 8970 6256 8970 6256 4 _1142_
rlabel metal1 s 8326 4658 8326 4658 4 _1143_
rlabel metal1 s 8786 3060 8786 3060 4 _1144_
rlabel metal1 s 8510 3026 8510 3026 4 _1145_
rlabel metal2 s 8510 2652 8510 2652 4 _1146_
rlabel metal2 s 8786 2176 8786 2176 4 _1147_
rlabel metal1 s 2208 12682 2208 12682 4 _1148_
rlabel metal1 s 8970 8398 8970 8398 4 _1149_
rlabel metal2 s 9890 5236 9890 5236 4 _1150_
rlabel metal1 s 6379 7310 6379 7310 4 _1151_
rlabel metal2 s 2070 8874 2070 8874 4 _1152_
rlabel metal2 s 6946 8364 6946 8364 4 _1153_
rlabel metal1 s 3312 2958 3312 2958 4 _1154_
rlabel metal1 s 1840 2958 1840 2958 4 _1155_
rlabel metal1 s 1288 5746 1288 5746 4 _1156_
rlabel metal1 s 1886 8058 1886 8058 4 _1157_
rlabel metal1 s 1426 12682 1426 12682 4 _1158_
rlabel metal2 s 874 6698 874 6698 4 _1159_
rlabel metal1 s 1886 3060 1886 3060 4 _1160_
rlabel metal1 s 2553 3094 2553 3094 4 _1161_
rlabel metal1 s 3864 3094 3864 3094 4 _1162_
rlabel metal1 s 8694 6732 8694 6732 4 _1163_
rlabel metal2 s 7406 18037 7406 18037 4 _1164_
rlabel metal2 s 8786 8058 8786 8058 4 _1165_
rlabel metal1 s 9568 3570 9568 3570 4 _1166_
rlabel metal1 s 10120 3366 10120 3366 4 _1167_
rlabel metal2 s 9430 1836 9430 1836 4 _1168_
rlabel metal1 s 17848 2618 17848 2618 4 _1169_
rlabel metal1 s 18354 4624 18354 4624 4 _1170_
rlabel metal3 s 21114 9605 21114 9605 4 _1171_
rlabel metal1 s 22034 7446 22034 7446 4 _1172_
rlabel metal2 s 22310 7548 22310 7548 4 _1173_
rlabel metal2 s 21942 6783 21942 6783 4 _1174_
rlabel metal1 s 17112 15470 17112 15470 4 _1175_
rlabel metal2 s 17710 14790 17710 14790 4 _1176_
rlabel metal1 s 17480 14790 17480 14790 4 _1177_
rlabel metal1 s 15318 17612 15318 17612 4 _1178_
rlabel metal1 s 15042 17646 15042 17646 4 _1179_
rlabel metal1 s 16330 17748 16330 17748 4 _1180_
rlabel metal1 s 16652 17646 16652 17646 4 _1181_
rlabel metal2 s 17848 14926 17848 14926 4 _1182_
rlabel metal1 s 18170 11322 18170 11322 4 _1183_
rlabel metal1 s 17710 10778 17710 10778 4 _1184_
rlabel metal2 s 17434 9180 17434 9180 4 _1185_
rlabel metal2 s 17342 8007 17342 8007 4 _1186_
rlabel metal1 s 9936 22746 9936 22746 4 b6
rlabel metal2 s 11822 23511 11822 23511 4 b7
rlabel metal2 s 5934 500 5934 500 4 b[0]
rlabel metal2 s 5198 636 5198 636 4 b[1]
rlabel metal2 s 4434 0 4490 400 4 b[2]
port 7 nsew
rlabel metal2 s 3726 500 3726 500 4 b[3]
rlabel metal2 s 2990 772 2990 772 4 b[4]
rlabel metal2 s 2254 942 2254 942 4 b[5]
rlabel metal2 s 1518 500 1518 500 4 b[6]
rlabel metal2 s 782 942 782 942 4 b[7]
rlabel metal2 s 5566 534 5566 534 4 bn[0]
rlabel metal2 s 4830 500 4830 500 4 bn[1]
rlabel metal2 s 4094 636 4094 636 4 bn[2]
rlabel metal2 s 3358 670 3358 670 4 bn[3]
rlabel metal2 s 2622 636 2622 636 4 bn[4]
rlabel metal2 s 1886 500 1886 500 4 bn[5]
rlabel metal2 s 1150 500 1150 500 4 bn[6]
rlabel metal2 s 414 483 414 483 4 bn[7]
rlabel metal2 s 13294 17901 13294 17901 4 clk
rlabel metal1 s 19458 17136 19458 17136 4 clknet_0_clk
rlabel metal1 s 1288 13838 1288 13838 4 clknet_3_0__leaf_clk
rlabel metal1 s 966 16694 966 16694 4 clknet_3_1__leaf_clk
rlabel metal1 s 2254 21556 2254 21556 4 clknet_3_2__leaf_clk
rlabel metal1 s 10258 20026 10258 20026 4 clknet_3_3__leaf_clk
rlabel metal2 s 16146 18768 16146 18768 4 clknet_3_4__leaf_clk
rlabel metal1 s 21574 12750 21574 12750 4 clknet_3_5__leaf_clk
rlabel metal1 s 14950 19278 14950 19278 4 clknet_3_6__leaf_clk
rlabel metal1 s 22586 22542 22586 22542 4 clknet_3_7__leaf_clk
rlabel metal1 s 20930 17646 20930 17646 4 divider\[0\]
rlabel metal1 s 20746 17034 20746 17034 4 divider\[1\]
rlabel metal1 s 10304 23290 10304 23290 4 g6
rlabel metal1 s 12926 21930 12926 21930 4 g7
rlabel metal2 s 14766 636 14766 636 4 g[0]
rlabel metal2 s 14030 500 14030 500 4 g[1]
rlabel metal2 s 13294 500 13294 500 4 g[2]
rlabel metal2 s 12558 500 12558 500 4 g[3]
rlabel metal2 s 11822 500 11822 500 4 g[4]
rlabel metal2 s 11086 415 11086 415 4 g[5]
rlabel metal2 s 10322 0 10378 400 4 g[6]
port 30 nsew
rlabel metal2 s 9614 636 9614 636 4 g[7]
rlabel metal1 s 23138 16762 23138 16762 4 gate
rlabel metal2 s 14398 534 14398 534 4 gn[0]
rlabel metal2 s 13662 500 13662 500 4 gn[1]
rlabel metal2 s 12926 500 12926 500 4 gn[2]
rlabel metal2 s 12190 500 12190 500 4 gn[3]
rlabel metal2 s 11454 500 11454 500 4 gn[4]
rlabel metal2 s 10690 0 10746 400 4 gn[5]
port 37 nsew
rlabel metal2 s 9982 670 9982 670 4 gn[6]
rlabel metal2 s 9246 1044 9246 1044 4 gn[7]
rlabel metal1 s 8234 23290 8234 23290 4 hblank
rlabel metal2 s 9522 23239 9522 23239 4 hsync
rlabel metal1 s 21390 11696 21390 11696 4 mode\[0\]
rlabel metal1 s 22448 12614 22448 12614 4 mode\[1\]
rlabel metal1 s 20884 18054 20884 18054 4 mode\[2\]
rlabel metal1 s 20286 17646 20286 17646 4 net1
rlabel metal2 s 1886 1700 1886 1700 4 net10
rlabel metal1 s 1058 1836 1058 1836 4 net11
rlabel metal1 s 5658 816 5658 816 4 net12
rlabel metal2 s 4922 1258 4922 1258 4 net13
rlabel metal2 s 4186 1258 4186 1258 4 net14
rlabel metal1 s 3220 782 3220 782 4 net15
rlabel metal2 s 2806 1564 2806 1564 4 net16
rlabel metal1 s 2254 1394 2254 1394 4 net17
rlabel metal1 s 1702 782 1702 782 4 net18
rlabel metal1 s 690 1394 690 1394 4 net19
rlabel metal1 s 21574 3604 21574 3604 4 net2
rlabel metal2 s 21666 1343 21666 1343 4 net20
rlabel metal2 s 18630 1003 18630 1003 4 net21
rlabel metal1 s 3818 748 3818 748 4 net22
rlabel metal1 s 2714 748 2714 748 4 net23
rlabel metal1 s 2346 816 2346 816 4 net24
rlabel metal2 s 1978 476 1978 476 4 net25
rlabel metal2 s 1242 578 1242 578 4 net26
rlabel metal1 s 1518 1428 1518 1428 4 net27
rlabel metal1 s 7912 1258 7912 1258 4 net28
rlabel metal3 s 12558 21845 12558 21845 4 net29
rlabel metal3 s 21574 18037 21574 18037 4 net3
rlabel metal1 s 15778 782 15778 782 4 net30
rlabel metal2 s 14674 1258 14674 1258 4 net31
rlabel metal2 s 13846 986 13846 986 4 net32
rlabel metal2 s 12650 1258 12650 1258 4 net33
rlabel metal2 s 11914 1326 11914 1326 4 net34
rlabel metal2 s 10166 986 10166 986 4 net35
rlabel metal1 s 9430 714 9430 714 4 net36
rlabel metal1 s 8694 850 8694 850 4 net37
rlabel metal1 s 15962 816 15962 816 4 net38
rlabel metal1 s 14352 782 14352 782 4 net39
rlabel metal2 s 19550 20128 19550 20128 4 net4
rlabel metal1 s 13846 1394 13846 1394 4 net40
rlabel metal1 s 12558 748 12558 748 4 net41
rlabel metal2 s 11592 714 11592 714 4 net42
rlabel metal1 s 10120 1394 10120 1394 4 net43
rlabel metal1 s 8970 782 8970 782 4 net44
rlabel metal1 s 9292 1530 9292 1530 4 net45
rlabel metal1 s 18906 19788 18906 19788 4 net46
rlabel metal1 s 9062 21590 9062 21590 4 net47
rlabel metal2 s 18722 1921 18722 1921 4 net48
rlabel metal3 s 14214 1003 14214 1003 4 net49
rlabel metal2 s 20746 17663 20746 17663 4 net5
rlabel metal1 s 22678 2992 22678 2992 4 net50
rlabel metal2 s 22770 3162 22770 3162 4 net51
rlabel metal2 s 22356 1938 22356 1938 4 net52
rlabel metal2 s 17710 510 17710 510 4 net53
rlabel metal1 s 21666 748 21666 748 4 net54
rlabel metal2 s 20746 901 20746 901 4 net55
rlabel metal1 s 19366 782 19366 782 4 net56
rlabel metal1 s 18722 748 18722 748 4 net57
rlabel metal2 s 22034 2057 22034 2057 4 net58
rlabel metal1 s 22816 1462 22816 1462 4 net59
rlabel metal2 s 20470 18105 20470 18105 4 net6
rlabel metal2 s 19918 1632 19918 1632 4 net60
rlabel metal1 s 19090 884 19090 884 4 net61
rlabel metal1 s 21298 816 21298 816 4 net62
rlabel metal2 s 20378 986 20378 986 4 net63
rlabel metal2 s 19090 1292 19090 1292 4 net64
rlabel metal1 s 18170 816 18170 816 4 net65
rlabel metal3 s 19550 5763 19550 5763 4 net66
rlabel metal1 s 9522 22678 9522 22678 4 net67
rlabel metal1 s 7360 22474 7360 22474 4 net68
rlabel metal1 s 17664 22474 17664 22474 4 net69
rlabel metal1 s 20470 19312 20470 19312 4 net7
rlabel metal1 s 14812 22542 14812 22542 4 net70
rlabel metal1 s 7544 18802 7544 18802 4 net71
rlabel metal2 s 19918 18683 19918 18683 4 net8
rlabel metal3 s 18032 21556 18032 21556 4 net9
rlabel metal1 s 10856 23290 10856 23290 4 r6
rlabel metal1 s 13340 21930 13340 21930 4 r7
rlabel metal1 s 23046 3094 23046 3094 4 r[0]
rlabel metal1 s 22908 2822 22908 2822 4 r[1]
rlabel metal2 s 22126 1180 22126 1180 4 r[2]
rlabel metal2 s 21390 500 21390 500 4 r[3]
rlabel metal2 s 20654 415 20654 415 4 r[4]
rlabel metal2 s 19890 0 19946 400 4 r[5]
port 49 nsew
rlabel metal2 s 19182 636 19182 636 4 r[6]
rlabel metal2 s 18446 500 18446 500 4 r[7]
rlabel metal2 s 23046 10778 23046 10778 4 registered
rlabel metal2 s 23230 1112 23230 1112 4 rn[0]
rlabel metal2 s 22466 0 22522 400 4 rn[1]
port 53 nsew
rlabel metal2 s 21758 636 21758 636 4 rn[2]
rlabel metal2 s 21022 636 21022 636 4 rn[3]
rlabel metal2 s 20258 0 20314 400 4 rn[4]
port 56 nsew
rlabel metal2 s 19550 534 19550 534 4 rn[5]
rlabel metal2 s 18814 534 18814 534 4 rn[6]
rlabel metal2 s 18078 500 18078 500 4 rn[7]
rlabel metal2 s 22954 22933 22954 22933 4 rst_n
rlabel metal1 s 22264 20774 22264 20774 4 ui_in[0]
rlabel metal2 s 21574 23470 21574 23470 4 ui_in[1]
rlabel metal1 s 21252 21046 21252 21046 4 ui_in[2]
rlabel metal2 s 20286 23443 20286 23443 4 ui_in[3]
rlabel metal2 s 19918 22586 19918 22586 4 ui_in[4]
rlabel metal1 s 21206 22576 21206 22576 4 ui_in[5]
rlabel metal1 s 18584 23222 18584 23222 4 ui_in[6]
rlabel metal1 s 17342 23222 17342 23222 4 ui_in[7]
rlabel metal1 s 8970 21658 8970 21658 4 vblank
rlabel metal1 s 13386 16694 13386 16694 4 vga_sync.hpos\[0\]
rlabel metal2 s 19918 17000 19918 17000 4 vga_sync.hpos\[1\]
rlabel metal1 s 14674 17136 14674 17136 4 vga_sync.hpos\[2\]
rlabel metal1 s 10350 16048 10350 16048 4 vga_sync.hpos\[3\]
rlabel metal2 s 7130 15980 7130 15980 4 vga_sync.hpos\[4\]
rlabel metal3 s 3358 15453 3358 15453 4 vga_sync.hpos\[5\]
rlabel metal2 s 2346 18122 2346 18122 4 vga_sync.hpos\[6\]
rlabel metal2 s 4186 18054 4186 18054 4 vga_sync.hpos\[7\]
rlabel metal2 s 5014 15657 5014 15657 4 vga_sync.hpos\[8\]
rlabel metal2 s 2346 16320 2346 16320 4 vga_sync.hpos\[9\]
rlabel metal2 s 8280 19142 8280 19142 4 vga_sync.hsync
rlabel metal1 s 5290 19278 5290 19278 4 vga_sync.mode
rlabel metal1 s 14490 21012 14490 21012 4 vga_sync.o_vpos\[0\]
rlabel metal1 s 13018 20570 13018 20570 4 vga_sync.o_vpos\[1\]
rlabel metal1 s 14306 23154 14306 23154 4 vga_sync.o_vpos\[2\]
rlabel metal1 s 13110 22474 13110 22474 4 vga_sync.o_vpos\[3\]
rlabel metal1 s 6394 22610 6394 22610 4 vga_sync.o_vpos\[4\]
rlabel metal1 s 3864 22066 3864 22066 4 vga_sync.o_vpos\[5\]
rlabel metal1 s 2116 22066 2116 22066 4 vga_sync.o_vpos\[6\]
rlabel metal1 s 5658 19924 5658 19924 4 vga_sync.o_vpos\[7\]
rlabel metal1 s 6440 18802 6440 18802 4 vga_sync.o_vpos\[8\]
rlabel metal2 s 6486 20149 6486 20149 4 vga_sync.o_vpos\[9\]
rlabel metal2 s 8142 22780 8142 22780 4 vga_sync.vsync
rlabel metal1 s 15686 21080 15686 21080 4 voffset\[0\]
rlabel metal2 s 17526 21080 17526 21080 4 voffset\[1\]
rlabel metal1 s 16974 22440 16974 22440 4 voffset\[2\]
rlabel metal1 s 13018 22610 13018 22610 4 voffset\[3\]
rlabel metal2 s 20102 23392 20102 23392 4 voffset\[4\]
rlabel metal1 s 17296 22202 17296 22202 4 voffset\[5\]
rlabel metal2 s 2254 23392 2254 23392 4 voffset\[6\]
rlabel metal3 s 2070 20349 2070 20349 4 voffset\[7\]
rlabel metal1 s 11546 23290 11546 23290 4 vsync
rlabel metal1 s 19182 18802 19182 18802 4 xor1.t\[0\]
rlabel metal2 s 2622 13600 2622 13600 4 xor1.t\[10\]
rlabel metal2 s 1610 14620 1610 14620 4 xor1.t\[11\]
rlabel metal2 s 20102 17102 20102 17102 4 xor1.t\[1\]
rlabel metal2 s 17710 18088 17710 18088 4 xor1.t\[2\]
rlabel metal1 s 15962 18190 15962 18190 4 xor1.t\[3\]
rlabel metal2 s 15134 18938 15134 18938 4 xor1.t\[4\]
rlabel metal1 s 13478 17034 13478 17034 4 xor1.t\[5\]
rlabel metal1 s 10534 16014 10534 16014 4 xor1.t\[6\]
rlabel metal1 s 3818 12138 3818 12138 4 xor1.t\[7\]
rlabel metal1 s 2254 10642 2254 10642 4 xor1.t\[8\]
rlabel metal2 s 2162 8908 2162 8908 4 xor1.t\[9\]
flabel metal4 s 22352 496 22752 23440 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 16352 496 16752 23440 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 10352 496 10752 23440 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 4352 496 4752 23440 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 19352 496 19752 23440 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 13352 496 13752 23440 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 7352 496 7752 23440 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 1352 496 1752 23440 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal2 s 9954 23600 10010 24000 0 FreeSans 280 90 0 0 b6
port 3 nsew
flabel metal2 s 12162 23600 12218 24000 0 FreeSans 280 90 0 0 b7
port 4 nsew
flabel metal2 s 5906 0 5962 400 0 FreeSans 280 90 0 0 b[0]
port 5 nsew
flabel metal2 s 5170 0 5226 400 0 FreeSans 280 90 0 0 b[1]
port 6 nsew
flabel metal2 s 4462 200 4462 200 0 FreeSans 280 90 0 0 b[2]
flabel metal2 s 3698 0 3754 400 0 FreeSans 280 90 0 0 b[3]
port 8 nsew
flabel metal2 s 2962 0 3018 400 0 FreeSans 280 90 0 0 b[4]
port 9 nsew
flabel metal2 s 2226 0 2282 400 0 FreeSans 280 90 0 0 b[5]
port 10 nsew
flabel metal2 s 1490 0 1546 400 0 FreeSans 280 90 0 0 b[6]
port 11 nsew
flabel metal2 s 754 0 810 400 0 FreeSans 280 90 0 0 b[7]
port 12 nsew
flabel metal2 s 5538 0 5594 400 0 FreeSans 280 90 0 0 bn[0]
port 13 nsew
flabel metal2 s 4802 0 4858 400 0 FreeSans 280 90 0 0 bn[1]
port 14 nsew
flabel metal2 s 4066 0 4122 400 0 FreeSans 280 90 0 0 bn[2]
port 15 nsew
flabel metal2 s 3330 0 3386 400 0 FreeSans 280 90 0 0 bn[3]
port 16 nsew
flabel metal2 s 2594 0 2650 400 0 FreeSans 280 90 0 0 bn[4]
port 17 nsew
flabel metal2 s 1858 0 1914 400 0 FreeSans 280 90 0 0 bn[5]
port 18 nsew
flabel metal2 s 1122 0 1178 400 0 FreeSans 280 90 0 0 bn[6]
port 19 nsew
flabel metal2 s 386 0 442 400 0 FreeSans 280 90 0 0 bn[7]
port 20 nsew
flabel metal2 s 23202 23600 23258 24000 0 FreeSans 280 90 0 0 clk
port 21 nsew
flabel metal2 s 10506 23600 10562 24000 0 FreeSans 280 90 0 0 g6
port 22 nsew
flabel metal2 s 12714 23600 12770 24000 0 FreeSans 280 90 0 0 g7
port 23 nsew
flabel metal2 s 14738 0 14794 400 0 FreeSans 280 90 0 0 g[0]
port 24 nsew
flabel metal2 s 14002 0 14058 400 0 FreeSans 280 90 0 0 g[1]
port 25 nsew
flabel metal2 s 13266 0 13322 400 0 FreeSans 280 90 0 0 g[2]
port 26 nsew
flabel metal2 s 12530 0 12586 400 0 FreeSans 280 90 0 0 g[3]
port 27 nsew
flabel metal2 s 11794 0 11850 400 0 FreeSans 280 90 0 0 g[4]
port 28 nsew
flabel metal2 s 11058 0 11114 400 0 FreeSans 280 90 0 0 g[5]
port 29 nsew
flabel metal2 s 10350 200 10350 200 0 FreeSans 280 90 0 0 g[6]
flabel metal2 s 9586 0 9642 400 0 FreeSans 280 90 0 0 g[7]
port 31 nsew
flabel metal2 s 14370 0 14426 400 0 FreeSans 280 90 0 0 gn[0]
port 32 nsew
flabel metal2 s 13634 0 13690 400 0 FreeSans 280 90 0 0 gn[1]
port 33 nsew
flabel metal2 s 12898 0 12954 400 0 FreeSans 280 90 0 0 gn[2]
port 34 nsew
flabel metal2 s 12162 0 12218 400 0 FreeSans 280 90 0 0 gn[3]
port 35 nsew
flabel metal2 s 11426 0 11482 400 0 FreeSans 280 90 0 0 gn[4]
port 36 nsew
flabel metal2 s 10718 200 10718 200 0 FreeSans 280 90 0 0 gn[5]
flabel metal2 s 9954 0 10010 400 0 FreeSans 280 90 0 0 gn[6]
port 38 nsew
flabel metal2 s 9218 0 9274 400 0 FreeSans 280 90 0 0 gn[7]
port 39 nsew
flabel metal2 s 8298 23600 8354 24000 0 FreeSans 280 90 0 0 hblank
port 40 nsew
flabel metal2 s 9402 23600 9458 24000 0 FreeSans 280 90 0 0 hsync
port 41 nsew
flabel metal2 s 11058 23600 11114 24000 0 FreeSans 280 90 0 0 r6
port 42 nsew
flabel metal2 s 13266 23600 13322 24000 0 FreeSans 280 90 0 0 r7
port 43 nsew
flabel metal2 s 23570 0 23626 400 0 FreeSans 280 90 0 0 r[0]
port 44 nsew
flabel metal2 s 22834 0 22890 400 0 FreeSans 280 90 0 0 r[1]
port 45 nsew
flabel metal2 s 22098 0 22154 400 0 FreeSans 280 90 0 0 r[2]
port 46 nsew
flabel metal2 s 21362 0 21418 400 0 FreeSans 280 90 0 0 r[3]
port 47 nsew
flabel metal2 s 20626 0 20682 400 0 FreeSans 280 90 0 0 r[4]
port 48 nsew
flabel metal2 s 19918 200 19918 200 0 FreeSans 280 90 0 0 r[5]
flabel metal2 s 19154 0 19210 400 0 FreeSans 280 90 0 0 r[6]
port 50 nsew
flabel metal2 s 18418 0 18474 400 0 FreeSans 280 90 0 0 r[7]
port 51 nsew
flabel metal2 s 23202 0 23258 400 0 FreeSans 280 90 0 0 rn[0]
port 52 nsew
flabel metal2 s 22494 200 22494 200 0 FreeSans 280 90 0 0 rn[1]
flabel metal2 s 21730 0 21786 400 0 FreeSans 280 90 0 0 rn[2]
port 54 nsew
flabel metal2 s 20994 0 21050 400 0 FreeSans 280 90 0 0 rn[3]
port 55 nsew
flabel metal2 s 20286 200 20286 200 0 FreeSans 280 90 0 0 rn[4]
flabel metal2 s 19522 0 19578 400 0 FreeSans 280 90 0 0 rn[5]
port 57 nsew
flabel metal2 s 18786 0 18842 400 0 FreeSans 280 90 0 0 rn[6]
port 58 nsew
flabel metal2 s 18050 0 18106 400 0 FreeSans 280 90 0 0 rn[7]
port 59 nsew
flabel metal2 s 22650 23600 22706 24000 0 FreeSans 280 90 0 0 rst_n
port 60 nsew
flabel metal2 s 22098 23600 22154 24000 0 FreeSans 280 90 0 0 ui_in[0]
port 61 nsew
flabel metal2 s 21546 23600 21602 24000 0 FreeSans 280 90 0 0 ui_in[1]
port 62 nsew
flabel metal2 s 20994 23600 21050 24000 0 FreeSans 280 90 0 0 ui_in[2]
port 63 nsew
flabel metal2 s 20442 23600 20498 24000 0 FreeSans 280 90 0 0 ui_in[3]
port 64 nsew
flabel metal2 s 19890 23600 19946 24000 0 FreeSans 280 90 0 0 ui_in[4]
port 65 nsew
flabel metal2 s 19338 23600 19394 24000 0 FreeSans 280 90 0 0 ui_in[5]
port 66 nsew
flabel metal2 s 18786 23600 18842 24000 0 FreeSans 280 90 0 0 ui_in[6]
port 67 nsew
flabel metal2 s 18234 23600 18290 24000 0 FreeSans 280 90 0 0 ui_in[7]
port 68 nsew
flabel metal2 s 8850 23600 8906 24000 0 FreeSans 280 90 0 0 vblank
port 69 nsew
flabel metal2 s 11610 23600 11666 24000 0 FreeSans 280 90 0 0 vsync
port 70 nsew
<< properties >>
string FIXED_BBOX 0 0 24000 24000
string GDS_END 3601306
string GDS_FILE ../gds/controller.gds
string GDS_START 435046
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1723601757
<< error_s >>
rect 11230 -7470 11239 -7461
rect 11421 -7470 11430 -7461
rect 11221 -7479 11230 -7470
rect 11430 -7479 11439 -7470
rect 11221 -7670 11230 -7661
rect 11430 -7670 11439 -7661
rect 11230 -7679 11239 -7670
rect 11421 -7679 11430 -7670
rect 5053 -8814 5088 -8780
rect 5054 -8833 5088 -8814
rect 4884 -8882 4942 -8876
rect 4884 -8916 4896 -8882
rect 4884 -8922 4942 -8916
rect 4884 -9092 4942 -9086
rect 4884 -9126 4896 -9092
rect 4884 -9132 4942 -9126
rect 5073 -9228 5088 -8833
rect 5107 -8867 5142 -8833
rect 5422 -8867 5457 -8833
rect 5107 -9228 5141 -8867
rect 5423 -8886 5457 -8867
rect 5253 -8935 5311 -8929
rect 5253 -8969 5265 -8935
rect 5253 -8975 5311 -8969
rect 5253 -9145 5311 -9139
rect 5253 -9179 5265 -9145
rect 5253 -9185 5311 -9179
rect 5107 -9262 5122 -9228
rect 5442 -9281 5457 -8886
rect 5476 -8920 5511 -8886
rect 7361 -8920 7396 -8886
rect 5476 -9281 5510 -8920
rect 7362 -8939 7396 -8920
rect 5476 -9315 5491 -9281
rect 7381 -9334 7396 -8939
rect 7415 -8973 7450 -8939
rect 7730 -8973 7765 -8939
rect 7415 -9334 7449 -8973
rect 7731 -8992 7765 -8973
rect 7561 -9041 7619 -9035
rect 7561 -9075 7573 -9041
rect 7561 -9081 7619 -9075
rect 7561 -9251 7619 -9245
rect 7561 -9285 7573 -9251
rect 7561 -9291 7619 -9285
rect 7415 -9368 7430 -9334
rect 7750 -9387 7765 -8992
rect 7784 -9026 7819 -8992
rect 8099 -9026 8134 -8992
rect 7784 -9387 7818 -9026
rect 8100 -9045 8134 -9026
rect 7930 -9094 7988 -9088
rect 7930 -9128 7942 -9094
rect 7930 -9134 7988 -9128
rect 7930 -9304 7988 -9298
rect 7930 -9338 7942 -9304
rect 7930 -9344 7988 -9338
rect 7784 -9421 7799 -9387
rect 8119 -9440 8134 -9045
rect 8153 -9079 8188 -9045
rect 9238 -9079 9273 -9045
rect 8153 -9440 8187 -9079
rect 9239 -9098 9273 -9079
rect 8153 -9474 8168 -9440
rect 9258 -9493 9273 -9098
rect 9292 -9132 9327 -9098
rect 9607 -9132 9642 -9098
rect 9292 -9493 9326 -9132
rect 9608 -9151 9642 -9132
rect 9438 -9200 9496 -9194
rect 9438 -9234 9450 -9200
rect 9438 -9240 9496 -9234
rect 9438 -9410 9496 -9404
rect 9438 -9444 9450 -9410
rect 9438 -9450 9496 -9444
rect 9292 -9527 9307 -9493
rect 9627 -9546 9642 -9151
rect 9661 -9185 9696 -9151
rect 9976 -9185 10011 -9151
rect 9661 -9546 9695 -9185
rect 9977 -9204 10011 -9185
rect 9807 -9253 9865 -9247
rect 9807 -9287 9819 -9253
rect 9807 -9293 9865 -9287
rect 9807 -9463 9865 -9457
rect 9807 -9497 9819 -9463
rect 9807 -9503 9865 -9497
rect 9661 -9580 9676 -9546
rect 9996 -9599 10011 -9204
rect 10030 -9238 10065 -9204
rect 10735 -9238 10770 -9204
rect 10030 -9599 10064 -9238
rect 10736 -9257 10770 -9238
rect 10030 -9633 10045 -9599
rect 10755 -9652 10770 -9257
rect 10789 -9291 10824 -9257
rect 11104 -9291 11139 -9257
rect 10789 -9652 10823 -9291
rect 11105 -9310 11139 -9291
rect 10935 -9359 10993 -9353
rect 10935 -9393 10947 -9359
rect 10935 -9399 10993 -9393
rect 10935 -9569 10993 -9563
rect 10935 -9603 10947 -9569
rect 10935 -9609 10993 -9603
rect 10789 -9686 10804 -9652
rect 11124 -9705 11139 -9310
rect 11158 -9344 11193 -9310
rect 11473 -9344 11508 -9310
rect 11158 -9705 11192 -9344
rect 11474 -9363 11508 -9344
rect 11304 -9412 11362 -9406
rect 11304 -9446 11316 -9412
rect 11304 -9452 11362 -9446
rect 11304 -9622 11362 -9616
rect 11304 -9656 11316 -9622
rect 11304 -9662 11362 -9656
rect 11158 -9739 11173 -9705
rect 11493 -9758 11508 -9363
rect 11527 -9397 11562 -9363
rect 12012 -9397 12047 -9363
rect 11527 -9758 11561 -9397
rect 12013 -9416 12047 -9397
rect 11527 -9792 11542 -9758
rect 12032 -9811 12047 -9416
rect 12066 -9450 12101 -9416
rect 12381 -9450 12416 -9416
rect 12066 -9811 12100 -9450
rect 12382 -9469 12416 -9450
rect 12212 -9518 12270 -9512
rect 12212 -9552 12224 -9518
rect 12212 -9558 12270 -9552
rect 12212 -9728 12270 -9722
rect 12212 -9762 12224 -9728
rect 12212 -9768 12270 -9762
rect 12066 -9845 12081 -9811
rect 12401 -9864 12416 -9469
rect 12435 -9503 12470 -9469
rect 12435 -9864 12469 -9503
rect 12581 -9571 12639 -9565
rect 12581 -9605 12593 -9571
rect 12581 -9611 12639 -9605
rect 12581 -9781 12639 -9775
rect 12581 -9815 12593 -9781
rect 12581 -9821 12639 -9815
rect 12435 -9898 12450 -9864
rect 12770 -9917 12785 -9469
rect 12804 -9917 12838 -9415
rect 13550 -9475 13584 -9421
rect 16272 -9427 16307 -9393
rect 15095 -9468 15130 -9434
rect 16273 -9446 16307 -9427
rect 12804 -9951 12819 -9917
rect 13569 -9970 13584 -9475
rect 13603 -9509 13638 -9475
rect 13918 -9509 13953 -9475
rect 15096 -9487 15130 -9468
rect 13603 -9970 13637 -9509
rect 13919 -9528 13953 -9509
rect 13749 -9577 13807 -9571
rect 13749 -9611 13761 -9577
rect 13749 -9617 13807 -9611
rect 13749 -9887 13807 -9881
rect 13749 -9921 13761 -9887
rect 13749 -9927 13807 -9921
rect 13603 -10004 13618 -9970
rect 13938 -10023 13953 -9528
rect 13972 -9562 14007 -9528
rect 14287 -9561 14322 -9528
rect 13972 -10023 14006 -9562
rect 14118 -9630 14176 -9624
rect 14118 -9664 14130 -9630
rect 14118 -9670 14176 -9664
rect 14118 -9940 14176 -9934
rect 14118 -9974 14130 -9940
rect 14118 -9980 14176 -9974
rect 13972 -10057 13987 -10023
rect 14307 -10076 14322 -9561
rect 14341 -9595 14376 -9561
rect 14341 -10076 14375 -9595
rect 14341 -10110 14356 -10076
rect 14746 -10129 14761 -9561
rect 14780 -10129 14814 -9507
rect 14926 -9536 14984 -9530
rect 14926 -9570 14938 -9536
rect 14926 -9576 14984 -9570
rect 14926 -10046 14984 -10040
rect 14926 -10080 14938 -10046
rect 14926 -10086 14984 -10080
rect 14780 -10163 14795 -10129
rect 15115 -10182 15130 -9487
rect 15149 -9521 15184 -9487
rect 15464 -9520 15499 -9487
rect 15149 -10182 15183 -9521
rect 15295 -9589 15353 -9583
rect 15295 -9623 15307 -9589
rect 15295 -9629 15353 -9623
rect 15295 -10099 15353 -10093
rect 15295 -10133 15307 -10099
rect 15295 -10139 15353 -10133
rect 15149 -10216 15164 -10182
rect 15484 -10235 15499 -9520
rect 15518 -9554 15553 -9520
rect 15518 -10235 15552 -9554
rect 15518 -10269 15533 -10235
rect 15923 -10288 15938 -9520
rect 15957 -10288 15991 -9466
rect 16103 -9495 16161 -9489
rect 16103 -9529 16115 -9495
rect 16103 -9535 16161 -9529
rect 16103 -10205 16161 -10199
rect 16103 -10239 16115 -10205
rect 16103 -10245 16161 -10239
rect 15957 -10322 15972 -10288
rect 16292 -10341 16307 -9446
rect 16326 -9480 16361 -9446
rect 16326 -10341 16360 -9480
rect 16472 -9548 16530 -9542
rect 16472 -9582 16484 -9548
rect 16472 -9588 16530 -9582
rect 16472 -10258 16530 -10252
rect 16472 -10292 16484 -10258
rect 16472 -10298 16530 -10292
rect 16326 -10375 16341 -10341
<< viali >>
rect 940 5060 1120 5110
rect 1380 5050 1630 5100
rect 850 4720 900 5010
rect 1280 4960 1330 5010
rect 1280 4730 1330 4780
rect 1680 4730 1720 5000
rect 940 4630 1120 4680
rect 1510 4640 1630 4680
rect 8560 -6085 8630 2855
rect 9940 -6090 10080 2850
rect 11390 -6085 11460 2855
<< metal1 >>
rect 1994 5696 2194 5896
rect 2394 5696 2594 5896
rect 2794 5696 2994 5896
rect 3194 5696 3394 5896
rect 3594 5696 3794 5896
rect 3994 5696 4194 5896
rect 4394 5696 4594 5896
rect 4794 5696 4994 5896
rect 5194 5696 5394 5896
rect 5594 5696 5794 5896
rect 5994 5696 6194 5896
rect 6394 5696 6594 5896
rect 6794 5696 6994 5896
rect 7194 5696 7394 5896
rect 7594 5696 7794 5896
rect 7994 5696 8194 5896
rect 840 5110 1140 5120
rect 840 5060 940 5110
rect 1120 5060 1140 5110
rect 840 5050 1140 5060
rect 1270 5100 1730 5110
rect 1270 5050 1380 5100
rect 1630 5050 1730 5100
rect 840 5010 910 5050
rect 1270 5040 1730 5050
rect 1270 5020 1350 5040
rect 840 4720 850 5010
rect 900 4920 910 5010
rect 990 4960 1280 5020
rect 1340 4960 1350 5020
rect 1670 5000 1730 5040
rect 990 4950 1350 4960
rect 1380 4950 1560 5000
rect 1380 4920 1460 4950
rect 1670 4920 1680 5000
rect 900 4820 1010 4920
rect 1050 4820 1460 4920
rect 1560 4820 1680 4920
rect 900 4720 910 4820
rect 990 4730 1280 4790
rect 1340 4730 1350 4790
rect 990 4720 1350 4730
rect 1380 4780 1460 4820
rect 1380 4730 1560 4780
rect 1670 4730 1680 4820
rect 1720 4730 1730 5000
rect 840 4690 910 4720
rect 840 4680 1140 4690
rect 840 4630 940 4680
rect 1120 4630 1140 4680
rect 0 4000 350 4200
rect 550 4000 556 4200
rect 840 4180 1140 4630
rect 840 4020 860 4180
rect 1120 4020 1140 4180
rect 840 4000 1140 4020
rect 0 3600 350 3800
rect 550 3600 556 3800
rect 1380 3370 1460 4730
rect 1670 4690 1730 4730
rect 1490 4680 1730 4690
rect 1490 4640 1510 4680
rect 1630 4640 1730 4680
rect 1490 4630 1730 4640
rect 1540 3780 1730 4630
rect 8970 4180 9590 4200
rect 8970 4020 8990 4180
rect 9570 4020 9590 4180
rect 1540 3620 1560 3780
rect 1710 3620 1730 3780
rect 1540 3600 1730 3620
rect 8470 3780 8650 3800
rect 8470 3620 8490 3780
rect 8630 3620 8650 3780
rect 1360 3350 1480 3370
rect 1360 3220 1380 3350
rect 1460 3220 1480 3350
rect 1360 3200 1480 3220
rect 8470 2855 8650 3620
rect 8470 -6085 8560 2855
rect 8630 -6085 8650 2855
rect 8970 2820 9590 4020
rect 10430 4180 11050 4200
rect 10430 4020 10450 4180
rect 11030 4020 11050 4180
rect 9920 3780 10100 3800
rect 9920 3620 9940 3780
rect 10080 3620 10100 3780
rect 9920 2850 10100 3620
rect 8690 2350 9870 2820
rect 8680 -6060 9880 -5580
rect 8470 -6260 8650 -6085
rect 8970 -7490 9590 -6060
rect 9920 -6090 9940 2850
rect 10080 -6090 10100 2850
rect 10430 2820 11050 4020
rect 11370 3780 11550 3800
rect 11370 3620 11390 3780
rect 11530 3620 11550 3780
rect 11370 2855 11550 3620
rect 10150 2350 11330 2820
rect 10140 -6060 11340 -5580
rect 9920 -6260 10100 -6090
rect 10430 -7090 11050 -6060
rect 11370 -6085 11390 2855
rect 11460 -6085 11550 2855
rect 11370 -6260 11550 -6085
rect 11224 -6870 11230 -6670
rect 11430 -6870 11710 -6670
rect 10430 -7250 10450 -7090
rect 11030 -7250 11050 -7090
rect 10430 -7270 11050 -7250
rect 11224 -7270 11230 -7070
rect 11430 -7270 11710 -7070
rect 8970 -7650 8990 -7490
rect 9570 -7650 9590 -7490
rect 8970 -7670 9590 -7650
rect 11430 -7670 11710 -7470
<< via1 >>
rect 1280 5010 1340 5020
rect 1280 4960 1330 5010
rect 1330 4960 1340 5010
rect 1280 4780 1340 4790
rect 1280 4730 1330 4780
rect 1330 4730 1340 4780
rect 350 4000 550 4200
rect 860 4020 1120 4180
rect 350 3600 550 3800
rect 8990 4020 9570 4180
rect 1560 3620 1710 3780
rect 8490 3620 8630 3780
rect 1380 3220 1460 3350
rect 10450 4020 11030 4180
rect 9940 3620 10080 3780
rect 11390 3620 11530 3780
rect 11230 -6870 11430 -6670
rect 10450 -7250 11030 -7090
rect 11230 -7270 11430 -7070
rect 8990 -7650 9570 -7490
rect 11230 -7670 11430 -7470
<< metal2 >>
rect 1270 5020 1350 5030
rect 1270 4960 1280 5020
rect 1340 4960 1350 5020
rect 1270 4790 1350 4960
rect 1270 4730 1280 4790
rect 1340 4730 1350 4790
rect 1270 4710 1350 4730
rect 330 4200 570 4220
rect 330 4000 350 4200
rect 550 4000 570 4200
rect 840 4180 1140 4200
rect 840 4020 860 4180
rect 1120 4020 1140 4180
rect 840 4000 1140 4020
rect 8970 4180 9590 4200
rect 8970 4020 8990 4180
rect 9570 4020 9590 4180
rect 8970 4000 9590 4020
rect 10430 4180 11050 4200
rect 10430 4020 10450 4180
rect 11030 4020 11050 4180
rect 10430 4000 11050 4020
rect 330 3980 570 4000
rect 330 3800 570 3820
rect 330 3600 350 3800
rect 550 3600 570 3800
rect 1540 3780 1730 3800
rect 1540 3620 1560 3780
rect 1710 3620 1730 3780
rect 1540 3600 1730 3620
rect 8470 3780 8650 3800
rect 8470 3620 8490 3780
rect 8630 3620 8650 3780
rect 8470 3600 8650 3620
rect 9920 3780 10100 3800
rect 9920 3620 9940 3780
rect 10080 3620 10100 3780
rect 9920 3600 10100 3620
rect 11370 3780 11550 3800
rect 11370 3620 11390 3780
rect 11530 3620 11550 3780
rect 11370 3600 11550 3620
rect 330 3580 570 3600
rect 260 3220 1380 3350
rect 1460 3220 8390 3350
rect 260 -6670 460 3220
rect 11230 -6670 11430 -6664
rect 260 -6870 11230 -6670
rect 11230 -6876 11430 -6870
rect 11230 -7070 11430 -7064
rect 10430 -7090 11050 -7070
rect 10430 -7250 10450 -7090
rect 11030 -7250 11050 -7090
rect 10430 -7270 11050 -7250
rect 11221 -7270 11230 -7070
rect 11430 -7270 11439 -7070
rect 11230 -7276 11430 -7270
rect 8970 -7490 9590 -7470
rect 8970 -7650 8990 -7490
rect 9570 -7650 9590 -7490
rect 8970 -7670 9590 -7650
<< via2 >>
rect 350 4000 550 4200
rect 860 4020 1120 4180
rect 8990 4020 9570 4180
rect 10450 4020 11030 4180
rect 350 3600 550 3800
rect 1560 3620 1710 3780
rect 8490 3620 8630 3780
rect 9940 3620 10080 3780
rect 11390 3620 11530 3780
rect 10450 -7250 11030 -7090
rect 11230 -7270 11430 -7070
rect 8990 -7650 9570 -7490
rect 11230 -7670 11430 -7470
<< metal3 >>
rect 330 4205 570 4220
rect 330 3995 345 4205
rect 555 3995 570 4205
rect 840 4180 1140 4200
rect 840 4020 860 4180
rect 1120 4020 1140 4180
rect 840 4000 1140 4020
rect 8970 4180 9590 4200
rect 8970 4020 8990 4180
rect 9570 4020 9590 4180
rect 8970 4000 9590 4020
rect 10430 4180 11050 4200
rect 10430 4020 10450 4180
rect 11030 4020 11050 4180
rect 10430 4000 11050 4020
rect 330 3980 570 3995
rect 345 3800 555 3805
rect 345 3600 350 3800
rect 550 3780 11550 3800
rect 550 3620 1560 3780
rect 1710 3620 8490 3780
rect 8630 3620 9940 3780
rect 10080 3620 11390 3780
rect 11530 3620 11550 3780
rect 550 3600 11550 3620
rect 345 3595 555 3600
rect 11225 -7070 11435 -7065
rect 260 -7090 11230 -7070
rect 260 -7250 10450 -7090
rect 11030 -7250 11230 -7090
rect 260 -7270 11230 -7250
rect 11430 -7270 11435 -7070
rect 11225 -7275 11435 -7270
rect 8970 -7490 9590 -7470
rect 8970 -7650 8990 -7490
rect 9570 -7650 9590 -7490
rect 8970 -7670 9590 -7650
rect 11219 -7675 11225 -7465
rect 11425 -7470 11435 -7465
rect 11430 -7670 11435 -7470
rect 11425 -7675 11435 -7670
<< via3 >>
rect 345 4200 555 4205
rect 345 4000 350 4200
rect 350 4000 550 4200
rect 550 4000 555 4200
rect 345 3995 555 4000
rect 860 4020 1120 4180
rect 8990 4020 9570 4180
rect 10450 4020 11030 4180
rect 8990 -7650 9570 -7490
rect 11225 -7470 11425 -7465
rect 11225 -7670 11230 -7470
rect 11230 -7670 11425 -7470
rect 11225 -7675 11425 -7670
<< metal4 >>
rect 344 4205 556 4206
rect 344 3995 345 4205
rect 555 4200 556 4205
rect 555 4180 11550 4200
rect 555 4020 860 4180
rect 1120 4020 8990 4180
rect 9570 4020 10450 4180
rect 11030 4020 11550 4180
rect 555 4000 11550 4020
rect 555 3995 556 4000
rect 344 3994 556 3995
rect 11224 -7465 11426 -7464
rect 11224 -7470 11225 -7465
rect 260 -7490 11225 -7470
rect 260 -7650 8990 -7490
rect 9570 -7650 11225 -7490
rect 260 -7670 11225 -7650
rect 11224 -7675 11225 -7670
rect 11425 -7675 11426 -7465
rect 11224 -7676 11426 -7675
use sky130_fd_pr__nfet_01v8_HZS9GD  XMB0 csdac_nom__devices
timestamp 1723498766
transform 1 0 2778 0 1 -8278
box -1796 -260 1796 260
use sky130_fd_pr__nfet_01v8_FMHZDY  XMB1 csdac_nom__devices
timestamp 1723498766
transform 1 0 6436 0 1 -9110
box -996 -260 996 260
use sky130_fd_pr__nfet_01v8_AHZR5K  XMB2 csdac_nom__devices
timestamp 1723498766
transform 1 0 8713 0 1 -9269
box -596 -260 596 260
use sky130_fd_pr__nfet_01v8_BHEWB6  XMB3 csdac_nom__devices
timestamp 1723498766
transform 1 0 10400 0 1 -9428
box -406 -260 406 260
use sky130_fd_pr__nfet_01v8_FMMQLY  XMB4 csdac_nom__devices
timestamp 1723498766
transform 1 0 11787 0 1 -9587
box -296 -260 296 260
use sky130_fd_pr__nfet_01v8_C4RU6Y  XMB5 csdac_nom__devices
timestamp 1723498766
transform 1 0 13194 0 1 -9606
box -426 -400 426 400
use sky130_fd_pr__nfet_01v8_N5FCK4  XMB6 csdac_nom__devices
timestamp 1723498766
transform 1 0 14551 0 1 -9845
box -246 -320 246 320
use sky130_fd_pr__nfet_01v8_8TEC39  XMB7 csdac_nom__devices
timestamp 1723498766
transform 1 0 15728 0 1 -9904
box -246 -420 246 420
use sky130_fd_pr__nfet_01v8_SMGLWN  XMmirror csdac_nom__devices
timestamp 1723498766
transform 1 0 1505 0 1 4867
box -246 -260 246 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMN0 csdac_nom__devices
timestamp 1723498766
transform 1 0 5282 0 1 -9057
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMN1
timestamp 1723498766
transform 1 0 7959 0 1 -9216
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMN2
timestamp 1723498766
transform 1 0 9836 0 1 -9375
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMN3
timestamp 1723498766
transform 1 0 11333 0 1 -9534
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMN4
timestamp 1723498766
transform 1 0 12610 0 1 -9693
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_648S5X  XMN5 csdac_nom__devices
timestamp 1723498766
transform 1 0 14147 0 1 -9802
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_ATLS57  XMN6 csdac_nom__devices
timestamp 1723498766
transform 1 0 15324 0 1 -9861
box -211 -410 211 410
use sky130_fd_pr__nfet_01v8_J2SMEF  XMN7 csdac_nom__devices
timestamp 1723498766
transform 1 0 16501 0 1 -9920
box -211 -510 211 510
use sky130_fd_pr__nfet_01v8_L9ESAD  XMP0
timestamp 1723498766
transform 1 0 4913 0 1 -9004
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMP1
timestamp 1723498766
transform 1 0 7590 0 1 -9163
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMP2
timestamp 1723498766
transform 1 0 9467 0 1 -9322
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMP3
timestamp 1723498766
transform 1 0 10964 0 1 -9481
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMP4
timestamp 1723498766
transform 1 0 12241 0 1 -9640
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_648S5X  XMP5
timestamp 1723498766
transform 1 0 13778 0 1 -9749
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_ATLS57  XMP6
timestamp 1723498766
transform 1 0 14955 0 1 -9808
box -211 -410 211 410
use sky130_fd_pr__nfet_01v8_J2SMEF  XMP7
timestamp 1723498766
transform 1 0 16132 0 1 -9867
box -211 -510 211 510
use sky130_fd_pr__pfet_01v8_XJ7GBL  XMprog csdac_nom__devices
timestamp 1723498766
transform 1 0 1031 0 1 4869
box -211 -269 211 269
use sky130_fd_pr__res_high_po_5p73_MRHKYZ  XR5 csdac_nom__devices
timestamp 1723498766
transform 1 0 9279 0 1 -1618
box -739 -4582 739 4582
use sky130_fd_pr__res_high_po_5p73_MRHKYZ  XR6
timestamp 1723498766
transform 1 0 10739 0 1 -1618
box -739 -4582 739 4582
<< labels >>
flabel metal1 7994 5696 8194 5896 0 FreeSans 256 90 0 0 p0
port 2 nsew
flabel metal1 7594 5696 7794 5896 0 FreeSans 256 90 0 0 n0
port 3 nsew
flabel metal1 7194 5696 7394 5896 0 FreeSans 256 90 0 0 p1
port 4 nsew
flabel metal1 6794 5696 6994 5896 0 FreeSans 256 90 0 0 n1
port 5 nsew
flabel metal1 6394 5696 6594 5896 0 FreeSans 256 90 0 0 p2
port 6 nsew
flabel metal1 5994 5696 6194 5896 0 FreeSans 256 90 0 0 n2
port 7 nsew
flabel metal1 5594 5696 5794 5896 0 FreeSans 256 90 0 0 p3
port 8 nsew
flabel metal1 5194 5696 5394 5896 0 FreeSans 256 90 0 0 n3
port 9 nsew
flabel metal1 4794 5696 4994 5896 0 FreeSans 256 90 0 0 p4
port 10 nsew
flabel metal1 4394 5696 4594 5896 0 FreeSans 256 90 0 0 n4
port 11 nsew
flabel metal1 3994 5696 4194 5896 0 FreeSans 256 90 0 0 p5
port 12 nsew
flabel metal1 3594 5696 3794 5896 0 FreeSans 256 90 0 0 n5
port 13 nsew
flabel metal1 3194 5696 3394 5896 0 FreeSans 256 90 0 0 p6
port 14 nsew
flabel metal1 2794 5696 2994 5896 0 FreeSans 256 90 0 0 n6
port 15 nsew
flabel metal1 2394 5696 2594 5896 0 FreeSans 256 90 0 0 p7
port 16 nsew
flabel metal1 1994 5696 2194 5896 0 FreeSans 256 90 0 0 n7
port 17 nsew
flabel metal1 0 4000 200 4200 0 FreeSans 256 0 0 0 vcc
port 0 nsew
flabel metal1 0 3600 200 3800 0 FreeSans 256 0 0 0 vss
port 1 nsew
flabel metal1 11510 -7670 11710 -7470 0 FreeSans 256 180 0 0 Vpos
port 18 nsew
flabel metal1 11510 -6870 11710 -6670 0 FreeSans 256 180 0 0 Vbias
port 20 nsew
flabel metal1 11510 -7270 11710 -7070 0 FreeSans 256 180 0 0 Vneg
port 19 nsew
<< end >>

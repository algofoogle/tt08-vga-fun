magic
tech sky130A
magscale 1 2
timestamp 1725609024
<< pwell >>
rect 1880 -1960 1930 -1760
<< viali >>
rect 930 -1140 1700 -1010
rect 830 -2310 870 -1650
rect 1640 -2060 1690 -1790
rect 1040 -2320 1190 -2260
rect 830 -2850 870 -2490
rect 1560 -2850 1600 -2490
rect 1550 -3240 1700 -3140
rect 1150 -3530 1280 -3280
rect 1140 -4250 1200 -4060
<< metal1 >>
rect 750 -610 810 -604
rect 730 -670 750 -610
rect 810 -660 1520 -610
rect 810 -670 980 -660
rect 750 -676 810 -670
rect 920 -900 980 -670
rect 1020 -760 1420 -750
rect 1020 -820 1030 -760
rect 1410 -820 1420 -760
rect 1020 -830 1420 -820
rect 1460 -900 1520 -660
rect 1790 -780 1870 -770
rect 1790 -840 1800 -780
rect 1860 -840 1870 -780
rect 1020 -1000 1420 -920
rect 800 -1010 1780 -1000
rect 800 -1140 860 -1010
rect 1700 -1140 1780 -1010
rect 800 -1150 1780 -1140
rect 1020 -1230 1420 -1150
rect 920 -1450 980 -1250
rect 1020 -1330 1420 -1320
rect 1020 -1390 1030 -1330
rect 1410 -1390 1420 -1330
rect 1020 -1400 1420 -1390
rect 1460 -1443 1520 -1250
rect 1880 -1280 1950 -880
rect 1790 -1370 1800 -1310
rect 1860 -1370 1870 -1310
rect 1790 -1380 1870 -1370
rect 1414 -1449 1520 -1443
rect 920 -1500 1414 -1450
rect 1466 -1500 1520 -1449
rect 1414 -1507 1466 -1501
rect 1020 -1540 1200 -1530
rect 1800 -1540 1860 -1380
rect 1020 -1600 1030 -1540
rect 1190 -1600 1860 -1540
rect 1020 -1620 1860 -1600
rect 800 -1650 880 -1630
rect 800 -2310 830 -1650
rect 870 -2250 880 -1650
rect 1020 -1670 1200 -1620
rect 910 -1690 980 -1680
rect 910 -1750 920 -1690
rect 910 -1760 980 -1750
rect 1240 -1690 1310 -1680
rect 1300 -1750 1310 -1690
rect 1800 -1720 1860 -1620
rect 1240 -1760 1310 -1750
rect 1910 -1760 1950 -1280
rect 910 -2080 980 -2070
rect 1020 -2080 1200 -1770
rect 1620 -1790 1800 -1770
rect 1620 -2060 1640 -1790
rect 1690 -1950 1800 -1790
rect 1690 -2060 1710 -1950
rect 1880 -1960 1950 -1760
rect 1780 -2050 1790 -1990
rect 1870 -2050 1880 -1990
rect 1780 -2060 1880 -2050
rect 1240 -2080 1310 -2070
rect 910 -2160 920 -2080
rect 910 -2170 980 -2160
rect 1300 -2160 1310 -2080
rect 1240 -2170 1310 -2160
rect 1020 -2250 1200 -2170
rect 870 -2260 1220 -2250
rect 1620 -2260 1710 -2060
rect 870 -2310 1040 -2260
rect 800 -2320 1040 -2310
rect 1190 -2270 1220 -2260
rect 1500 -2270 1710 -2260
rect 1190 -2320 1510 -2270
rect 800 -2340 1510 -2320
rect 800 -2490 880 -2340
rect 1500 -2350 1510 -2340
rect 1620 -2340 1710 -2270
rect 1620 -2350 1630 -2340
rect 1500 -2360 1630 -2350
rect 800 -2850 830 -2490
rect 870 -2580 880 -2490
rect 970 -2480 1050 -2460
rect 970 -2540 980 -2480
rect 1040 -2540 1050 -2480
rect 1380 -2480 1460 -2460
rect 1380 -2540 1390 -2480
rect 1450 -2540 1460 -2480
rect 1550 -2490 1630 -2360
rect 1550 -2580 1560 -2490
rect 870 -2760 980 -2580
rect 1060 -2760 1370 -2580
rect 1450 -2760 1560 -2580
rect 870 -2850 880 -2760
rect 800 -2870 880 -2850
rect 970 -2860 980 -2800
rect 1040 -2860 1050 -2800
rect 970 -2880 1050 -2860
rect 1240 -2975 1290 -2760
rect 1380 -2860 1390 -2800
rect 1450 -2860 1460 -2800
rect 1380 -2880 1460 -2860
rect 1550 -2850 1560 -2760
rect 1600 -2850 1630 -2490
rect 1550 -2870 1630 -2850
rect 1910 -2902 1950 -1960
rect 1910 -2942 2030 -2902
rect 1240 -3025 1945 -2975
rect 1240 -3030 1290 -3025
rect 960 -3130 1060 -3110
rect 960 -3190 980 -3130
rect 1040 -3190 1060 -3130
rect 1360 -3120 1480 -3110
rect 1770 -3120 1860 -3110
rect 1360 -3190 1380 -3120
rect 1460 -3190 1480 -3120
rect 1360 -3200 1480 -3190
rect 1530 -3130 1720 -3120
rect 1530 -3250 1540 -3130
rect 1710 -3250 1720 -3130
rect 1770 -3180 1780 -3120
rect 1850 -3180 1860 -3120
rect 1770 -3190 1860 -3180
rect 1530 -3260 1720 -3250
rect 1050 -3280 1370 -3260
rect 1050 -3400 1150 -3280
rect 880 -3560 980 -3440
rect 1130 -3530 1150 -3400
rect 1280 -3400 1370 -3280
rect 1280 -3530 1300 -3400
rect 1130 -3550 1300 -3530
rect 1460 -3540 1790 -3300
rect 880 -3640 960 -3560
rect 1895 -3590 1945 -3025
rect 1895 -3620 1950 -3590
rect 1880 -3630 1950 -3620
rect 1890 -3640 1950 -3630
rect 880 -4080 920 -3640
rect 1820 -3670 1860 -3660
rect 960 -3730 980 -3670
rect 1040 -3730 1060 -3670
rect 960 -3750 1060 -3730
rect 1360 -3740 1370 -3670
rect 1470 -3740 1480 -3670
rect 1360 -3750 1480 -3740
rect 1770 -3740 1780 -3670
rect 1870 -3740 1880 -3670
rect 1770 -3750 1880 -3740
rect 1598 -3896 1604 -3844
rect 1656 -3850 1662 -3844
rect 1910 -3850 1950 -3640
rect 1656 -3890 1950 -3850
rect 1656 -3896 1662 -3890
rect 1120 -3940 1220 -3930
rect 960 -3990 1060 -3970
rect 960 -4050 980 -3990
rect 1040 -4050 1060 -3990
rect 1120 -4040 1130 -3940
rect 1210 -4040 1220 -3940
rect 1990 -4040 2030 -2942
rect 1120 -4060 1220 -4040
rect 1120 -4080 1140 -4060
rect 880 -4160 960 -4080
rect 860 -4240 960 -4160
rect 860 -4480 910 -4240
rect 1060 -4250 1140 -4080
rect 1200 -4250 1220 -4060
rect 1060 -4270 1220 -4250
rect 1960 -4080 2030 -4040
rect 960 -4370 980 -4310
rect 1040 -4370 1060 -4310
rect 960 -4390 1060 -4370
rect 1960 -4478 2000 -4080
rect 860 -4490 950 -4480
rect 860 -4560 870 -4490
rect 940 -4560 950 -4490
rect 1954 -4484 2006 -4478
rect 1954 -4542 2006 -4536
rect 860 -4570 950 -4560
<< via1 >>
rect 750 -670 810 -610
rect 1030 -820 1410 -760
rect 1800 -840 1860 -780
rect 860 -1140 930 -1010
rect 930 -1140 970 -1010
rect 1030 -1390 1410 -1330
rect 1800 -1370 1860 -1310
rect 1414 -1501 1466 -1449
rect 1030 -1600 1190 -1540
rect 920 -1750 980 -1690
rect 1240 -1750 1300 -1690
rect 1790 -2050 1870 -1990
rect 920 -2160 980 -2080
rect 1240 -2160 1300 -2080
rect 1510 -2350 1620 -2270
rect 980 -2540 1040 -2480
rect 1390 -2540 1450 -2480
rect 980 -2860 1040 -2800
rect 1390 -2860 1450 -2800
rect 980 -3190 1040 -3130
rect 1380 -3190 1460 -3120
rect 1540 -3140 1710 -3130
rect 1540 -3240 1550 -3140
rect 1550 -3240 1700 -3140
rect 1700 -3240 1710 -3140
rect 1540 -3250 1710 -3240
rect 1780 -3180 1850 -3120
rect 1160 -3530 1270 -3280
rect 980 -3730 1040 -3670
rect 1370 -3740 1470 -3670
rect 1780 -3740 1870 -3670
rect 1604 -3896 1656 -3844
rect 980 -4050 1040 -3990
rect 1130 -4040 1210 -3940
rect 980 -4370 1040 -4310
rect 870 -4560 940 -4490
rect 1954 -4536 2006 -4484
<< metal2 >>
rect 720 -330 840 -210
rect 1510 -330 1630 -210
rect 750 -610 810 -330
rect 744 -670 750 -610
rect 810 -670 816 -610
rect 750 -1530 810 -670
rect 1020 -760 1420 -750
rect 1020 -820 1030 -760
rect 1410 -820 1420 -760
rect 850 -1010 980 -1000
rect 850 -1140 860 -1010
rect 970 -1140 980 -1010
rect 850 -1150 980 -1140
rect 1020 -1330 1420 -820
rect 1020 -1390 1030 -1330
rect 1410 -1390 1420 -1330
rect 1020 -1400 1420 -1390
rect 750 -1590 980 -1530
rect 750 -2380 810 -1590
rect 920 -1690 980 -1590
rect 1020 -1540 1200 -1400
rect 1408 -1501 1414 -1449
rect 1466 -1501 1472 -1449
rect 1545 -1501 1595 -330
rect 1020 -1600 1030 -1540
rect 1190 -1600 1200 -1540
rect 1020 -1610 1200 -1600
rect 1415 -1551 1595 -1501
rect 920 -1800 980 -1750
rect 1240 -1690 1300 -1670
rect 1240 -1800 1300 -1750
rect 920 -1860 1300 -1800
rect 1415 -1945 1465 -1551
rect 1245 -1995 1465 -1945
rect 1245 -2070 1295 -1995
rect 910 -2080 980 -2070
rect 910 -2160 920 -2080
rect 910 -2170 980 -2160
rect 1240 -2080 1310 -2070
rect 1300 -2160 1310 -2080
rect 1240 -2170 1310 -2160
rect 925 -2215 975 -2170
rect 1245 -2215 1295 -2170
rect 1545 -2175 1595 -1551
rect 1670 -780 1880 -770
rect 1670 -840 1800 -780
rect 1860 -840 1880 -780
rect 1670 -1300 1740 -840
rect 1670 -1310 1880 -1300
rect 1670 -1370 1800 -1310
rect 1860 -1370 1880 -1310
rect 1670 -1985 1740 -1370
rect 1780 -1985 1880 -1980
rect 1670 -1990 1880 -1985
rect 1670 -2050 1790 -1990
rect 1870 -2050 1880 -1990
rect 1670 -2055 1880 -2050
rect 1780 -2060 1880 -2055
rect 925 -2265 1295 -2215
rect 1395 -2225 1595 -2175
rect 750 -2440 1040 -2380
rect 980 -2470 1040 -2440
rect 1395 -2470 1445 -2225
rect 1500 -2270 1630 -2260
rect 1500 -2350 1510 -2270
rect 1620 -2350 1630 -2270
rect 1500 -2360 1630 -2350
rect 970 -2480 1050 -2470
rect 970 -2540 980 -2480
rect 1040 -2540 1050 -2480
rect 970 -2550 1050 -2540
rect 1380 -2480 1460 -2470
rect 1380 -2540 1390 -2480
rect 1450 -2540 1460 -2480
rect 1380 -2550 1460 -2540
rect 980 -2790 1040 -2550
rect 1395 -2790 1445 -2550
rect 970 -2800 1050 -2790
rect 970 -2860 980 -2800
rect 1040 -2860 1050 -2800
rect 970 -2940 1050 -2860
rect 1380 -2800 1460 -2790
rect 1380 -2860 1390 -2800
rect 1450 -2860 1460 -2800
rect 1380 -2940 1460 -2860
rect 1600 -2940 1710 -2930
rect 970 -3020 1230 -2940
rect 1380 -2950 1870 -2940
rect 1380 -3020 1620 -2950
rect 1690 -3020 1870 -2950
rect 960 -3130 1060 -3110
rect 960 -3190 980 -3130
rect 1040 -3190 1060 -3130
rect 960 -3670 1060 -3190
rect 1150 -3120 1230 -3020
rect 1600 -3040 1710 -3020
rect 1790 -3110 1870 -3020
rect 1360 -3120 1480 -3110
rect 1770 -3120 1890 -3110
rect 1150 -3190 1380 -3120
rect 1460 -3190 1480 -3120
rect 1150 -3200 1480 -3190
rect 1530 -3130 1720 -3120
rect 1140 -3280 1290 -3260
rect 1140 -3530 1160 -3280
rect 1270 -3530 1290 -3280
rect 1140 -3550 1290 -3530
rect 1380 -3660 1460 -3200
rect 1530 -3250 1540 -3130
rect 1710 -3250 1720 -3130
rect 1770 -3180 1780 -3120
rect 1850 -3180 1890 -3120
rect 1770 -3200 1890 -3180
rect 1530 -3260 1720 -3250
rect 1790 -3660 1870 -3200
rect 960 -3730 980 -3670
rect 1040 -3730 1060 -3670
rect 960 -3850 1060 -3730
rect 1360 -3670 1480 -3660
rect 1360 -3740 1370 -3670
rect 1470 -3740 1480 -3670
rect 1360 -3750 1480 -3740
rect 1770 -3670 1890 -3660
rect 1770 -3740 1780 -3670
rect 1870 -3740 1890 -3670
rect 1770 -3750 1890 -3740
rect 1604 -3844 1656 -3838
rect 960 -3890 1604 -3850
rect 960 -3990 1060 -3890
rect 1604 -3902 1656 -3896
rect 960 -4050 980 -3990
rect 1040 -4050 1060 -3990
rect 1120 -3940 1220 -3930
rect 1120 -4040 1130 -3940
rect 1210 -4040 1220 -3940
rect 1120 -4050 1220 -4040
rect 960 -4310 1060 -4050
rect 960 -4370 980 -4310
rect 1040 -4370 1060 -4310
rect 960 -4390 1060 -4370
rect 860 -4560 870 -4490
rect 940 -4560 980 -4490
rect 860 -4700 980 -4560
rect 1381 -4570 1390 -4450
rect 1510 -4570 1519 -4450
rect 1948 -4536 1954 -4484
rect 2006 -4536 2012 -4484
rect 1390 -4700 1510 -4570
rect 1960 -4580 2000 -4536
rect 1920 -4700 2040 -4580
<< via2 >>
rect 860 -1140 970 -1010
rect 1510 -2350 1620 -2270
rect 1620 -3020 1690 -2950
rect 1160 -3530 1270 -3280
rect 1540 -3250 1710 -3130
rect 1130 -4040 1210 -3940
rect 1390 -4570 1510 -4450
<< metal3 >>
rect 950 -400 1070 -210
rect 850 -540 1070 -400
rect 1240 -415 1360 -210
rect 1240 -540 1385 -415
rect 850 -1010 980 -540
rect 850 -1140 860 -1010
rect 970 -1140 980 -1010
rect 850 -3725 980 -1140
rect 1255 -1545 1385 -540
rect 1255 -1675 1630 -1545
rect 1500 -2140 1630 -1675
rect 1500 -2270 1905 -2140
rect 1500 -2350 1510 -2270
rect 1620 -2350 1630 -2270
rect 1500 -2360 1630 -2350
rect 1775 -2920 1905 -2270
rect 1600 -2950 1710 -2930
rect 1600 -3020 1620 -2950
rect 1690 -3020 1710 -2950
rect 1600 -3040 1710 -3020
rect 1530 -3125 1720 -3120
rect 1415 -3130 1720 -3125
rect 1415 -3250 1540 -3130
rect 1710 -3250 1720 -3130
rect 1415 -3260 1720 -3250
rect 1140 -3280 1290 -3260
rect 1140 -3530 1160 -3280
rect 1270 -3530 1290 -3280
rect 1140 -3725 1290 -3530
rect 1415 -3725 1545 -3260
rect 1780 -3340 1905 -2920
rect 850 -3855 1545 -3725
rect 1775 -3925 1905 -3340
rect 1115 -3940 1905 -3925
rect 1115 -4040 1130 -3940
rect 1210 -4040 1905 -3940
rect 1115 -4055 1905 -4040
rect 1385 -4450 1515 -4445
rect 1385 -4570 1390 -4450
rect 1510 -4570 1590 -4450
rect 1710 -4570 1716 -4450
rect 1385 -4575 1515 -4570
<< via3 >>
rect 1620 -3020 1690 -2950
rect 1590 -4570 1710 -4450
<< metal4 >>
rect 1600 -2950 1710 -2930
rect 1600 -3020 1620 -2950
rect 1690 -3020 1710 -2950
rect 1600 -4120 1710 -3020
rect 1590 -4390 1710 -4360
rect 1550 -4450 1750 -4390
rect 1550 -4560 1590 -4450
rect 1589 -4570 1590 -4560
rect 1710 -4560 1750 -4450
rect 1710 -4570 1711 -4560
rect 1589 -4571 1711 -4570
use sky130_fd_pr__res_generic_m4_VRQADB  R1
timestamp 1725602025
transform 1 0 1650 0 1 -4243
box -100 -157 100 157
use sky130_fd_pr__pfet_01v8_XLV5ZZ  XMA1
timestamp 1725602025
transform 0 1 1219 -1 0 -869
box -211 -419 211 419
use sky130_fd_pr__pfet_01v8_XLV5ZZ  XMA2
timestamp 1725602025
transform 0 1 1219 -1 0 -1279
box -211 -419 211 419
use sky130_fd_pr__nfet_01v8_V8CAV6  XMA3
timestamp 1725602025
transform 0 1 1110 -1 0 -1719
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_V8CAV6  XMA4
timestamp 1725602025
transform 0 1 1110 -1 0 -2129
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XLV5ZZ  XMA5
timestamp 1725602025
transform 1 0 1831 0 1 -1071
box -211 -419 211 419
use sky130_fd_pr__nfet_01v8_V8CAV6  XMA6
timestamp 1725602025
transform 1 0 1831 0 1 -1860
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XLV5ZZ  XMO1
timestamp 1725602025
transform -1 0 1421 0 -1 -3431
box -211 -419 211 419
use sky130_fd_pr__pfet_01v8_XLV5ZZ  XMO2
timestamp 1725602025
transform 1 0 1831 0 1 -3431
box -211 -419 211 419
use sky130_fd_pr__nfet_01v8_V8CAV6  XMO3
timestamp 1725602025
transform 1 0 1011 0 1 -2670
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_V8CAV6  XMO4
timestamp 1725602025
transform 1 0 1421 0 1 -2670
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XLV5ZZ  XMO5
timestamp 1725602025
transform 1 0 1011 0 1 -3431
box -211 -419 211 419
use sky130_fd_pr__nfet_01v8_V8CAV6  XMO6
timestamp 1725602025
transform 1 0 1011 0 1 -4180
box -211 -310 211 310
<< labels >>
flabel metal2 720 -330 840 -210 0 FreeSans 640 0 0 0 b0
port 7 nsew
flabel metal2 1510 -330 1630 -210 0 FreeSans 640 0 0 0 b1
port 8 nsew
flabel metal3 950 -330 1070 -210 0 FreeSans 640 0 0 0 VCC
port 10 nsew
flabel metal3 1240 -330 1360 -210 0 FreeSans 640 0 0 0 VSS
port 11 nsew
flabel metal2 860 -4700 980 -4580 0 FreeSans 640 0 0 0 s1
port 12 nsew
flabel metal2 1920 -4700 2040 -4580 0 FreeSans 640 0 0 0 s3
port 9 nsew
flabel metal2 1390 -4700 1510 -4580 0 FreeSans 640 0 0 0 s2
port 13 nsew
<< end >>

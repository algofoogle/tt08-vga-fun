magic
tech sky130A
magscale 1 2
timestamp 1724297220
<< metal1 >>
rect 11648 15062 11654 15118
rect 11710 15062 11716 15118
rect 12016 15062 12022 15118
rect 12078 15062 12084 15118
rect 12384 15062 12390 15118
rect 12446 15062 12452 15118
rect 12752 15062 12758 15118
rect 12814 15062 12820 15118
rect 13120 15062 13126 15118
rect 13182 15062 13188 15118
rect 13488 15062 13494 15118
rect 13550 15062 13556 15118
rect 13856 15062 13862 15118
rect 13918 15062 13924 15118
rect 14224 15062 14230 15118
rect 14286 15062 14292 15118
rect 14592 15062 14598 15118
rect 14654 15062 14660 15118
rect 14960 15062 14966 15118
rect 15022 15062 15028 15118
rect 15328 15062 15334 15118
rect 15390 15062 15396 15118
rect 15696 15062 15702 15118
rect 15758 15062 15764 15118
rect 16064 15062 16070 15118
rect 16126 15062 16132 15118
rect 16432 15062 16438 15118
rect 16494 15062 16500 15118
rect 16800 15062 16806 15118
rect 16862 15062 16868 15118
rect 17168 15062 17174 15118
rect 17230 15062 17236 15118
<< via1 >>
rect 20494 18672 20550 18728
rect 20862 18672 20918 18728
rect 21230 18672 21286 18728
rect 21598 18672 21654 18728
rect 21966 18672 22022 18728
rect 22334 18672 22390 18728
rect 22702 18672 22758 18728
rect 23070 18672 23126 18728
rect 23438 18672 23494 18728
rect 23806 18672 23862 18728
rect 24174 18672 24230 18728
rect 24542 18672 24598 18728
rect 24910 18672 24966 18728
rect 25278 18672 25334 18728
rect 25646 18672 25702 18728
rect 26014 18672 26070 18728
rect 11654 15062 11710 15118
rect 12022 15062 12078 15118
rect 12390 15062 12446 15118
rect 12758 15062 12814 15118
rect 13126 15062 13182 15118
rect 13494 15062 13550 15118
rect 13862 15062 13918 15118
rect 14230 15062 14286 15118
rect 14598 15062 14654 15118
rect 14966 15062 15022 15118
rect 15334 15062 15390 15118
rect 15702 15062 15758 15118
rect 16070 15062 16126 15118
rect 16438 15062 16494 15118
rect 16806 15062 16862 15118
rect 17174 15062 17230 15118
<< metal2 >>
rect 10704 44870 10824 44900
rect 10704 44810 10732 44870
rect 10792 44810 10824 44870
rect 10704 44780 10824 44810
rect 11256 44870 11376 44900
rect 11256 44810 11284 44870
rect 11344 44810 11376 44870
rect 11256 44780 11376 44810
rect 11808 44870 11928 44900
rect 11808 44810 11836 44870
rect 11896 44810 11928 44870
rect 11808 44780 11928 44810
rect 12360 44870 12480 44900
rect 12360 44810 12388 44870
rect 12448 44810 12480 44870
rect 12360 44780 12480 44810
rect 12912 44870 13032 44900
rect 12912 44810 12940 44870
rect 13000 44810 13032 44870
rect 12912 44780 13032 44810
rect 13464 44870 13584 44900
rect 13464 44810 13492 44870
rect 13552 44810 13584 44870
rect 13464 44780 13584 44810
rect 14016 44870 14136 44900
rect 14016 44810 14044 44870
rect 14104 44810 14136 44870
rect 14016 44780 14136 44810
rect 14568 44870 14688 44900
rect 14568 44810 14596 44870
rect 14656 44810 14688 44870
rect 14568 44780 14688 44810
rect 15120 44870 15240 44900
rect 15120 44810 15148 44870
rect 15208 44810 15240 44870
rect 15120 44780 15240 44810
rect 15672 44870 15792 44900
rect 15672 44810 15700 44870
rect 15760 44810 15792 44870
rect 15672 44780 15792 44810
rect 20640 44870 20760 44900
rect 20640 44810 20668 44870
rect 20728 44810 20760 44870
rect 20640 44780 20760 44810
rect 21192 44870 21312 44900
rect 21192 44810 21220 44870
rect 21280 44810 21312 44870
rect 21192 44780 21312 44810
rect 21744 44870 21864 44900
rect 21744 44810 21772 44870
rect 21832 44810 21864 44870
rect 21744 44780 21864 44810
rect 22296 44870 22416 44900
rect 22296 44810 22324 44870
rect 22384 44810 22416 44870
rect 22296 44780 22416 44810
rect 22848 44870 22968 44900
rect 22848 44810 22876 44870
rect 22936 44810 22968 44870
rect 22848 44780 22968 44810
rect 23400 44870 23520 44900
rect 23400 44810 23428 44870
rect 23488 44810 23520 44870
rect 23400 44780 23520 44810
rect 23952 44870 24072 44900
rect 23952 44810 23980 44870
rect 24040 44810 24072 44870
rect 23952 44780 24072 44810
rect 24504 44870 24624 44900
rect 24504 44810 24532 44870
rect 24592 44810 24624 44870
rect 24504 44780 24624 44810
rect 25056 44870 25176 44900
rect 25056 44810 25084 44870
rect 25144 44810 25176 44870
rect 25056 44780 25176 44810
rect 25608 44870 25728 44900
rect 25608 44810 25636 44870
rect 25696 44810 25728 44870
rect 25608 44780 25728 44810
rect 10734 44162 10790 44780
rect 11286 44162 11342 44780
rect 11838 44162 11894 44780
rect 12390 44162 12446 44780
rect 12942 44162 12998 44780
rect 13494 44162 13550 44780
rect 14046 44162 14102 44780
rect 14598 44162 14654 44780
rect 15150 44162 15206 44780
rect 15702 44162 15758 44780
rect 20670 44162 20726 44780
rect 21222 44162 21278 44780
rect 21774 44162 21830 44780
rect 22326 44162 22382 44780
rect 22878 44162 22934 44780
rect 23430 44162 23486 44780
rect 23982 44162 24038 44780
rect 24534 44162 24590 44780
rect 25086 44162 25142 44780
rect 25638 44162 25694 44780
rect 11654 15118 11710 20448
rect 11654 15056 11710 15062
rect 12022 15118 12078 20448
rect 12022 15056 12078 15062
rect 12390 15118 12446 20448
rect 12390 15056 12446 15062
rect 12758 15118 12814 20448
rect 12758 15056 12814 15062
rect 13126 15118 13182 20448
rect 13126 15056 13182 15062
rect 13494 15118 13550 20448
rect 13494 15056 13550 15062
rect 13862 15118 13918 20448
rect 13862 15056 13918 15062
rect 14230 15118 14286 20448
rect 14230 15056 14286 15062
rect 14598 15118 14654 20448
rect 14598 15056 14654 15062
rect 14966 15118 15022 20448
rect 14966 15056 15022 15062
rect 15334 15118 15390 20448
rect 15334 15056 15390 15062
rect 15702 15118 15758 20448
rect 15702 15056 15758 15062
rect 16070 15118 16126 20448
rect 16070 15056 16126 15062
rect 16438 15118 16494 20448
rect 16438 15056 16494 15062
rect 16806 15118 16862 20448
rect 16806 15056 16862 15062
rect 17174 15118 17230 20448
rect 20494 18728 20550 20580
rect 20494 18666 20550 18672
rect 20862 18728 20918 20580
rect 20862 18666 20918 18672
rect 21230 18728 21286 20580
rect 21230 18666 21286 18672
rect 21598 18728 21654 20580
rect 21598 18666 21654 18672
rect 21966 18728 22022 20580
rect 21966 18666 22022 18672
rect 22334 18728 22390 20580
rect 22334 18666 22390 18672
rect 22702 18728 22758 20580
rect 22702 18666 22758 18672
rect 23070 18728 23126 20580
rect 23070 18666 23126 18672
rect 23438 18728 23494 20580
rect 23438 18666 23494 18672
rect 23806 18728 23862 20580
rect 23806 18666 23862 18672
rect 24174 18728 24230 20580
rect 24174 18666 24230 18672
rect 24542 18728 24598 20580
rect 24542 18666 24598 18672
rect 24910 18728 24966 20580
rect 24910 18666 24966 18672
rect 25278 18728 25334 20580
rect 25278 18666 25334 18672
rect 25646 18728 25702 20580
rect 25646 18666 25702 18672
rect 26014 18728 26070 20580
rect 26014 18666 26070 18672
rect 17174 15056 17230 15062
<< via2 >>
rect 10732 44810 10792 44870
rect 11284 44810 11344 44870
rect 11836 44810 11896 44870
rect 12388 44810 12448 44870
rect 12940 44810 13000 44870
rect 13492 44810 13552 44870
rect 14044 44810 14104 44870
rect 14596 44810 14656 44870
rect 15148 44810 15208 44870
rect 15700 44810 15760 44870
rect 20668 44810 20728 44870
rect 21220 44810 21280 44870
rect 21772 44810 21832 44870
rect 22324 44810 22384 44870
rect 22876 44810 22936 44870
rect 23428 44810 23488 44870
rect 23980 44810 24040 44870
rect 24532 44810 24592 44870
rect 25084 44810 25144 44870
rect 25636 44810 25696 44870
<< metal3 >>
rect 10704 44875 10824 44900
rect 6310 44798 6316 44862
rect 6380 44798 6386 44862
rect 6862 44798 6868 44862
rect 6932 44798 6938 44862
rect 10704 44805 10727 44875
rect 10797 44805 10824 44875
rect 926 44703 1074 44704
rect 921 44557 927 44703
rect 1073 44557 1079 44703
rect 926 44064 1074 44557
rect 6318 44408 6378 44798
rect 6870 44408 6930 44798
rect 10704 44780 10824 44805
rect 11256 44875 11376 44900
rect 11256 44805 11279 44875
rect 11349 44805 11376 44875
rect 11256 44780 11376 44805
rect 11808 44875 11928 44900
rect 11808 44805 11831 44875
rect 11901 44805 11928 44875
rect 11808 44780 11928 44805
rect 12360 44875 12480 44900
rect 12360 44805 12383 44875
rect 12453 44805 12480 44875
rect 12360 44780 12480 44805
rect 12912 44875 13032 44900
rect 12912 44805 12935 44875
rect 13005 44805 13032 44875
rect 12912 44780 13032 44805
rect 13464 44875 13584 44900
rect 13464 44805 13487 44875
rect 13557 44805 13584 44875
rect 13464 44780 13584 44805
rect 14016 44875 14136 44900
rect 14016 44805 14039 44875
rect 14109 44805 14136 44875
rect 14016 44780 14136 44805
rect 14568 44875 14688 44900
rect 14568 44805 14591 44875
rect 14661 44805 14688 44875
rect 14568 44780 14688 44805
rect 15120 44875 15240 44900
rect 15120 44805 15143 44875
rect 15213 44805 15240 44875
rect 15120 44780 15240 44805
rect 15672 44875 15792 44900
rect 15672 44805 15695 44875
rect 15765 44805 15792 44875
rect 15672 44780 15792 44805
rect 20640 44875 20760 44900
rect 20640 44805 20663 44875
rect 20733 44805 20760 44875
rect 20640 44780 20760 44805
rect 21192 44875 21312 44900
rect 21192 44805 21215 44875
rect 21285 44805 21312 44875
rect 21192 44780 21312 44805
rect 21744 44875 21864 44900
rect 21744 44805 21767 44875
rect 21837 44805 21864 44875
rect 21744 44780 21864 44805
rect 22296 44875 22416 44900
rect 22296 44805 22319 44875
rect 22389 44805 22416 44875
rect 22296 44780 22416 44805
rect 22848 44875 22968 44900
rect 22848 44805 22871 44875
rect 22941 44805 22968 44875
rect 22848 44780 22968 44805
rect 23400 44875 23520 44900
rect 23400 44805 23423 44875
rect 23493 44805 23520 44875
rect 23400 44780 23520 44805
rect 23952 44875 24072 44900
rect 23952 44805 23975 44875
rect 24045 44805 24072 44875
rect 23952 44780 24072 44805
rect 24504 44875 24624 44900
rect 24504 44805 24527 44875
rect 24597 44805 24624 44875
rect 24504 44780 24624 44805
rect 25056 44875 25176 44900
rect 25056 44805 25079 44875
rect 25149 44805 25176 44875
rect 25056 44780 25176 44805
rect 25608 44875 25728 44900
rect 25608 44805 25631 44875
rect 25701 44805 25728 44875
rect 25608 44780 25728 44805
rect 6316 44402 6380 44408
rect 6316 44332 6380 44338
rect 6868 44402 6932 44408
rect 6868 44332 6932 44338
rect 926 43910 1074 43916
rect 3789 20070 4187 20075
rect 200 20069 22190 20070
rect 200 20050 3789 20069
rect 200 19690 220 20050
rect 580 19690 3789 20050
rect 200 19671 3789 19690
rect 4187 20050 22190 20069
rect 4187 19690 9830 20050
rect 10170 19690 15810 20050
rect 16170 19690 21810 20050
rect 22170 19690 22190 20050
rect 4187 19671 22190 19690
rect 200 19670 22190 19671
rect 3789 19665 4187 19670
rect 6783 19091 6789 19489
rect 7187 19091 7193 19489
rect 9520 14189 9720 19670
rect 12783 19091 12789 19489
rect 13187 19091 13193 19489
rect 18490 17769 18690 19670
rect 18783 19091 18789 19489
rect 19187 19091 19193 19489
rect 24783 19091 24789 19489
rect 25187 19091 25193 19489
rect 18490 17571 18491 17769
rect 18689 17571 18690 17769
rect 18490 17570 18690 17571
rect 18491 17565 18689 17570
rect 9520 13991 9521 14189
rect 9719 13991 9720 14189
rect 9520 13990 9720 13991
rect 9521 13985 9719 13990
<< via3 >>
rect 6316 44798 6380 44862
rect 6868 44798 6932 44862
rect 10727 44870 10797 44875
rect 10727 44810 10732 44870
rect 10732 44810 10792 44870
rect 10792 44810 10797 44870
rect 10727 44805 10797 44810
rect 927 44557 1073 44703
rect 11279 44870 11349 44875
rect 11279 44810 11284 44870
rect 11284 44810 11344 44870
rect 11344 44810 11349 44870
rect 11279 44805 11349 44810
rect 11831 44870 11901 44875
rect 11831 44810 11836 44870
rect 11836 44810 11896 44870
rect 11896 44810 11901 44870
rect 11831 44805 11901 44810
rect 12383 44870 12453 44875
rect 12383 44810 12388 44870
rect 12388 44810 12448 44870
rect 12448 44810 12453 44870
rect 12383 44805 12453 44810
rect 12935 44870 13005 44875
rect 12935 44810 12940 44870
rect 12940 44810 13000 44870
rect 13000 44810 13005 44870
rect 12935 44805 13005 44810
rect 13487 44870 13557 44875
rect 13487 44810 13492 44870
rect 13492 44810 13552 44870
rect 13552 44810 13557 44870
rect 13487 44805 13557 44810
rect 14039 44870 14109 44875
rect 14039 44810 14044 44870
rect 14044 44810 14104 44870
rect 14104 44810 14109 44870
rect 14039 44805 14109 44810
rect 14591 44870 14661 44875
rect 14591 44810 14596 44870
rect 14596 44810 14656 44870
rect 14656 44810 14661 44870
rect 14591 44805 14661 44810
rect 15143 44870 15213 44875
rect 15143 44810 15148 44870
rect 15148 44810 15208 44870
rect 15208 44810 15213 44870
rect 15143 44805 15213 44810
rect 15695 44870 15765 44875
rect 15695 44810 15700 44870
rect 15700 44810 15760 44870
rect 15760 44810 15765 44870
rect 15695 44805 15765 44810
rect 20663 44870 20733 44875
rect 20663 44810 20668 44870
rect 20668 44810 20728 44870
rect 20728 44810 20733 44870
rect 20663 44805 20733 44810
rect 21215 44870 21285 44875
rect 21215 44810 21220 44870
rect 21220 44810 21280 44870
rect 21280 44810 21285 44870
rect 21215 44805 21285 44810
rect 21767 44870 21837 44875
rect 21767 44810 21772 44870
rect 21772 44810 21832 44870
rect 21832 44810 21837 44870
rect 21767 44805 21837 44810
rect 22319 44870 22389 44875
rect 22319 44810 22324 44870
rect 22324 44810 22384 44870
rect 22384 44810 22389 44870
rect 22319 44805 22389 44810
rect 22871 44870 22941 44875
rect 22871 44810 22876 44870
rect 22876 44810 22936 44870
rect 22936 44810 22941 44870
rect 22871 44805 22941 44810
rect 23423 44870 23493 44875
rect 23423 44810 23428 44870
rect 23428 44810 23488 44870
rect 23488 44810 23493 44870
rect 23423 44805 23493 44810
rect 23975 44870 24045 44875
rect 23975 44810 23980 44870
rect 23980 44810 24040 44870
rect 24040 44810 24045 44870
rect 23975 44805 24045 44810
rect 24527 44870 24597 44875
rect 24527 44810 24532 44870
rect 24532 44810 24592 44870
rect 24592 44810 24597 44870
rect 24527 44805 24597 44810
rect 25079 44870 25149 44875
rect 25079 44810 25084 44870
rect 25084 44810 25144 44870
rect 25144 44810 25149 44870
rect 25079 44805 25149 44810
rect 25631 44870 25701 44875
rect 25631 44810 25636 44870
rect 25636 44810 25696 44870
rect 25696 44810 25701 44870
rect 25631 44805 25701 44810
rect 6316 44338 6380 44402
rect 6868 44338 6932 44402
rect 926 43916 1074 44064
rect 220 19690 580 20050
rect 3789 19671 4187 20069
rect 9830 19690 10170 20050
rect 15810 19690 16170 20050
rect 21810 19690 22170 20050
rect 6789 19091 7187 19489
rect 12789 19091 13187 19489
rect 18789 19091 19187 19489
rect 24789 19091 25187 19489
rect 18491 17571 18689 17769
rect 9521 13991 9719 14189
<< metal4 >>
rect 926 44703 1074 44704
rect 926 44557 927 44703
rect 1073 44696 1074 44703
rect 3006 44696 3066 45152
rect 3558 44696 3618 45152
rect 4110 44696 4170 45152
rect 4662 44696 4722 45152
rect 5214 44696 5274 45152
rect 5766 44696 5826 45152
rect 6318 44863 6378 45152
rect 6870 44863 6930 45152
rect 6315 44862 6381 44863
rect 6315 44798 6316 44862
rect 6380 44798 6381 44862
rect 6315 44797 6381 44798
rect 6867 44862 6933 44863
rect 6867 44798 6868 44862
rect 6932 44798 6933 44862
rect 6867 44797 6933 44798
rect 7422 44696 7482 45152
rect 7974 44696 8034 45152
rect 8526 44696 8586 45152
rect 9078 44696 9138 45152
rect 9630 44696 9690 45152
rect 10182 44696 10242 45152
rect 10734 45010 10794 45152
rect 11286 45010 11346 45152
rect 11838 45010 11898 45152
rect 12390 45010 12450 45152
rect 12942 45010 13002 45152
rect 13494 45010 13554 45152
rect 14046 45010 14106 45152
rect 14598 45010 14658 45152
rect 15150 45010 15210 45152
rect 15702 45010 15762 45152
rect 10724 44900 10804 45010
rect 11276 44900 11356 45010
rect 11828 44900 11908 45010
rect 12380 44900 12460 45010
rect 12932 44900 13012 45010
rect 13484 44900 13564 45010
rect 14036 44900 14116 45010
rect 14588 44900 14668 45010
rect 15140 44900 15220 45010
rect 15692 44900 15772 45010
rect 16254 44952 16314 45152
rect 16806 44952 16866 45152
rect 17358 44952 17418 45152
rect 17910 44952 17970 45152
rect 18462 44952 18522 45152
rect 19014 44952 19074 45152
rect 19566 44952 19626 45152
rect 20118 44952 20178 45152
rect 20670 45010 20730 45152
rect 21222 45010 21282 45152
rect 21774 45010 21834 45152
rect 22326 45010 22386 45152
rect 22878 45010 22938 45152
rect 23430 45010 23490 45152
rect 23982 45010 24042 45152
rect 24534 45010 24594 45152
rect 25086 45010 25146 45152
rect 25638 45010 25698 45152
rect 20660 44900 20740 45010
rect 21212 44900 21292 45010
rect 21764 44900 21844 45010
rect 22316 44900 22396 45010
rect 22868 44900 22948 45010
rect 23420 44900 23500 45010
rect 23972 44900 24052 45010
rect 24524 44900 24604 45010
rect 25076 44900 25156 45010
rect 25628 44900 25708 45010
rect 26190 44952 26250 45152
rect 10704 44875 10824 44900
rect 10704 44805 10727 44875
rect 10797 44805 10824 44875
rect 10704 44780 10824 44805
rect 11256 44875 11376 44900
rect 11256 44805 11279 44875
rect 11349 44805 11376 44875
rect 11256 44780 11376 44805
rect 11808 44875 11928 44900
rect 11808 44805 11831 44875
rect 11901 44805 11928 44875
rect 11808 44780 11928 44805
rect 12360 44875 12480 44900
rect 12360 44805 12383 44875
rect 12453 44805 12480 44875
rect 12360 44780 12480 44805
rect 12912 44875 13032 44900
rect 12912 44805 12935 44875
rect 13005 44805 13032 44875
rect 12912 44780 13032 44805
rect 13464 44875 13584 44900
rect 13464 44805 13487 44875
rect 13557 44805 13584 44875
rect 13464 44780 13584 44805
rect 14016 44875 14136 44900
rect 14016 44805 14039 44875
rect 14109 44805 14136 44875
rect 14016 44780 14136 44805
rect 14568 44875 14688 44900
rect 14568 44805 14591 44875
rect 14661 44805 14688 44875
rect 14568 44780 14688 44805
rect 15120 44875 15240 44900
rect 15120 44805 15143 44875
rect 15213 44805 15240 44875
rect 15120 44780 15240 44805
rect 15672 44875 15792 44900
rect 15672 44805 15695 44875
rect 15765 44805 15792 44875
rect 15672 44780 15792 44805
rect 20640 44875 20760 44900
rect 20640 44805 20663 44875
rect 20733 44805 20760 44875
rect 20640 44780 20760 44805
rect 21192 44875 21312 44900
rect 21192 44805 21215 44875
rect 21285 44805 21312 44875
rect 21192 44780 21312 44805
rect 21744 44875 21864 44900
rect 21744 44805 21767 44875
rect 21837 44805 21864 44875
rect 21744 44780 21864 44805
rect 22296 44875 22416 44900
rect 22296 44805 22319 44875
rect 22389 44805 22416 44875
rect 22296 44780 22416 44805
rect 22848 44875 22968 44900
rect 22848 44805 22871 44875
rect 22941 44805 22968 44875
rect 22848 44780 22968 44805
rect 23400 44875 23520 44900
rect 23400 44805 23423 44875
rect 23493 44805 23520 44875
rect 23400 44780 23520 44805
rect 23952 44875 24072 44900
rect 23952 44805 23975 44875
rect 24045 44805 24072 44875
rect 23952 44780 24072 44805
rect 24504 44875 24624 44900
rect 24504 44805 24527 44875
rect 24597 44805 24624 44875
rect 24504 44780 24624 44805
rect 25056 44875 25176 44900
rect 25056 44805 25079 44875
rect 25149 44805 25176 44875
rect 25056 44780 25176 44805
rect 25608 44875 25728 44900
rect 25608 44805 25631 44875
rect 25701 44805 25728 44875
rect 25608 44780 25728 44805
rect 1073 44564 10316 44696
rect 1073 44557 1074 44564
rect 926 44556 1074 44557
rect 321 44442 479 44449
rect 321 44402 7092 44442
rect 321 44338 6316 44402
rect 6380 44338 6868 44402
rect 6932 44338 7092 44402
rect 321 44298 7092 44338
rect 321 44152 479 44298
rect 928 44152 1072 44160
rect 200 20050 600 44152
rect 200 19690 220 20050
rect 580 19690 600 20050
rect 200 1000 600 19690
rect 800 44064 1200 44152
rect 800 43916 926 44064
rect 1074 43916 1200 44064
rect 800 19490 1200 43916
rect 3788 20069 4188 21180
rect 3788 19671 3789 20069
rect 4187 19671 4188 20069
rect 3788 19670 4188 19671
rect 6788 19490 7188 21260
rect 9788 20050 10188 21180
rect 9788 19690 9830 20050
rect 10170 19690 10188 20050
rect 9788 19670 10188 19690
rect 12788 19490 13188 21260
rect 15788 20050 16188 21180
rect 15788 19690 15810 20050
rect 16170 19690 16188 20050
rect 15788 19670 16188 19690
rect 18788 19490 19188 21260
rect 21788 20050 22188 21180
rect 21788 19690 21810 20050
rect 22170 19690 22188 20050
rect 21788 19670 22188 19690
rect 24788 19490 25188 21260
rect 800 19489 25200 19490
rect 800 19091 6789 19489
rect 7187 19091 12789 19489
rect 13187 19091 18789 19489
rect 19187 19091 24789 19489
rect 25187 19091 25200 19489
rect 800 19090 25200 19091
rect 800 1000 1200 19090
rect 9140 13790 9340 19090
rect 18160 17370 18360 19090
rect 18490 17769 19280 17770
rect 18490 17571 18491 17769
rect 18689 17571 19280 17769
rect 18490 17570 19280 17571
rect 18160 17170 19320 17370
rect 9520 14189 10440 14190
rect 9520 13991 9521 14189
rect 9719 13991 10440 14189
rect 9520 13990 10440 13991
rect 9140 13590 10450 13790
rect 19186 4096 23544 4264
rect 25158 4198 27402 4362
rect 16338 618 19682 782
rect 186 0 366 200
rect 4050 0 4230 200
rect 7914 0 8094 200
rect 11778 0 11958 200
rect 15642 0 15822 220
rect 19518 200 19682 618
rect 23376 200 23544 4096
rect 27238 200 27402 4198
rect 28560 1000 28960 44152
rect 19506 0 19686 200
rect 23370 0 23550 200
rect 27234 0 27414 200
use controller  controller_0
timestamp 1724295482
transform 1 0 2436 0 1 20284
box 386 0 23630 24000
use csdac_nom  green_dac
timestamp 1724297071
transform 1 0 10230 0 1 9990
box 0 -9390 9210 5196
use csdac_nom  red_dac
timestamp 1724297071
transform 1 0 19070 0 1 13570
box 0 -9390 9210 5196
<< labels >>
flabel metal4 s 25638 44952 25698 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 26190 44952 26250 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 27234 0 27414 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 23370 0 23550 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 19506 0 19686 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 15642 0 15822 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 11778 0 11958 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 7914 0 8094 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4050 0 4230 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 186 0 366 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 24534 44952 24594 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 23982 44952 24042 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 23430 44952 23490 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 22326 44952 22386 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 21774 44952 21834 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 21222 44952 21282 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 20118 44952 20178 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 19566 44952 19626 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 19014 44952 19074 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 17910 44952 17970 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 17358 44952 17418 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 16806 44952 16866 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 6870 44952 6930 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 6318 44952 6378 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 5766 44952 5826 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 4662 44952 4722 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 4110 44952 4170 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3558 44952 3618 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11286 44952 11346 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 10734 44952 10794 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10182 44952 10242 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 9078 44952 9138 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8526 44952 8586 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7974 44952 8034 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 15702 44952 15762 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 15150 44952 15210 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 14598 44952 14658 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 13494 44952 13554 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 12942 44952 13002 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 12390 44952 12450 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 28560 1000 28960 44152 1 FreeSans 400 0 0 0 VAPWR
port 53 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 29072 45152
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1723353804
<< error_p >>
rect -29 122 29 128
rect -29 88 -17 122
rect -29 82 29 88
rect -29 -88 29 -82
rect -29 -122 -17 -88
rect -29 -128 29 -122
<< pwell >>
rect -211 -260 211 260
<< nmos >>
rect -15 -50 15 50
<< ndiff >>
rect -73 38 -15 50
rect -73 -38 -61 38
rect -27 -38 -15 38
rect -73 -50 -15 -38
rect 15 38 73 50
rect 15 -38 27 38
rect 61 -38 73 38
rect 15 -50 73 -38
<< ndiffc >>
rect -61 -38 -27 38
rect 27 -38 61 38
<< psubdiff >>
rect -175 190 -79 224
rect 79 190 175 224
rect -175 128 -141 190
rect 141 128 175 190
rect -175 -190 -141 -128
rect 141 -190 175 -128
rect -175 -224 -79 -190
rect 79 -224 175 -190
<< psubdiffcont >>
rect -79 190 79 224
rect -175 -128 -141 128
rect 141 -128 175 128
rect -79 -224 79 -190
<< poly >>
rect -33 122 33 138
rect -33 88 -17 122
rect 17 88 33 122
rect -33 72 33 88
rect -15 50 15 72
rect -15 -72 15 -50
rect -33 -88 33 -72
rect -33 -122 -17 -88
rect 17 -122 33 -88
rect -33 -138 33 -122
<< polycont >>
rect -17 88 17 122
rect -17 -122 17 -88
<< locali >>
rect -175 190 -79 224
rect 79 190 175 224
rect -175 128 -141 190
rect 141 128 175 190
rect -33 88 -17 122
rect 17 88 33 122
rect -61 38 -27 54
rect -61 -54 -27 -38
rect 27 38 61 54
rect 27 -54 61 -38
rect -33 -122 -17 -88
rect 17 -122 33 -88
rect -175 -190 -141 -128
rect 141 -190 175 -128
rect -175 -224 -79 -190
rect 79 -224 175 -190
<< viali >>
rect -17 88 17 122
rect -61 -38 -27 38
rect 27 -38 61 38
rect -17 -122 17 -88
<< metal1 >>
rect -29 122 29 128
rect -29 88 -17 122
rect 17 88 29 122
rect -29 82 29 88
rect -67 38 -21 50
rect -67 -38 -61 38
rect -27 -38 -21 38
rect -67 -50 -21 -38
rect 21 38 67 50
rect 21 -38 27 38
rect 61 -38 67 38
rect 21 -50 67 -38
rect -29 -88 29 -82
rect -29 -122 -17 -88
rect 17 -122 29 -88
rect -29 -128 29 -122
<< properties >>
string FIXED_BBOX -158 -207 158 207
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.5 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

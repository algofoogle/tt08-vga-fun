magic
tech sky130A
magscale 1 2
timestamp 1723498766
<< error_p >>
rect -29 131 29 137
rect -29 97 -17 131
rect -29 91 29 97
rect -29 -97 29 -91
rect -29 -131 -17 -97
rect -29 -137 29 -131
<< nwell >>
rect -211 -269 211 269
<< pmos >>
rect -15 -50 15 50
<< pdiff >>
rect -73 38 -15 50
rect -73 -38 -61 38
rect -27 -38 -15 38
rect -73 -50 -15 -38
rect 15 38 73 50
rect 15 -38 27 38
rect 61 -38 73 38
rect 15 -50 73 -38
<< pdiffc >>
rect -61 -38 -27 38
rect 27 -38 61 38
<< nsubdiff >>
rect -175 199 -79 233
rect 79 199 175 233
rect -175 137 -141 199
rect 141 137 175 199
rect -175 -199 -141 -137
rect 141 -199 175 -137
rect -175 -233 -79 -199
rect 79 -233 175 -199
<< nsubdiffcont >>
rect -79 199 79 233
rect -175 -137 -141 137
rect 141 -137 175 137
rect -79 -233 79 -199
<< poly >>
rect -33 131 33 147
rect -33 97 -17 131
rect 17 97 33 131
rect -33 81 33 97
rect -15 50 15 81
rect -15 -81 15 -50
rect -33 -97 33 -81
rect -33 -131 -17 -97
rect 17 -131 33 -97
rect -33 -147 33 -131
<< polycont >>
rect -17 97 17 131
rect -17 -131 17 -97
<< locali >>
rect -175 199 -79 233
rect 79 199 175 233
rect -175 137 -141 199
rect 141 137 175 199
rect -33 97 -17 131
rect 17 97 33 131
rect -61 38 -27 54
rect -61 -54 -27 -38
rect 27 38 61 54
rect 27 -54 61 -38
rect -33 -131 -17 -97
rect 17 -131 33 -97
rect -175 -199 -141 -137
rect 141 -199 175 -137
rect -175 -233 -79 -199
rect 79 -233 175 -199
<< viali >>
rect -17 97 17 131
rect -61 -38 -27 38
rect 27 -38 61 38
rect -17 -131 17 -97
<< metal1 >>
rect -29 131 29 137
rect -29 97 -17 131
rect 17 97 29 131
rect -29 91 29 97
rect -67 38 -21 50
rect -67 -38 -61 38
rect -27 -38 -21 38
rect -67 -50 -21 -38
rect 21 38 67 50
rect 21 -38 27 38
rect 61 -38 67 38
rect 21 -50 67 -38
rect -29 -97 29 -91
rect -29 -131 -17 -97
rect 17 -131 29 -97
rect -29 -137 29 -131
<< properties >>
string FIXED_BBOX -158 -216 158 216
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.5 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1724386042
<< metal1 >>
rect 2808 17462 2814 17518
rect 2870 17462 2876 17518
rect 3176 17462 3182 17518
rect 3238 17462 3244 17518
rect 3544 17462 3550 17518
rect 3606 17462 3612 17518
rect 3912 17462 3918 17518
rect 3974 17462 3980 17518
rect 4280 17462 4286 17518
rect 4342 17462 4348 17518
rect 4648 17462 4654 17518
rect 4710 17462 4716 17518
rect 5016 17462 5022 17518
rect 5078 17462 5084 17518
rect 5384 17462 5390 17518
rect 5446 17462 5452 17518
rect 5752 17462 5758 17518
rect 5814 17462 5820 17518
rect 6120 17462 6126 17518
rect 6182 17462 6188 17518
rect 6488 17462 6494 17518
rect 6550 17462 6556 17518
rect 6856 17462 6862 17518
rect 6918 17462 6924 17518
rect 7224 17462 7230 17518
rect 7286 17462 7292 17518
rect 7592 17462 7598 17518
rect 7654 17462 7660 17518
rect 7960 17462 7966 17518
rect 8022 17462 8028 17518
rect 8328 17462 8334 17518
rect 8390 17462 8396 17518
rect 11648 17462 11654 17518
rect 11710 17462 11716 17518
rect 12016 17462 12022 17518
rect 12078 17462 12084 17518
rect 12384 17462 12390 17518
rect 12446 17462 12452 17518
rect 12752 17462 12758 17518
rect 12814 17462 12820 17518
rect 13120 17462 13126 17518
rect 13182 17462 13188 17518
rect 13488 17462 13494 17518
rect 13550 17462 13556 17518
rect 13856 17462 13862 17518
rect 13918 17462 13924 17518
rect 14224 17462 14230 17518
rect 14286 17462 14292 17518
rect 14592 17462 14598 17518
rect 14654 17462 14660 17518
rect 14960 17462 14966 17518
rect 15022 17462 15028 17518
rect 15328 17462 15334 17518
rect 15390 17462 15396 17518
rect 15696 17462 15702 17518
rect 15758 17462 15764 17518
rect 16064 17462 16070 17518
rect 16126 17462 16132 17518
rect 16432 17462 16438 17518
rect 16494 17462 16500 17518
rect 16800 17462 16806 17518
rect 16862 17462 16868 17518
rect 17168 17462 17174 17518
rect 17230 17462 17236 17518
<< via1 >>
rect 2814 17462 2870 17518
rect 3182 17462 3238 17518
rect 3550 17462 3606 17518
rect 3918 17462 3974 17518
rect 4286 17462 4342 17518
rect 4654 17462 4710 17518
rect 5022 17462 5078 17518
rect 5390 17462 5446 17518
rect 5758 17462 5814 17518
rect 6126 17462 6182 17518
rect 6494 17462 6550 17518
rect 6862 17462 6918 17518
rect 7230 17462 7286 17518
rect 7598 17462 7654 17518
rect 7966 17462 8022 17518
rect 8334 17462 8390 17518
rect 11654 17462 11710 17518
rect 12022 17462 12078 17518
rect 12390 17462 12446 17518
rect 12758 17462 12814 17518
rect 13126 17462 13182 17518
rect 13494 17462 13550 17518
rect 13862 17462 13918 17518
rect 14230 17462 14286 17518
rect 14598 17462 14654 17518
rect 14966 17462 15022 17518
rect 15334 17462 15390 17518
rect 15702 17462 15758 17518
rect 16070 17462 16126 17518
rect 16438 17462 16494 17518
rect 16806 17462 16862 17518
rect 17174 17462 17230 17518
rect 20494 17472 20550 17528
rect 20862 17472 20918 17528
rect 21230 17472 21286 17528
rect 21598 17472 21654 17528
rect 21966 17472 22022 17528
rect 22334 17472 22390 17528
rect 22702 17472 22758 17528
rect 23070 17472 23126 17528
rect 23438 17472 23494 17528
rect 23806 17472 23862 17528
rect 24174 17472 24230 17528
rect 24542 17472 24598 17528
rect 24910 17472 24966 17528
rect 25278 17472 25334 17528
rect 25646 17472 25702 17528
rect 26014 17472 26070 17528
<< metal2 >>
rect 10704 44870 10824 44900
rect 10704 44810 10732 44870
rect 10792 44810 10824 44870
rect 10704 44780 10824 44810
rect 11256 44870 11376 44900
rect 11256 44810 11284 44870
rect 11344 44810 11376 44870
rect 11256 44780 11376 44810
rect 11808 44870 11928 44900
rect 11808 44810 11836 44870
rect 11896 44810 11928 44870
rect 11808 44780 11928 44810
rect 12360 44870 12480 44900
rect 12360 44810 12388 44870
rect 12448 44810 12480 44870
rect 12360 44780 12480 44810
rect 12912 44870 13032 44900
rect 12912 44810 12940 44870
rect 13000 44810 13032 44870
rect 12912 44780 13032 44810
rect 13464 44870 13584 44900
rect 13464 44810 13492 44870
rect 13552 44810 13584 44870
rect 13464 44780 13584 44810
rect 14016 44870 14136 44900
rect 14016 44810 14044 44870
rect 14104 44810 14136 44870
rect 14016 44780 14136 44810
rect 14568 44870 14688 44900
rect 14568 44810 14596 44870
rect 14656 44810 14688 44870
rect 14568 44780 14688 44810
rect 15120 44870 15240 44900
rect 15120 44810 15148 44870
rect 15208 44810 15240 44870
rect 15120 44780 15240 44810
rect 15672 44870 15792 44900
rect 15672 44810 15700 44870
rect 15760 44810 15792 44870
rect 15672 44780 15792 44810
rect 20640 44870 20760 44900
rect 20640 44810 20668 44870
rect 20728 44810 20760 44870
rect 20640 44780 20760 44810
rect 21192 44870 21312 44900
rect 21192 44810 21220 44870
rect 21280 44810 21312 44870
rect 21192 44780 21312 44810
rect 21744 44870 21864 44900
rect 21744 44810 21772 44870
rect 21832 44810 21864 44870
rect 21744 44780 21864 44810
rect 22296 44870 22416 44900
rect 22296 44810 22324 44870
rect 22384 44810 22416 44870
rect 22296 44780 22416 44810
rect 22848 44870 22968 44900
rect 22848 44810 22876 44870
rect 22936 44810 22968 44870
rect 22848 44780 22968 44810
rect 23400 44870 23520 44900
rect 23400 44810 23428 44870
rect 23488 44810 23520 44870
rect 23400 44780 23520 44810
rect 23952 44870 24072 44900
rect 23952 44810 23980 44870
rect 24040 44810 24072 44870
rect 23952 44780 24072 44810
rect 24504 44870 24624 44900
rect 24504 44810 24532 44870
rect 24592 44810 24624 44870
rect 24504 44780 24624 44810
rect 25056 44870 25176 44900
rect 25056 44810 25084 44870
rect 25144 44810 25176 44870
rect 25056 44780 25176 44810
rect 25608 44870 25728 44900
rect 25608 44810 25636 44870
rect 25696 44810 25728 44870
rect 25608 44780 25728 44810
rect 10734 42962 10790 44780
rect 11286 42962 11342 44780
rect 11838 42962 11894 44780
rect 12390 42962 12446 44780
rect 12942 42962 12998 44780
rect 13494 42962 13550 44780
rect 14046 42962 14102 44780
rect 14598 42962 14654 44780
rect 15150 42962 15206 44780
rect 15702 42962 15758 44780
rect 20670 42962 20726 44780
rect 21222 42962 21278 44780
rect 21774 42962 21830 44780
rect 22326 42962 22382 44780
rect 22878 42962 22934 44780
rect 23430 42962 23486 44780
rect 23982 42962 24038 44780
rect 24534 42962 24590 44780
rect 25086 42962 25142 44780
rect 25638 42962 25694 44780
rect 2814 17518 2870 19248
rect 2814 17456 2870 17462
rect 3182 17518 3238 19248
rect 3182 17456 3238 17462
rect 3550 17518 3606 19248
rect 3550 17456 3606 17462
rect 3918 17518 3974 19248
rect 3918 17456 3974 17462
rect 4286 17518 4342 19248
rect 4286 17456 4342 17462
rect 4654 17518 4710 19248
rect 4654 17456 4710 17462
rect 5022 17518 5078 19248
rect 5022 17456 5078 17462
rect 5390 17518 5446 19248
rect 5390 17456 5446 17462
rect 5758 17518 5814 19248
rect 5758 17456 5814 17462
rect 6126 17518 6182 19248
rect 6126 17456 6182 17462
rect 6494 17518 6550 19248
rect 6494 17456 6550 17462
rect 6862 17518 6918 19248
rect 6862 17456 6918 17462
rect 7230 17518 7286 19248
rect 7230 17456 7286 17462
rect 7598 17518 7654 19248
rect 7598 17456 7654 17462
rect 7966 17518 8022 19248
rect 7966 17456 8022 17462
rect 8334 17518 8390 19248
rect 8334 17456 8390 17462
rect 11654 17518 11710 19248
rect 11654 17456 11710 17462
rect 12022 17518 12078 19248
rect 12022 17456 12078 17462
rect 12390 17518 12446 19248
rect 12390 17456 12446 17462
rect 12758 17518 12814 19248
rect 12758 17456 12814 17462
rect 13126 17518 13182 19248
rect 13126 17456 13182 17462
rect 13494 17518 13550 19248
rect 13494 17456 13550 17462
rect 13862 17518 13918 19248
rect 13862 17456 13918 17462
rect 14230 17518 14286 19248
rect 14230 17456 14286 17462
rect 14598 17518 14654 19248
rect 14598 17456 14654 17462
rect 14966 17518 15022 19248
rect 14966 17456 15022 17462
rect 15334 17518 15390 19248
rect 15334 17456 15390 17462
rect 15702 17518 15758 19248
rect 15702 17456 15758 17462
rect 16070 17518 16126 19248
rect 16070 17456 16126 17462
rect 16438 17518 16494 19248
rect 16438 17456 16494 17462
rect 16806 17518 16862 19248
rect 16806 17456 16862 17462
rect 17174 17518 17230 19248
rect 20494 17528 20550 19380
rect 20494 17466 20550 17472
rect 20862 17528 20918 19380
rect 20862 17466 20918 17472
rect 21230 17528 21286 19380
rect 21230 17466 21286 17472
rect 21598 17528 21654 19380
rect 21598 17466 21654 17472
rect 21966 17528 22022 19380
rect 21966 17466 22022 17472
rect 22334 17528 22390 19380
rect 22334 17466 22390 17472
rect 22702 17528 22758 19380
rect 22702 17466 22758 17472
rect 23070 17528 23126 19380
rect 23070 17466 23126 17472
rect 23438 17528 23494 19380
rect 23438 17466 23494 17472
rect 23806 17528 23862 19380
rect 23806 17466 23862 17472
rect 24174 17528 24230 19380
rect 24174 17466 24230 17472
rect 24542 17528 24598 19380
rect 24542 17466 24598 17472
rect 24910 17528 24966 19380
rect 24910 17466 24966 17472
rect 25278 17528 25334 19380
rect 25278 17466 25334 17472
rect 25646 17528 25702 19380
rect 25646 17466 25702 17472
rect 26014 17528 26070 19380
rect 26014 17466 26070 17472
rect 17174 17456 17230 17462
<< via2 >>
rect 10732 44810 10792 44870
rect 11284 44810 11344 44870
rect 11836 44810 11896 44870
rect 12388 44810 12448 44870
rect 12940 44810 13000 44870
rect 13492 44810 13552 44870
rect 14044 44810 14104 44870
rect 14596 44810 14656 44870
rect 15148 44810 15208 44870
rect 15700 44810 15760 44870
rect 20668 44810 20728 44870
rect 21220 44810 21280 44870
rect 21772 44810 21832 44870
rect 22324 44810 22384 44870
rect 22876 44810 22936 44870
rect 23428 44810 23488 44870
rect 23980 44810 24040 44870
rect 24532 44810 24592 44870
rect 25084 44810 25144 44870
rect 25636 44810 25696 44870
<< metal3 >>
rect 10704 44875 10824 44900
rect 6310 44798 6316 44862
rect 6380 44798 6386 44862
rect 6862 44798 6868 44862
rect 6932 44798 6938 44862
rect 10704 44805 10727 44875
rect 10797 44805 10824 44875
rect 6318 43528 6378 44798
rect 6870 43528 6930 44798
rect 10704 44780 10824 44805
rect 11256 44875 11376 44900
rect 11256 44805 11279 44875
rect 11349 44805 11376 44875
rect 11256 44780 11376 44805
rect 11808 44875 11928 44900
rect 11808 44805 11831 44875
rect 11901 44805 11928 44875
rect 11808 44780 11928 44805
rect 12360 44875 12480 44900
rect 12360 44805 12383 44875
rect 12453 44805 12480 44875
rect 12360 44780 12480 44805
rect 12912 44875 13032 44900
rect 12912 44805 12935 44875
rect 13005 44805 13032 44875
rect 12912 44780 13032 44805
rect 13464 44875 13584 44900
rect 13464 44805 13487 44875
rect 13557 44805 13584 44875
rect 13464 44780 13584 44805
rect 14016 44875 14136 44900
rect 14016 44805 14039 44875
rect 14109 44805 14136 44875
rect 14016 44780 14136 44805
rect 14568 44875 14688 44900
rect 14568 44805 14591 44875
rect 14661 44805 14688 44875
rect 14568 44780 14688 44805
rect 15120 44875 15240 44900
rect 15120 44805 15143 44875
rect 15213 44805 15240 44875
rect 15120 44780 15240 44805
rect 15672 44875 15792 44900
rect 15672 44805 15695 44875
rect 15765 44805 15792 44875
rect 15672 44780 15792 44805
rect 20640 44875 20760 44900
rect 20640 44805 20663 44875
rect 20733 44805 20760 44875
rect 20640 44780 20760 44805
rect 21192 44875 21312 44900
rect 21192 44805 21215 44875
rect 21285 44805 21312 44875
rect 21192 44780 21312 44805
rect 21744 44875 21864 44900
rect 21744 44805 21767 44875
rect 21837 44805 21864 44875
rect 21744 44780 21864 44805
rect 22296 44875 22416 44900
rect 22296 44805 22319 44875
rect 22389 44805 22416 44875
rect 22296 44780 22416 44805
rect 22848 44875 22968 44900
rect 22848 44805 22871 44875
rect 22941 44805 22968 44875
rect 22848 44780 22968 44805
rect 23400 44875 23520 44900
rect 23400 44805 23423 44875
rect 23493 44805 23520 44875
rect 23400 44780 23520 44805
rect 23952 44875 24072 44900
rect 23952 44805 23975 44875
rect 24045 44805 24072 44875
rect 23952 44780 24072 44805
rect 24504 44875 24624 44900
rect 24504 44805 24527 44875
rect 24597 44805 24624 44875
rect 24504 44780 24624 44805
rect 25056 44875 25176 44900
rect 25056 44805 25079 44875
rect 25149 44805 25176 44875
rect 25056 44780 25176 44805
rect 25608 44875 25728 44900
rect 25608 44805 25631 44875
rect 25701 44805 25728 44875
rect 25608 44780 25728 44805
rect 7220 44660 7620 44666
rect 6316 43522 6380 43528
rect 6316 43452 6380 43458
rect 6868 43522 6932 43528
rect 6868 43452 6932 43458
rect 7220 43099 7620 44260
rect 12788 44660 13188 44666
rect 12788 43099 13188 44260
rect 18788 44660 19188 44666
rect 18788 43099 19188 44260
rect 24788 44660 25188 44666
rect 24788 43099 25188 44260
rect 7220 42701 7221 43099
rect 7619 42701 7620 43099
rect 12783 42701 12789 43099
rect 13187 42701 13193 43099
rect 18783 42701 18789 43099
rect 19187 42701 19193 43099
rect 24783 42701 24789 43099
rect 25187 42701 25193 43099
rect 7220 42700 7620 42701
rect 12788 42700 13188 42701
rect 18788 42700 19188 42701
rect 24788 42700 25188 42701
rect 7221 42695 7619 42700
rect 3789 18870 4187 18875
rect 1070 18869 27360 18870
rect 1070 18471 3789 18869
rect 4187 18850 27360 18869
rect 4187 18490 9830 18850
rect 10170 18490 15810 18850
rect 16170 18490 21810 18850
rect 22170 18490 26980 18850
rect 27340 18490 27360 18850
rect 4187 18471 27360 18490
rect 1070 18470 27360 18471
rect 1070 16569 1270 18470
rect 3789 18465 4187 18470
rect 1070 16371 1071 16569
rect 1269 16371 1270 16569
rect 1070 16370 1270 16371
rect 9520 16569 9720 18470
rect 9520 16371 9521 16569
rect 9719 16371 9720 16569
rect 9520 16370 9720 16371
rect 18490 16569 18690 18470
rect 26450 18270 28360 18290
rect 26450 17910 26470 18270
rect 26830 17910 27980 18270
rect 28340 17910 28360 18270
rect 26450 17890 28360 17910
rect 18490 16371 18491 16569
rect 18689 16371 18690 16569
rect 18490 16370 18690 16371
rect 1071 16365 1269 16370
rect 9521 16365 9719 16370
rect 18491 16365 18689 16370
<< via3 >>
rect 6316 44798 6380 44862
rect 6868 44798 6932 44862
rect 10727 44870 10797 44875
rect 10727 44810 10732 44870
rect 10732 44810 10792 44870
rect 10792 44810 10797 44870
rect 10727 44805 10797 44810
rect 11279 44870 11349 44875
rect 11279 44810 11284 44870
rect 11284 44810 11344 44870
rect 11344 44810 11349 44870
rect 11279 44805 11349 44810
rect 11831 44870 11901 44875
rect 11831 44810 11836 44870
rect 11836 44810 11896 44870
rect 11896 44810 11901 44870
rect 11831 44805 11901 44810
rect 12383 44870 12453 44875
rect 12383 44810 12388 44870
rect 12388 44810 12448 44870
rect 12448 44810 12453 44870
rect 12383 44805 12453 44810
rect 12935 44870 13005 44875
rect 12935 44810 12940 44870
rect 12940 44810 13000 44870
rect 13000 44810 13005 44870
rect 12935 44805 13005 44810
rect 13487 44870 13557 44875
rect 13487 44810 13492 44870
rect 13492 44810 13552 44870
rect 13552 44810 13557 44870
rect 13487 44805 13557 44810
rect 14039 44870 14109 44875
rect 14039 44810 14044 44870
rect 14044 44810 14104 44870
rect 14104 44810 14109 44870
rect 14039 44805 14109 44810
rect 14591 44870 14661 44875
rect 14591 44810 14596 44870
rect 14596 44810 14656 44870
rect 14656 44810 14661 44870
rect 14591 44805 14661 44810
rect 15143 44870 15213 44875
rect 15143 44810 15148 44870
rect 15148 44810 15208 44870
rect 15208 44810 15213 44870
rect 15143 44805 15213 44810
rect 15695 44870 15765 44875
rect 15695 44810 15700 44870
rect 15700 44810 15760 44870
rect 15760 44810 15765 44870
rect 15695 44805 15765 44810
rect 20663 44870 20733 44875
rect 20663 44810 20668 44870
rect 20668 44810 20728 44870
rect 20728 44810 20733 44870
rect 20663 44805 20733 44810
rect 21215 44870 21285 44875
rect 21215 44810 21220 44870
rect 21220 44810 21280 44870
rect 21280 44810 21285 44870
rect 21215 44805 21285 44810
rect 21767 44870 21837 44875
rect 21767 44810 21772 44870
rect 21772 44810 21832 44870
rect 21832 44810 21837 44870
rect 21767 44805 21837 44810
rect 22319 44870 22389 44875
rect 22319 44810 22324 44870
rect 22324 44810 22384 44870
rect 22384 44810 22389 44870
rect 22319 44805 22389 44810
rect 22871 44870 22941 44875
rect 22871 44810 22876 44870
rect 22876 44810 22936 44870
rect 22936 44810 22941 44870
rect 22871 44805 22941 44810
rect 23423 44870 23493 44875
rect 23423 44810 23428 44870
rect 23428 44810 23488 44870
rect 23488 44810 23493 44870
rect 23423 44805 23493 44810
rect 23975 44870 24045 44875
rect 23975 44810 23980 44870
rect 23980 44810 24040 44870
rect 24040 44810 24045 44870
rect 23975 44805 24045 44810
rect 24527 44870 24597 44875
rect 24527 44810 24532 44870
rect 24532 44810 24592 44870
rect 24592 44810 24597 44870
rect 24527 44805 24597 44810
rect 25079 44870 25149 44875
rect 25079 44810 25084 44870
rect 25084 44810 25144 44870
rect 25144 44810 25149 44870
rect 25079 44805 25149 44810
rect 25631 44870 25701 44875
rect 25631 44810 25636 44870
rect 25636 44810 25696 44870
rect 25696 44810 25701 44870
rect 25631 44805 25701 44810
rect 7220 44260 7620 44660
rect 6316 43458 6380 43522
rect 6868 43458 6932 43522
rect 12788 44260 13188 44660
rect 18788 44260 19188 44660
rect 24788 44260 25188 44660
rect 7221 42701 7619 43099
rect 12789 42701 13187 43099
rect 18789 42701 19187 43099
rect 24789 42701 25187 43099
rect 3789 18471 4187 18869
rect 9830 18490 10170 18850
rect 15810 18490 16170 18850
rect 21810 18490 22170 18850
rect 26980 18490 27340 18850
rect 1071 16371 1269 16569
rect 9521 16371 9719 16569
rect 26470 17910 26830 18270
rect 27980 17910 28340 18270
rect 18491 16371 18689 16569
<< metal4 >>
rect 3006 44660 3066 45152
rect 3558 44660 3618 45152
rect 4110 44660 4170 45152
rect 4662 44660 4722 45152
rect 5214 44660 5274 45152
rect 5766 44660 5826 45152
rect 6318 44863 6378 45152
rect 6870 44863 6930 45152
rect 6315 44862 6381 44863
rect 6315 44798 6316 44862
rect 6380 44798 6381 44862
rect 6315 44797 6381 44798
rect 6867 44862 6933 44863
rect 6867 44798 6868 44862
rect 6932 44798 6933 44862
rect 6867 44797 6933 44798
rect 7422 44661 7482 45152
rect 7219 44660 7621 44661
rect 7974 44660 8034 45152
rect 8526 44660 8586 45152
rect 9078 44660 9138 45152
rect 9630 44660 9690 45152
rect 10182 44660 10242 45152
rect 10734 45010 10794 45152
rect 11286 45010 11346 45152
rect 11838 45010 11898 45152
rect 12390 45010 12450 45152
rect 12942 45010 13002 45152
rect 13494 45010 13554 45152
rect 14046 45010 14106 45152
rect 14598 45010 14658 45152
rect 15150 45010 15210 45152
rect 15702 45010 15762 45152
rect 10724 44900 10804 45010
rect 11276 44900 11356 45010
rect 11828 44900 11908 45010
rect 12380 44900 12460 45010
rect 12932 44900 13012 45010
rect 13484 44900 13564 45010
rect 14036 44900 14116 45010
rect 14588 44900 14668 45010
rect 15140 44900 15220 45010
rect 15692 44900 15772 45010
rect 16254 44952 16314 45152
rect 16806 44952 16866 45152
rect 17358 44952 17418 45152
rect 17910 44952 17970 45152
rect 18462 44952 18522 45152
rect 19014 44952 19074 45152
rect 19566 44952 19626 45152
rect 20118 44952 20178 45152
rect 20670 45010 20730 45152
rect 21222 45010 21282 45152
rect 21774 45010 21834 45152
rect 22326 45010 22386 45152
rect 22878 45010 22938 45152
rect 23430 45010 23490 45152
rect 23982 45010 24042 45152
rect 24534 45010 24594 45152
rect 25086 45010 25146 45152
rect 25638 45010 25698 45152
rect 20660 44900 20740 45010
rect 21212 44900 21292 45010
rect 21764 44900 21844 45010
rect 22316 44900 22396 45010
rect 22868 44900 22948 45010
rect 23420 44900 23500 45010
rect 23972 44900 24052 45010
rect 24524 44900 24604 45010
rect 25076 44900 25156 45010
rect 25628 44900 25708 45010
rect 26190 44952 26250 45152
rect 10704 44875 10824 44900
rect 10704 44805 10727 44875
rect 10797 44805 10824 44875
rect 10704 44780 10824 44805
rect 11256 44875 11376 44900
rect 11256 44805 11279 44875
rect 11349 44805 11376 44875
rect 11256 44780 11376 44805
rect 11808 44875 11928 44900
rect 11808 44805 11831 44875
rect 11901 44805 11928 44875
rect 11808 44780 11928 44805
rect 12360 44875 12480 44900
rect 12360 44805 12383 44875
rect 12453 44805 12480 44875
rect 12360 44780 12480 44805
rect 12912 44875 13032 44900
rect 12912 44805 12935 44875
rect 13005 44805 13032 44875
rect 12912 44780 13032 44805
rect 13464 44875 13584 44900
rect 13464 44805 13487 44875
rect 13557 44805 13584 44875
rect 13464 44780 13584 44805
rect 14016 44875 14136 44900
rect 14016 44805 14039 44875
rect 14109 44805 14136 44875
rect 14016 44780 14136 44805
rect 14568 44875 14688 44900
rect 14568 44805 14591 44875
rect 14661 44805 14688 44875
rect 14568 44780 14688 44805
rect 15120 44875 15240 44900
rect 15120 44805 15143 44875
rect 15213 44805 15240 44875
rect 15120 44780 15240 44805
rect 15672 44875 15792 44900
rect 15672 44805 15695 44875
rect 15765 44805 15792 44875
rect 15672 44780 15792 44805
rect 20640 44875 20760 44900
rect 20640 44805 20663 44875
rect 20733 44805 20760 44875
rect 20640 44780 20760 44805
rect 21192 44875 21312 44900
rect 21192 44805 21215 44875
rect 21285 44805 21312 44875
rect 21192 44780 21312 44805
rect 21744 44875 21864 44900
rect 21744 44805 21767 44875
rect 21837 44805 21864 44875
rect 21744 44780 21864 44805
rect 22296 44875 22416 44900
rect 22296 44805 22319 44875
rect 22389 44805 22416 44875
rect 22296 44780 22416 44805
rect 22848 44875 22968 44900
rect 22848 44805 22871 44875
rect 22941 44805 22968 44875
rect 22848 44780 22968 44805
rect 23400 44875 23520 44900
rect 23400 44805 23423 44875
rect 23493 44805 23520 44875
rect 23400 44780 23520 44805
rect 23952 44875 24072 44900
rect 23952 44805 23975 44875
rect 24045 44805 24072 44875
rect 23952 44780 24072 44805
rect 24504 44875 24624 44900
rect 24504 44805 24527 44875
rect 24597 44805 24624 44875
rect 24504 44780 24624 44805
rect 25056 44875 25176 44900
rect 25056 44805 25079 44875
rect 25149 44805 25176 44875
rect 25056 44780 25176 44805
rect 25608 44875 25728 44900
rect 25608 44805 25631 44875
rect 25701 44805 25728 44875
rect 25608 44780 25728 44805
rect 12787 44660 13189 44661
rect 18787 44660 19189 44661
rect 24787 44660 25189 44661
rect 26330 44660 28360 44860
rect 2950 44260 7220 44660
rect 7620 44260 12788 44660
rect 13188 44260 18788 44660
rect 19188 44260 24788 44660
rect 25188 44460 28360 44660
rect 25188 44260 26730 44460
rect 7219 44259 7621 44260
rect 12787 44259 13189 44260
rect 18787 44259 19189 44260
rect 24787 44259 25189 44260
rect 26960 43620 27560 44160
rect 3790 43522 27560 43620
rect 3790 43458 6316 43522
rect 6380 43458 6868 43522
rect 6932 43458 27560 43522
rect 3790 43400 27560 43458
rect 3788 43220 27560 43400
rect 3788 42060 4188 43220
rect 6788 43099 7620 43100
rect 6788 42701 7221 43099
rect 7619 42701 7620 43099
rect 6788 42700 7620 42701
rect 6788 42030 7188 42700
rect 9788 42040 10188 43220
rect 12788 43099 13188 43100
rect 12788 42701 12789 43099
rect 13187 42701 13188 43099
rect 12788 42040 13188 42701
rect 15788 42030 16188 43220
rect 18788 43099 19188 43100
rect 18788 42701 18789 43099
rect 19187 42701 19188 43099
rect 18788 42044 19188 42701
rect 21788 42050 22188 43220
rect 24788 43099 25188 43100
rect 24788 42701 24789 43099
rect 25187 42701 25188 43099
rect 24788 42044 25188 42701
rect 3788 18869 4188 19980
rect 3788 18471 3789 18869
rect 4187 18471 4188 18869
rect 3788 18470 4188 18471
rect 6788 18290 7188 20060
rect 9788 18850 10188 19980
rect 9788 18490 9830 18850
rect 10170 18490 10188 18850
rect 9788 18470 10188 18490
rect 12788 18290 13188 20060
rect 15788 18850 16188 19980
rect 15788 18490 15810 18850
rect 16170 18490 16188 18850
rect 15788 18470 16188 18490
rect 18788 18290 19188 20060
rect 21788 18850 22188 19980
rect 21788 18490 21810 18850
rect 22170 18490 22188 18850
rect 21788 18470 22188 18490
rect 24788 18290 25188 20060
rect 26960 18850 27560 43220
rect 26960 18490 26980 18850
rect 27340 18490 27560 18850
rect 680 18270 26850 18290
rect 680 17910 26470 18270
rect 26830 17910 26850 18270
rect 680 17890 26850 17910
rect 680 16170 880 17890
rect 1070 16569 1650 16570
rect 1070 16371 1071 16569
rect 1269 16371 1650 16569
rect 1070 16370 1650 16371
rect 9140 16170 9340 17890
rect 9520 16569 10440 16570
rect 9520 16371 9521 16569
rect 9719 16371 10440 16569
rect 9520 16370 10440 16371
rect 18160 16170 18360 17890
rect 18490 16569 19280 16570
rect 18490 16371 18491 16569
rect 18689 16371 19280 16569
rect 18490 16370 19280 16371
rect 680 15970 1730 16170
rect 9140 15970 10450 16170
rect 18160 15970 19320 16170
rect 25928 7188 26742 7352
rect 8230 700 8410 1600
rect 8230 520 15822 700
rect 17078 692 17242 1602
rect 25916 694 26084 1604
rect 17078 528 19682 692
rect 186 0 366 200
rect 4050 0 4230 200
rect 7914 0 8094 200
rect 11778 0 11958 200
rect 15642 0 15822 520
rect 19518 200 19682 528
rect 23376 526 26084 694
rect 26578 688 26742 7188
rect 26960 990 27560 18490
rect 27760 18270 28360 44460
rect 27760 17910 27980 18270
rect 28340 17910 28360 18270
rect 27760 1000 28360 17910
rect 28560 1000 28960 44152
rect 23376 200 23544 526
rect 26566 524 27402 688
rect 27238 200 27402 524
rect 19506 0 19686 200
rect 23370 0 23550 200
rect 27234 0 27414 200
use csdac_nom  B_dac
timestamp 1724369829
transform 1 0 1450 0 1 12370
box 0 -10950 6992 5196
use controller  controller_0
timestamp 1724295482
transform 1 0 2436 0 1 19084
box 386 0 23630 24000
use csdac_nom  G_dac
timestamp 1724369829
transform 1 0 10290 0 1 12370
box 0 -10950 6992 5196
use csdac_nom  R_dac
timestamp 1724369829
transform 1 0 19130 0 1 12370
box 0 -10950 6992 5196
<< labels >>
flabel metal4 s 25638 44952 25698 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 26190 44952 26250 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 27234 0 27414 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 23370 0 23550 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 19506 0 19686 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 15642 0 15822 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 11778 0 11958 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 7914 0 8094 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4050 0 4230 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 186 0 366 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 24534 44952 24594 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 23982 44952 24042 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 23430 44952 23490 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 22326 44952 22386 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 21774 44952 21834 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 21222 44952 21282 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 20118 44952 20178 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 19566 44952 19626 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 19014 44952 19074 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 17910 44952 17970 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 17358 44952 17418 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 16806 44952 16866 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 6870 44952 6930 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 6318 44952 6378 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 5766 44952 5826 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 4662 44952 4722 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 4110 44952 4170 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3558 44952 3618 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11286 44952 11346 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 10734 44952 10794 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10182 44952 10242 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 9078 44952 9138 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8526 44952 8586 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7974 44952 8034 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 15702 44952 15762 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 15150 44952 15210 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 14598 44952 14658 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 13494 44952 13554 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 12942 44952 13002 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 12390 44952 12450 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 27760 1000 28360 44152 1 FreeSans 1600 90 0 0 VGND
port 54 nsew ground bidirectional
flabel metal4 28560 1000 28960 44152 1 FreeSans 1600 90 0 0 VAPWR
port 55 nsew power bidirectional
flabel metal4 26960 1000 27560 44152 1 FreeSans 1600 90 0 0 VDPWR
port 51 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 29072 45152
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1723607196
<< error_s >>
rect 11230 -7470 11239 -7461
rect 11421 -7470 11430 -7461
rect 11221 -7479 11230 -7470
rect 11430 -7479 11439 -7470
rect 11221 -7670 11230 -7661
rect 11430 -7670 11439 -7661
rect 11230 -7679 11239 -7670
rect 11421 -7679 11430 -7670
rect 5053 -8814 5088 -8780
rect 5054 -8833 5088 -8814
rect 4884 -8882 4942 -8876
rect 4884 -8916 4896 -8882
rect 4884 -8922 4942 -8916
rect 4884 -9092 4942 -9086
rect 4884 -9126 4896 -9092
rect 4884 -9132 4942 -9126
rect 5073 -9228 5088 -8833
rect 5107 -8867 5142 -8833
rect 5422 -8867 5457 -8833
rect 5107 -9228 5141 -8867
rect 5423 -8886 5457 -8867
rect 5253 -8935 5311 -8929
rect 5253 -8969 5265 -8935
rect 5253 -8975 5311 -8969
rect 5253 -9145 5311 -9139
rect 5253 -9179 5265 -9145
rect 5253 -9185 5311 -9179
rect 5107 -9262 5122 -9228
rect 5442 -9281 5457 -8886
rect 5476 -8920 5511 -8886
rect 7361 -8920 7396 -8886
rect 5476 -9281 5510 -8920
rect 7362 -8939 7396 -8920
rect 5476 -9315 5491 -9281
rect 7381 -9334 7396 -8939
rect 7415 -8973 7450 -8939
rect 7730 -8973 7765 -8939
rect 7415 -9334 7449 -8973
rect 7731 -8992 7765 -8973
rect 7561 -9041 7619 -9035
rect 7561 -9075 7573 -9041
rect 7561 -9081 7619 -9075
rect 7561 -9251 7619 -9245
rect 7561 -9285 7573 -9251
rect 7561 -9291 7619 -9285
rect 7415 -9368 7430 -9334
rect 7750 -9387 7765 -8992
rect 7784 -9026 7819 -8992
rect 8099 -9026 8134 -8992
rect 7784 -9387 7818 -9026
rect 8100 -9045 8134 -9026
rect 7930 -9094 7988 -9088
rect 7930 -9128 7942 -9094
rect 7930 -9134 7988 -9128
rect 7930 -9304 7988 -9298
rect 7930 -9338 7942 -9304
rect 7930 -9344 7988 -9338
rect 7784 -9421 7799 -9387
rect 8119 -9440 8134 -9045
rect 8153 -9079 8188 -9045
rect 9238 -9079 9273 -9045
rect 8153 -9440 8187 -9079
rect 9239 -9098 9273 -9079
rect 8153 -9474 8168 -9440
rect 9258 -9493 9273 -9098
rect 9292 -9132 9327 -9098
rect 9607 -9132 9642 -9098
rect 9292 -9493 9326 -9132
rect 9608 -9151 9642 -9132
rect 9438 -9200 9496 -9194
rect 9438 -9234 9450 -9200
rect 9438 -9240 9496 -9234
rect 9438 -9410 9496 -9404
rect 9438 -9444 9450 -9410
rect 9438 -9450 9496 -9444
rect 9292 -9527 9307 -9493
rect 9627 -9546 9642 -9151
rect 9661 -9185 9696 -9151
rect 9976 -9185 10011 -9151
rect 9661 -9546 9695 -9185
rect 9977 -9204 10011 -9185
rect 9807 -9253 9865 -9247
rect 9807 -9287 9819 -9253
rect 9807 -9293 9865 -9287
rect 9807 -9463 9865 -9457
rect 9807 -9497 9819 -9463
rect 9807 -9503 9865 -9497
rect 9661 -9580 9676 -9546
rect 9996 -9599 10011 -9204
rect 10030 -9238 10065 -9204
rect 10735 -9238 10770 -9204
rect 10030 -9599 10064 -9238
rect 10736 -9257 10770 -9238
rect 10030 -9633 10045 -9599
rect 10755 -9652 10770 -9257
rect 10789 -9291 10824 -9257
rect 11104 -9291 11139 -9257
rect 10789 -9652 10823 -9291
rect 11105 -9310 11139 -9291
rect 10935 -9359 10993 -9353
rect 10935 -9393 10947 -9359
rect 10935 -9399 10993 -9393
rect 10935 -9569 10993 -9563
rect 10935 -9603 10947 -9569
rect 10935 -9609 10993 -9603
rect 10789 -9686 10804 -9652
rect 11124 -9705 11139 -9310
rect 11158 -9344 11193 -9310
rect 11473 -9344 11508 -9310
rect 11158 -9705 11192 -9344
rect 11474 -9363 11508 -9344
rect 11304 -9412 11362 -9406
rect 11304 -9446 11316 -9412
rect 11304 -9452 11362 -9446
rect 11304 -9622 11362 -9616
rect 11304 -9656 11316 -9622
rect 11304 -9662 11362 -9656
rect 11158 -9739 11173 -9705
rect 11493 -9758 11508 -9363
rect 11527 -9397 11562 -9363
rect 12012 -9397 12047 -9363
rect 11527 -9758 11561 -9397
rect 12013 -9416 12047 -9397
rect 11527 -9792 11542 -9758
rect 12032 -9811 12047 -9416
rect 12066 -9450 12101 -9416
rect 12381 -9450 12416 -9416
rect 12066 -9811 12100 -9450
rect 12382 -9469 12416 -9450
rect 12212 -9518 12270 -9512
rect 12212 -9552 12224 -9518
rect 12212 -9558 12270 -9552
rect 12212 -9728 12270 -9722
rect 12212 -9762 12224 -9728
rect 12212 -9768 12270 -9762
rect 12066 -9845 12081 -9811
rect 12401 -9864 12416 -9469
rect 12435 -9503 12470 -9469
rect 12435 -9864 12469 -9503
rect 12581 -9571 12639 -9565
rect 12581 -9605 12593 -9571
rect 12581 -9611 12639 -9605
rect 12581 -9781 12639 -9775
rect 12581 -9815 12593 -9781
rect 12581 -9821 12639 -9815
rect 12435 -9898 12450 -9864
rect 12770 -9917 12785 -9469
rect 12804 -9917 12838 -9415
rect 13550 -9475 13584 -9421
rect 12804 -9951 12819 -9917
rect 13569 -9970 13584 -9475
rect 13603 -9509 13638 -9475
rect 13918 -9509 13953 -9475
rect 13603 -9970 13637 -9509
rect 13919 -9528 13953 -9509
rect 13749 -9577 13807 -9571
rect 13749 -9611 13761 -9577
rect 13749 -9617 13807 -9611
rect 13749 -9887 13807 -9881
rect 13749 -9921 13761 -9887
rect 13749 -9927 13807 -9921
rect 13603 -10004 13618 -9970
rect 13938 -10023 13953 -9528
rect 13972 -9562 14007 -9528
rect 13972 -10023 14006 -9562
rect 14118 -9630 14176 -9624
rect 14118 -9664 14130 -9630
rect 14118 -9670 14176 -9664
rect 14118 -9940 14176 -9934
rect 14118 -9974 14130 -9940
rect 14118 -9980 14176 -9974
rect 13972 -10057 13987 -10023
<< viali >>
rect 940 5060 1120 5110
rect 1380 5050 1630 5100
rect 850 4720 900 5010
rect 1280 4960 1330 5010
rect 1280 4730 1330 4780
rect 1680 4730 1720 5000
rect 940 4630 1120 4680
rect 1510 4640 1630 4680
rect 2040 3050 2350 3100
rect 1790 2760 1840 3010
rect 1890 2570 2090 2710
rect 1890 1560 2050 1690
rect 1890 630 2050 680
rect 8560 -6085 8630 2855
rect 9940 -6090 10080 2850
rect 11390 -6085 11460 2855
<< metal1 >>
rect 1994 5696 2194 5896
rect 2394 5696 2594 5896
rect 2794 5696 2994 5896
rect 3194 5696 3394 5896
rect 3594 5696 3794 5896
rect 3994 5696 4194 5896
rect 4394 5696 4594 5896
rect 4794 5696 4994 5896
rect 5194 5696 5394 5896
rect 5594 5696 5794 5896
rect 5994 5696 6194 5896
rect 6394 5696 6594 5896
rect 6794 5696 6994 5896
rect 7194 5696 7394 5896
rect 7594 5696 7794 5896
rect 7994 5696 8194 5896
rect 840 5110 1140 5120
rect 840 5060 940 5110
rect 1120 5060 1140 5110
rect 840 5050 1140 5060
rect 1270 5100 1730 5110
rect 1270 5050 1380 5100
rect 1630 5050 1730 5100
rect 840 5010 910 5050
rect 1270 5040 1730 5050
rect 1270 5020 1350 5040
rect 840 4720 850 5010
rect 900 4920 910 5010
rect 990 4960 1280 5020
rect 1340 4960 1350 5020
rect 1670 5000 1730 5040
rect 990 4950 1350 4960
rect 1380 4950 1560 5000
rect 1380 4920 1460 4950
rect 1670 4920 1680 5000
rect 900 4820 1010 4920
rect 1050 4820 1460 4920
rect 1560 4820 1680 4920
rect 900 4720 910 4820
rect 990 4730 1280 4790
rect 1340 4730 1350 4790
rect 990 4720 1350 4730
rect 1380 4780 1460 4820
rect 1380 4730 1560 4780
rect 1670 4730 1680 4820
rect 1720 4730 1730 5000
rect 840 4690 910 4720
rect 840 4680 1140 4690
rect 840 4630 940 4680
rect 1120 4630 1140 4680
rect 0 4000 350 4200
rect 550 4000 556 4200
rect 840 4180 1140 4630
rect 840 4020 860 4180
rect 1120 4020 1140 4180
rect 840 4000 1140 4020
rect 0 3600 350 3800
rect 550 3600 556 3800
rect 1380 3370 1460 4730
rect 1670 4690 1730 4730
rect 1490 4680 1730 4690
rect 1490 4640 1510 4680
rect 1630 4640 1730 4680
rect 1490 4630 1730 4640
rect 1540 3800 1730 4630
rect 2060 4350 2120 5696
rect 2460 4500 2520 5696
rect 2460 4440 2860 4500
rect 2060 4290 2710 4350
rect 1540 3780 1850 3800
rect 1540 3620 1560 3780
rect 1820 3620 1850 3780
rect 1360 3350 1480 3370
rect 1360 3220 1380 3350
rect 1460 3220 1480 3350
rect 1360 3200 1480 3220
rect 1540 3010 1850 3620
rect 2030 3780 2360 3800
rect 2030 3620 2050 3780
rect 2340 3620 2360 3780
rect 1880 3340 1980 3350
rect 1880 3230 1890 3340
rect 1970 3230 1980 3340
rect 1880 3220 1980 3230
rect 1540 2760 1790 3010
rect 1840 2760 1850 3010
rect 1890 2830 1940 3220
rect 2030 3100 2360 3620
rect 2410 3340 2510 3350
rect 2410 3230 2420 3340
rect 2500 3230 2510 3340
rect 2410 3220 2510 3230
rect 2030 3050 2040 3100
rect 2350 3050 2360 3100
rect 2030 3000 2360 3050
rect 1970 2940 2390 3000
rect 2420 2830 2470 3220
rect 2650 3130 2710 4290
rect 2800 3130 2860 4440
rect 8970 4180 9590 4200
rect 8970 4020 8990 4180
rect 9570 4020 9590 4180
rect 8470 3780 8650 3800
rect 8470 3620 8490 3780
rect 8630 3620 8650 3780
rect 2644 3070 2650 3130
rect 2710 3070 2716 3130
rect 2794 3070 2800 3130
rect 2860 3070 2866 3130
rect 8470 2855 8650 3620
rect 1970 2770 2390 2830
rect 1540 2730 1850 2760
rect 1540 2710 2110 2730
rect 1540 2690 1890 2710
rect 1540 2580 1560 2690
rect 1670 2580 1890 2690
rect 1540 2570 1890 2580
rect 2090 2570 2110 2710
rect 1540 2560 2110 2570
rect 1930 2460 2030 2520
rect 2090 2460 2100 2520
rect 2170 2420 2380 2770
rect 690 2400 1950 2420
rect 690 1860 710 2400
rect 870 1860 1950 2400
rect 690 1840 1950 1860
rect 1990 1840 2380 2420
rect 1930 1740 2030 1800
rect 2090 1740 2100 1800
rect 1540 1690 2110 1700
rect 1540 1680 1890 1690
rect 1540 1570 1560 1680
rect 1670 1570 1890 1680
rect 1540 1560 1890 1570
rect 2050 1560 2110 1690
rect 1540 1550 2110 1560
rect 1930 1450 2030 1510
rect 2090 1450 2100 1510
rect 2170 1410 2380 1840
rect 290 1390 1950 1410
rect 290 850 310 1390
rect 470 850 1950 1390
rect 290 830 1950 850
rect 1990 830 2380 1410
rect 1540 750 1690 770
rect 1540 640 1560 750
rect 1670 690 1690 750
rect 1930 730 2030 790
rect 2090 730 2100 790
rect 1670 680 2110 690
rect 1670 640 1890 680
rect 1540 630 1890 640
rect 2050 630 2110 680
rect 1540 620 2110 630
rect 1670 360 1750 370
rect 1670 300 1680 360
rect 1740 340 1750 360
rect 1740 300 2250 340
rect 1670 290 2250 300
rect 690 240 1940 260
rect 690 -110 710 240
rect 870 -110 1940 240
rect 690 -130 1940 -110
rect 1990 240 2190 250
rect 1990 -120 2100 240
rect 2180 -120 2190 240
rect 1990 -130 2190 -120
rect 1670 -180 2000 -170
rect 1670 -240 1680 -180
rect 1740 -220 2000 -180
rect 1740 -240 1750 -220
rect 1670 -250 1750 -240
rect 2230 -270 2700 -220
rect 2230 -350 2280 -270
rect 1090 -370 2280 -350
rect 1090 -460 1110 -370
rect 1270 -460 2280 -370
rect 1090 -480 2280 -460
rect 2230 -550 2280 -480
rect 2320 -320 2600 -310
rect 2320 -500 2330 -320
rect 2460 -500 2600 -320
rect 2320 -510 2600 -500
rect 1670 -590 1750 -580
rect 1670 -650 1680 -590
rect 1740 -610 1750 -590
rect 2230 -600 2700 -550
rect 1740 -650 2000 -610
rect 1670 -660 2000 -650
rect 290 -710 1940 -690
rect 290 -1060 310 -710
rect 470 -1060 1940 -710
rect 290 -1080 1940 -1060
rect 1990 -710 2190 -700
rect 1990 -1070 2100 -710
rect 2180 -1070 2190 -710
rect 1990 -1080 2190 -1070
rect 1670 -1130 2250 -1120
rect 1670 -1190 1680 -1130
rect 1740 -1170 2250 -1130
rect 1740 -1190 1750 -1170
rect 1670 -1200 1750 -1190
rect 8470 -6085 8560 2855
rect 8630 -6085 8650 2855
rect 8970 2820 9590 4020
rect 10430 4180 11050 4200
rect 10430 4020 10450 4180
rect 11030 4020 11050 4180
rect 9920 3780 10100 3800
rect 9920 3620 9940 3780
rect 10080 3620 10100 3780
rect 9920 2850 10100 3620
rect 8690 2350 9870 2820
rect 8680 -6060 9880 -5580
rect 8470 -6260 8650 -6085
rect 8970 -7490 9590 -6060
rect 9920 -6090 9940 2850
rect 10080 -6090 10100 2850
rect 10430 2820 11050 4020
rect 11370 3780 11550 3800
rect 11370 3620 11390 3780
rect 11530 3620 11550 3780
rect 11370 2855 11550 3620
rect 10150 2350 11330 2820
rect 10140 -6060 11340 -5580
rect 9920 -6260 10100 -6090
rect 10430 -7090 11050 -6060
rect 11370 -6085 11390 2855
rect 11460 -6085 11550 2855
rect 11370 -6260 11550 -6085
rect 11224 -6870 11230 -6670
rect 11430 -6870 11710 -6670
rect 10430 -7250 10450 -7090
rect 11030 -7250 11050 -7090
rect 10430 -7270 11050 -7250
rect 11224 -7270 11230 -7070
rect 11430 -7270 11710 -7070
rect 8970 -7650 8990 -7490
rect 9570 -7650 9590 -7490
rect 8970 -7670 9590 -7650
rect 11430 -7670 11710 -7470
<< via1 >>
rect 1280 5010 1340 5020
rect 1280 4960 1330 5010
rect 1330 4960 1340 5010
rect 1280 4780 1340 4790
rect 1280 4730 1330 4780
rect 1330 4730 1340 4780
rect 350 4000 550 4200
rect 860 4020 1120 4180
rect 350 3600 550 3800
rect 1560 3620 1820 3780
rect 1380 3220 1460 3350
rect 2050 3620 2340 3780
rect 1890 3230 1970 3340
rect 2420 3230 2500 3340
rect 8990 4020 9570 4180
rect 8490 3620 8630 3780
rect 2650 3070 2710 3130
rect 2800 3070 2860 3130
rect 1560 2580 1670 2690
rect 2030 2460 2090 2520
rect 710 1860 870 2400
rect 2030 1740 2090 1800
rect 1560 1570 1670 1680
rect 2030 1450 2090 1510
rect 310 850 470 1390
rect 1560 640 1670 750
rect 2030 730 2090 790
rect 1680 300 1740 360
rect 710 -110 870 240
rect 2100 -120 2180 240
rect 1680 -240 1740 -180
rect 1110 -460 1270 -370
rect 2330 -500 2460 -320
rect 1680 -650 1740 -590
rect 310 -1060 470 -710
rect 2100 -1070 2180 -710
rect 1680 -1190 1740 -1130
rect 10450 4020 11030 4180
rect 9940 3620 10080 3780
rect 11390 3620 11530 3780
rect 11230 -6870 11430 -6670
rect 10450 -7250 11030 -7090
rect 11230 -7270 11430 -7070
rect 8990 -7650 9570 -7490
rect 11230 -7670 11430 -7470
<< metal2 >>
rect 1270 5020 1350 5030
rect 1270 4960 1280 5020
rect 1340 4960 1350 5020
rect 1270 4790 1350 4960
rect 1270 4730 1280 4790
rect 1340 4730 1350 4790
rect 1270 4710 1350 4730
rect 330 4200 570 4220
rect 330 4000 350 4200
rect 550 4000 570 4200
rect 840 4180 1140 4200
rect 840 4020 860 4180
rect 1120 4020 1140 4180
rect 840 4000 1140 4020
rect 8970 4180 9590 4200
rect 8970 4020 8990 4180
rect 9570 4020 9590 4180
rect 8970 4000 9590 4020
rect 10430 4180 11050 4200
rect 10430 4020 10450 4180
rect 11030 4020 11050 4180
rect 10430 4000 11050 4020
rect 330 3980 570 4000
rect 330 3800 570 3820
rect 330 3600 350 3800
rect 550 3600 570 3800
rect 1540 3780 1840 3800
rect 1540 3620 1560 3780
rect 1820 3620 1840 3780
rect 1540 3600 1840 3620
rect 2030 3780 2360 3800
rect 2030 3620 2050 3780
rect 2340 3620 2360 3780
rect 2030 3600 2360 3620
rect 8470 3780 8650 3800
rect 8470 3620 8490 3780
rect 8630 3620 8650 3780
rect 8470 3600 8650 3620
rect 9920 3780 10100 3800
rect 9920 3620 9940 3780
rect 10080 3620 10100 3780
rect 9920 3600 10100 3620
rect 11370 3780 11550 3800
rect 11370 3620 11390 3780
rect 11530 3620 11550 3780
rect 11370 3600 11550 3620
rect 330 3580 570 3600
rect 1090 3220 1380 3350
rect 1460 3340 8390 3350
rect 1460 3230 1890 3340
rect 1970 3230 2420 3340
rect 2500 3230 8390 3340
rect 1460 3220 8390 3230
rect 690 2400 890 2420
rect 690 1860 710 2400
rect 870 1860 890 2400
rect 690 1840 890 1860
rect 290 1390 490 1410
rect 290 850 310 1390
rect 470 850 490 1390
rect 290 830 490 850
rect 690 240 890 260
rect 690 -110 710 240
rect 870 -110 890 240
rect 690 -130 890 -110
rect 1090 -370 1290 3220
rect 2650 3130 2710 3136
rect 1540 2690 1690 2710
rect 1540 2580 1560 2690
rect 1670 2580 1690 2690
rect 1540 1680 1690 2580
rect 2650 2520 2710 3070
rect 2020 2460 2030 2520
rect 2090 2460 2710 2520
rect 2800 3130 2860 3136
rect 2440 1800 2500 2460
rect 2800 2370 2860 3070
rect 2020 1740 2030 1800
rect 2090 1740 2500 1800
rect 2580 2310 2860 2370
rect 1540 1570 1560 1680
rect 1670 1570 1690 1680
rect 1540 750 1690 1570
rect 2580 1510 2640 2310
rect 2020 1450 2030 1510
rect 2090 1450 2640 1510
rect 2440 790 2500 1450
rect 1540 640 1560 750
rect 1670 640 1690 750
rect 2020 730 2030 790
rect 2090 730 2500 790
rect 1540 620 1690 640
rect 1670 360 1750 370
rect 1670 300 1680 360
rect 1740 300 1750 360
rect 1670 -180 1750 300
rect 2090 240 2470 250
rect 2090 -120 2100 240
rect 2180 -120 2470 240
rect 2090 -130 2470 -120
rect 1670 -240 1680 -180
rect 1740 -240 1750 -180
rect 1670 -250 1750 -240
rect 1090 -460 1110 -370
rect 1270 -460 1290 -370
rect 290 -710 490 -690
rect 290 -1060 310 -710
rect 470 -1060 490 -710
rect 290 -1080 490 -1060
rect 1090 -6670 1290 -460
rect 2320 -320 2470 -130
rect 2320 -500 2330 -320
rect 2460 -500 2470 -320
rect 1670 -590 1750 -580
rect 1670 -650 1680 -590
rect 1740 -650 1750 -590
rect 1670 -1130 1750 -650
rect 2320 -700 2470 -500
rect 2090 -710 2470 -700
rect 2090 -1070 2100 -710
rect 2180 -1070 2470 -710
rect 2090 -1080 2470 -1070
rect 1670 -1190 1680 -1130
rect 1740 -1190 1750 -1130
rect 1670 -1200 1750 -1190
rect 11230 -6670 11430 -6664
rect 1090 -6870 11230 -6670
rect 11230 -6876 11430 -6870
rect 11230 -7070 11430 -7064
rect 10430 -7090 11050 -7070
rect 10430 -7250 10450 -7090
rect 11030 -7250 11050 -7090
rect 10430 -7270 11050 -7250
rect 11221 -7270 11230 -7070
rect 11430 -7270 11439 -7070
rect 11230 -7276 11430 -7270
rect 8970 -7490 9590 -7470
rect 8970 -7650 8990 -7490
rect 9570 -7650 9590 -7490
rect 8970 -7670 9590 -7650
<< via2 >>
rect 350 4000 550 4200
rect 860 4020 1120 4180
rect 8990 4020 9570 4180
rect 10450 4020 11030 4180
rect 350 3600 550 3800
rect 1560 3620 1820 3780
rect 2050 3620 2340 3780
rect 8490 3620 8630 3780
rect 9940 3620 10080 3780
rect 11390 3620 11530 3780
rect 710 1860 870 2400
rect 310 850 470 1390
rect 710 -110 870 240
rect 310 -1060 470 -710
rect 10450 -7250 11030 -7090
rect 11230 -7270 11430 -7070
rect 8990 -7650 9570 -7490
rect 11230 -7670 11430 -7470
<< metal3 >>
rect 330 4205 570 4220
rect 330 3995 345 4205
rect 555 3995 570 4205
rect 840 4180 1140 4200
rect 840 4020 860 4180
rect 1120 4020 1140 4180
rect 840 4000 1140 4020
rect 8970 4180 9590 4200
rect 8970 4020 8990 4180
rect 9570 4020 9590 4180
rect 8970 4000 9590 4020
rect 10430 4180 11050 4200
rect 10430 4020 10450 4180
rect 11030 4020 11050 4180
rect 10430 4000 11050 4020
rect 330 3980 570 3995
rect 345 3800 555 3805
rect 345 3600 350 3800
rect 550 3780 11550 3800
rect 550 3620 1560 3780
rect 1820 3620 2050 3780
rect 2340 3620 8490 3780
rect 8630 3620 9940 3780
rect 10080 3620 11390 3780
rect 11530 3620 11550 3780
rect 550 3600 11550 3620
rect 345 3595 555 3600
rect 690 2400 890 2980
rect 690 1860 710 2400
rect 870 1860 890 2400
rect 290 1390 490 1410
rect 290 850 310 1390
rect 470 850 490 1390
rect 290 830 490 850
rect 690 240 890 1860
rect 690 -110 710 240
rect 870 -110 890 240
rect 290 -710 490 -690
rect 290 -1060 310 -710
rect 470 -1060 490 -710
rect 290 -1080 490 -1060
rect 690 -7070 890 -110
rect 11225 -7070 11435 -7065
rect 690 -7090 11230 -7070
rect 690 -7250 10450 -7090
rect 11030 -7250 11230 -7090
rect 690 -7270 11230 -7250
rect 11430 -7270 11435 -7070
rect 11225 -7275 11435 -7270
rect 8970 -7490 9590 -7470
rect 8970 -7650 8990 -7490
rect 9570 -7650 9590 -7490
rect 8970 -7670 9590 -7650
rect 11219 -7675 11225 -7465
rect 11425 -7470 11435 -7465
rect 11430 -7670 11435 -7470
rect 11425 -7675 11435 -7670
<< via3 >>
rect 345 4200 555 4205
rect 345 4000 350 4200
rect 350 4000 550 4200
rect 550 4000 555 4200
rect 345 3995 555 4000
rect 860 4020 1120 4180
rect 8990 4020 9570 4180
rect 10450 4020 11030 4180
rect 310 850 470 1390
rect 310 -1060 470 -710
rect 8990 -7650 9570 -7490
rect 11225 -7470 11425 -7465
rect 11225 -7670 11230 -7470
rect 11230 -7670 11425 -7470
rect 11225 -7675 11425 -7670
<< metal4 >>
rect 344 4205 556 4206
rect 344 3995 345 4205
rect 555 4200 556 4205
rect 555 4180 11550 4200
rect 555 4020 860 4180
rect 1120 4020 8990 4180
rect 9570 4020 10450 4180
rect 11030 4020 11550 4180
rect 555 4000 11550 4020
rect 555 3995 556 4000
rect 344 3994 556 3995
rect 290 1390 490 2980
rect 290 850 310 1390
rect 470 850 490 1390
rect 290 -710 490 850
rect 290 -1060 310 -710
rect 470 -1060 490 -710
rect 290 -7470 490 -1060
rect 11224 -7465 11426 -7464
rect 11224 -7470 11225 -7465
rect 290 -7490 11225 -7470
rect 290 -7650 8990 -7490
rect 9570 -7650 11225 -7490
rect 290 -7670 11225 -7650
rect 11224 -7675 11225 -7670
rect 11425 -7675 11426 -7465
rect 11224 -7676 11426 -7675
use sky130_fd_pr__nfet_01v8_ATLS57  sky130_fd_pr__nfet_01v8_ATLS57_0 csdac_nom__devices
timestamp 1723498766
transform -1 0 1971 0 -1 -890
box -211 -410 211 410
use sky130_fd_pr__nfet_01v8_HZS9GD  XMB0 csdac_nom__devices
timestamp 1723498766
transform 1 0 2778 0 1 -8278
box -1796 -260 1796 260
use sky130_fd_pr__nfet_01v8_FMHZDY  XMB1 csdac_nom__devices
timestamp 1723498766
transform 1 0 6436 0 1 -9110
box -996 -260 996 260
use sky130_fd_pr__nfet_01v8_AHZR5K  XMB2 csdac_nom__devices
timestamp 1723498766
transform 1 0 8713 0 1 -9269
box -596 -260 596 260
use sky130_fd_pr__nfet_01v8_BHEWB6  XMB3 csdac_nom__devices
timestamp 1723498766
transform 1 0 10400 0 1 -9428
box -406 -260 406 260
use sky130_fd_pr__nfet_01v8_FMMQLY  XMB4 csdac_nom__devices
timestamp 1723498766
transform 1 0 11787 0 1 -9587
box -296 -260 296 260
use sky130_fd_pr__nfet_01v8_C4RU6Y  XMB5 csdac_nom__devices
timestamp 1723498766
transform 1 0 13194 0 1 -9606
box -426 -400 426 400
use sky130_fd_pr__nfet_01v8_N5FCK4  XMB6 csdac_nom__devices
timestamp 1723498766
transform 1 0 2656 0 1 -410
box -246 -320 246 320
use sky130_fd_pr__nfet_01v8_8TEC39  XMB7 csdac_nom__devices
timestamp 1723498766
transform 0 -1 2180 1 0 2886
box -246 -420 246 420
use sky130_fd_pr__nfet_01v8_SMGLWN  XMmirror csdac_nom__devices
timestamp 1723498766
transform 1 0 1505 0 1 4867
box -246 -260 246 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMN0 csdac_nom__devices
timestamp 1723498766
transform 1 0 5282 0 1 -9057
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMN1
timestamp 1723498766
transform 1 0 7959 0 1 -9216
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMN2
timestamp 1723498766
transform 1 0 9836 0 1 -9375
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMN3
timestamp 1723498766
transform 1 0 11333 0 1 -9534
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMN4
timestamp 1723498766
transform 1 0 12610 0 1 -9693
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_648S5X  XMN5 csdac_nom__devices
timestamp 1723498766
transform 1 0 14147 0 1 -9802
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_ATLS57  XMN6
timestamp 1723498766
transform -1 0 1971 0 -1 60
box -211 -410 211 410
use sky130_fd_pr__nfet_01v8_J2SMEF  XMN7 csdac_nom__devices
timestamp 1723498766
transform 1 0 1971 0 1 2130
box -211 -510 211 510
use sky130_fd_pr__nfet_01v8_L9ESAD  XMP0
timestamp 1723498766
transform 1 0 4913 0 1 -9004
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMP1
timestamp 1723498766
transform 1 0 7590 0 1 -9163
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMP2
timestamp 1723498766
transform 1 0 9467 0 1 -9322
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMP3
timestamp 1723498766
transform 1 0 10964 0 1 -9481
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMP4
timestamp 1723498766
transform 1 0 12241 0 1 -9640
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_648S5X  XMP5
timestamp 1723498766
transform 1 0 13778 0 1 -9749
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_J2SMEF  XMP7
timestamp 1723498766
transform 1 0 1971 0 1 1120
box -211 -510 211 510
use sky130_fd_pr__pfet_01v8_XJ7GBL  XMprog csdac_nom__devices
timestamp 1723498766
transform 1 0 1031 0 1 4869
box -211 -269 211 269
use sky130_fd_pr__res_high_po_5p73_MRHKYZ  XR5 csdac_nom__devices
timestamp 1723498766
transform 1 0 9279 0 1 -1618
box -739 -4582 739 4582
use sky130_fd_pr__res_high_po_5p73_MRHKYZ  XR6
timestamp 1723498766
transform 1 0 10739 0 1 -1618
box -739 -4582 739 4582
<< labels >>
flabel metal1 7994 5696 8194 5896 0 FreeSans 256 90 0 0 p0
port 2 nsew
flabel metal1 7594 5696 7794 5896 0 FreeSans 256 90 0 0 n0
port 3 nsew
flabel metal1 7194 5696 7394 5896 0 FreeSans 256 90 0 0 p1
port 4 nsew
flabel metal1 6794 5696 6994 5896 0 FreeSans 256 90 0 0 n1
port 5 nsew
flabel metal1 6394 5696 6594 5896 0 FreeSans 256 90 0 0 p2
port 6 nsew
flabel metal1 5994 5696 6194 5896 0 FreeSans 256 90 0 0 n2
port 7 nsew
flabel metal1 5594 5696 5794 5896 0 FreeSans 256 90 0 0 p3
port 8 nsew
flabel metal1 5194 5696 5394 5896 0 FreeSans 256 90 0 0 n3
port 9 nsew
flabel metal1 4794 5696 4994 5896 0 FreeSans 256 90 0 0 p4
port 10 nsew
flabel metal1 4394 5696 4594 5896 0 FreeSans 256 90 0 0 n4
port 11 nsew
flabel metal1 3994 5696 4194 5896 0 FreeSans 256 90 0 0 p5
port 12 nsew
flabel metal1 3594 5696 3794 5896 0 FreeSans 256 90 0 0 n5
port 13 nsew
flabel metal1 3194 5696 3394 5896 0 FreeSans 256 90 0 0 p6
port 14 nsew
flabel metal1 2794 5696 2994 5896 0 FreeSans 256 90 0 0 n6
port 15 nsew
flabel metal1 2394 5696 2594 5896 0 FreeSans 256 90 0 0 p7
port 16 nsew
flabel metal1 1994 5696 2194 5896 0 FreeSans 256 90 0 0 n7
port 17 nsew
flabel metal1 0 4000 200 4200 0 FreeSans 256 0 0 0 vcc
port 0 nsew
flabel metal1 0 3600 200 3800 0 FreeSans 256 0 0 0 vss
port 1 nsew
flabel metal1 11510 -7670 11710 -7470 0 FreeSans 256 180 0 0 Vpos
port 18 nsew
flabel metal1 11510 -6870 11710 -6670 0 FreeSans 256 180 0 0 Vbias
port 20 nsew
flabel metal1 11510 -7270 11710 -7070 0 FreeSans 256 180 0 0 Vneg
port 19 nsew
flabel metal1 2170 830 2380 2830 0 FreeSans 800 0 0 0 IS7
<< end >>

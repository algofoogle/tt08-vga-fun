magic
tech sky130A
magscale 1 2
timestamp 1723412611
<< error_s >>
rect 5552 4902 5610 4908
rect 5962 4902 6020 4908
rect 5552 4868 5564 4902
rect 5962 4868 5974 4902
rect 5552 4862 5610 4868
rect 5962 4862 6020 4868
rect 5552 4692 5610 4698
rect 5962 4692 6020 4698
rect 5552 4658 5564 4692
rect 5962 4658 5974 4692
rect 5552 4652 5610 4658
rect 5962 4652 6020 4658
rect 9199 520 9234 554
rect 9200 501 9234 520
rect 9030 452 9088 458
rect 9030 418 9042 452
rect 9030 412 9088 418
rect 9030 242 9088 248
rect 9030 208 9042 242
rect 9030 202 9088 208
rect 9219 106 9234 501
rect 9253 467 9288 501
rect 9568 467 9603 501
rect 9253 106 9287 467
rect 9569 448 9603 467
rect 9399 399 9457 405
rect 9399 365 9411 399
rect 9399 359 9457 365
rect 9399 189 9457 195
rect 9399 155 9411 189
rect 9399 149 9457 155
rect 9253 72 9268 106
rect 9588 53 9603 448
rect 9622 414 9657 448
rect 10327 414 10362 448
rect 9622 53 9656 414
rect 10328 395 10362 414
rect 9622 19 9637 53
rect 10347 0 10362 395
rect 10381 361 10416 395
rect 10696 361 10731 395
rect 10381 0 10415 361
rect 10697 342 10731 361
rect 10527 293 10585 299
rect 10527 259 10539 293
rect 10527 253 10585 259
rect 10527 83 10585 89
rect 10527 49 10539 83
rect 10527 43 10585 49
rect 10381 -34 10396 0
rect 10716 -53 10731 342
rect 10750 308 10785 342
rect 11065 308 11100 342
rect 10750 -53 10784 308
rect 11066 289 11100 308
rect 10896 240 10954 246
rect 10896 206 10908 240
rect 10896 200 10954 206
rect 10896 30 10954 36
rect 10896 -4 10908 30
rect 10896 -10 10954 -4
rect 10750 -87 10765 -53
rect 11085 -106 11100 289
rect 11119 255 11154 289
rect 11604 255 11639 289
rect 11119 -106 11153 255
rect 11605 236 11639 255
rect 11119 -140 11134 -106
rect 11624 -159 11639 236
rect 11658 202 11693 236
rect 11973 202 12008 236
rect 11658 -159 11692 202
rect 11974 183 12008 202
rect 11804 134 11862 140
rect 11804 100 11816 134
rect 11804 94 11862 100
rect 11804 -76 11862 -70
rect 11804 -110 11816 -76
rect 11804 -116 11862 -110
rect 11658 -193 11673 -159
rect 11993 -212 12008 183
rect 12027 149 12062 183
rect 12027 -212 12061 149
rect 12173 81 12231 87
rect 12173 47 12185 81
rect 12173 41 12231 47
rect 12173 -129 12231 -123
rect 12173 -163 12185 -129
rect 12173 -169 12231 -163
rect 12027 -246 12042 -212
rect 12362 -265 12377 183
rect 12396 -265 12430 237
rect 13142 177 13176 231
rect 15864 225 15899 259
rect 14687 184 14722 218
rect 15865 206 15899 225
rect 12396 -299 12411 -265
rect 13161 -318 13176 177
rect 13195 143 13230 177
rect 13510 143 13545 177
rect 14688 165 14722 184
rect 13195 -318 13229 143
rect 13511 124 13545 143
rect 13341 75 13399 81
rect 13341 41 13353 75
rect 13341 35 13399 41
rect 13341 -235 13399 -229
rect 13341 -269 13353 -235
rect 13341 -275 13399 -269
rect 13195 -352 13210 -318
rect 13530 -371 13545 124
rect 13564 90 13599 124
rect 13879 91 13914 124
rect 13564 -371 13598 90
rect 13710 22 13768 28
rect 13710 -12 13722 22
rect 13710 -18 13768 -12
rect 13710 -288 13768 -282
rect 13710 -322 13722 -288
rect 13710 -328 13768 -322
rect 13564 -405 13579 -371
rect 13899 -424 13914 91
rect 13933 57 13968 91
rect 13933 -424 13967 57
rect 13933 -458 13948 -424
rect 14338 -477 14353 91
rect 14372 -477 14406 145
rect 14518 116 14576 122
rect 14518 82 14530 116
rect 14518 76 14576 82
rect 14518 -394 14576 -388
rect 14518 -428 14530 -394
rect 14518 -434 14576 -428
rect 14372 -511 14387 -477
rect 14707 -530 14722 165
rect 14741 131 14776 165
rect 15056 132 15091 165
rect 14741 -530 14775 131
rect 14887 63 14945 69
rect 14887 29 14899 63
rect 14887 23 14945 29
rect 14887 -447 14945 -441
rect 14887 -481 14899 -447
rect 14887 -487 14945 -481
rect 14741 -564 14756 -530
rect 15076 -583 15091 132
rect 15110 98 15145 132
rect 15110 -583 15144 98
rect 15110 -617 15125 -583
rect 15515 -636 15530 132
rect 15549 -636 15583 186
rect 15695 157 15753 163
rect 15695 123 15707 157
rect 15695 117 15753 123
rect 15695 -553 15753 -547
rect 15695 -587 15707 -553
rect 15695 -593 15753 -587
rect 15549 -670 15564 -636
rect 15884 -689 15899 206
rect 15918 172 15953 206
rect 15918 -689 15952 172
rect 16064 104 16122 110
rect 16064 70 16076 104
rect 16064 64 16122 70
rect 16064 -606 16122 -600
rect 16064 -640 16076 -606
rect 16064 -646 16122 -640
rect 15918 -723 15933 -689
<< viali >>
rect 7360 6170 7610 6220
rect 7890 6180 8060 6230
rect 7270 5850 7320 6130
rect 7650 6070 7710 6120
rect 7650 5860 7710 5910
rect 8100 5840 8160 6140
rect 7360 5760 7410 5810
rect 7560 5760 7610 5810
rect 7890 5750 8060 5800
rect 6130 5340 6180 5620
rect 6850 5340 6900 5620
rect 6220 5250 6400 5300
rect 6640 5250 6820 5300
rect 6390 1570 6440 4930
rect 6800 1570 6850 4820
rect 6470 1490 6770 1540
<< metal1 >>
rect 592 7110 792 7310
rect 992 7110 1192 7310
rect 1392 7110 1592 7310
rect 1792 7110 1992 7310
rect 2192 7110 2392 7310
rect 2592 7110 2792 7310
rect 2992 7110 3192 7310
rect 3392 7110 3592 7310
rect 3792 7110 3992 7310
rect 4192 7110 4392 7310
rect 4592 7110 4792 7310
rect 4992 7110 5192 7310
rect 5392 7110 5592 7310
rect 5792 7110 5992 7310
rect 6192 7110 6392 7310
rect 6592 7110 6792 7310
rect 6120 5620 6190 5640
rect 6280 5620 6340 7110
rect 6690 5620 6750 7110
rect 7392 6335 7592 7310
rect 7874 7308 8072 7310
rect 7872 7110 8072 7308
rect 7235 6230 7592 6335
rect 7874 6270 8072 7110
rect 7860 6240 8080 6270
rect 7860 6230 8170 6240
rect 7235 6220 7720 6230
rect 7235 6170 7360 6220
rect 7610 6170 7720 6220
rect 7860 6180 7890 6230
rect 8060 6180 8170 6230
rect 7860 6170 8170 6180
rect 7235 6160 7720 6170
rect 7235 6130 7345 6160
rect 7640 6130 7720 6160
rect 8090 6140 8170 6170
rect 7235 5850 7270 6130
rect 7320 5850 7345 6130
rect 7430 6070 7600 6130
rect 7540 6020 7600 6070
rect 7640 6120 8010 6130
rect 7640 6070 7650 6120
rect 7710 6080 8010 6120
rect 7710 6070 7720 6080
rect 7640 6050 7720 6070
rect 7900 6020 7950 6050
rect 8090 6040 8100 6140
rect 7540 5960 7950 6020
rect 7540 5910 7600 5960
rect 7900 5930 7950 5960
rect 7990 5940 8100 6040
rect 7430 5850 7600 5910
rect 7640 5910 7720 5930
rect 7640 5860 7650 5910
rect 7710 5900 7720 5910
rect 7710 5860 8010 5900
rect 7640 5850 8010 5860
rect 7235 5820 7345 5850
rect 7235 5810 7430 5820
rect 7235 5760 7360 5810
rect 7410 5760 7430 5810
rect 7235 5750 7430 5760
rect 6840 5620 6910 5640
rect 6120 5340 6130 5620
rect 6180 5340 6190 5620
rect 6270 5560 6370 5620
rect 6430 5560 6440 5620
rect 6590 5560 6600 5620
rect 6660 5560 6760 5620
rect 6330 5430 6700 5530
rect 6270 5340 6370 5400
rect 6430 5340 6440 5400
rect 6120 5310 6190 5340
rect 6120 5300 6450 5310
rect 6120 5250 6220 5300
rect 6400 5250 6450 5300
rect 6120 5240 6450 5250
rect 6380 5175 6450 5240
rect 6380 4930 6450 5105
rect 6380 1570 6390 4930
rect 6440 1570 6450 4930
rect 6490 1635 6540 5430
rect 6590 5340 6600 5400
rect 6660 5340 6760 5400
rect 6840 5340 6850 5620
rect 6900 5340 6910 5620
rect 6840 5310 6910 5340
rect 6620 5300 6910 5310
rect 6620 5250 6640 5300
rect 6820 5250 6910 5300
rect 6620 5240 6910 5250
rect 6840 5190 6910 5240
rect 7235 5190 7345 5750
rect 6820 5170 7345 5190
rect 6820 5110 6840 5170
rect 6910 5110 7345 5170
rect 6820 5080 7345 5110
rect 7460 4950 7510 5850
rect 7640 5820 7720 5850
rect 7540 5810 7720 5820
rect 8090 5840 8100 5940
rect 8160 5840 8170 6140
rect 8090 5810 8170 5840
rect 7540 5760 7560 5810
rect 7610 5760 7720 5810
rect 7540 5750 7720 5760
rect 7870 5800 8170 5810
rect 7870 5750 7890 5800
rect 8060 5750 8170 5800
rect 7870 5740 8170 5750
rect 6570 4900 7515 4950
rect 6570 1600 6670 4900
rect 6700 4820 6860 4850
rect 6700 1670 6800 4820
rect 6380 1560 6450 1570
rect 6790 1570 6800 1670
rect 6850 4805 6860 4820
rect 6850 4735 6995 4805
rect 7065 4735 7071 4805
rect 6850 1570 6860 4735
rect 6790 1560 6860 1570
rect 6380 1540 6860 1560
rect 6380 1490 6470 1540
rect 6770 1490 6860 1540
rect 6380 1480 6860 1490
rect 7465 -5385 7515 4900
rect 7015 -5435 7515 -5385
rect 7015 -7482 7065 -5435
rect 6940 -7682 7140 -7482
rect 7340 -7682 7540 -7482
rect 7740 -7682 7940 -7482
<< via1 >>
rect 6370 5560 6430 5620
rect 6600 5560 6660 5620
rect 6370 5340 6430 5400
rect 6380 5105 6450 5175
rect 6600 5340 6660 5400
rect 6840 5110 6910 5170
rect 6995 4735 7065 4805
<< metal2 >>
rect 6360 5620 6440 5630
rect 6360 5560 6370 5620
rect 6430 5560 6440 5620
rect 6360 5400 6440 5560
rect 6360 5340 6370 5400
rect 6430 5340 6440 5400
rect 6360 5330 6440 5340
rect 6590 5620 6670 5630
rect 6590 5560 6600 5620
rect 6660 5560 6670 5620
rect 6590 5400 6670 5560
rect 6590 5340 6600 5400
rect 6660 5340 6670 5400
rect 6590 5330 6670 5340
rect 6370 5175 6460 5180
rect 6370 5105 6380 5175
rect 6450 5170 7065 5175
rect 6450 5110 6840 5170
rect 6910 5110 7065 5170
rect 6450 5105 7065 5110
rect 6370 5100 6460 5105
rect 6995 4805 7065 5105
rect 6995 4729 7065 4735
use sky130_fd_pr__nfet_01v8_HZS9GD  XMB0 csdac_nom__devices
timestamp 1723353804
transform 0 1 6620 -1 0 3256
box -1796 -260 1796 260
use sky130_fd_pr__nfet_01v8_FMHZDY  XMB1 csdac_nom__devices
timestamp 1723353804
transform 0 1 5900 -1 0 3266
box -996 -260 996 260
use sky130_fd_pr__nfet_01v8_AHZR5K  XMB2 csdac_nom__devices
timestamp 1723353804
transform 1 0 3256 0 1 2820
box -596 -260 596 260
use sky130_fd_pr__nfet_01v8_BHEWB6  XMB3 csdac_nom__devices
timestamp 1723353804
transform 1 0 9992 0 1 224
box -406 -260 406 260
use sky130_fd_pr__nfet_01v8_FMMQLY  XMB4 csdac_nom__devices
timestamp 1723353804
transform 1 0 11379 0 1 65
box -296 -260 296 260
use sky130_fd_pr__nfet_01v8_C4RU6Y  XMB5 csdac_nom__devices
timestamp 1723353804
transform 1 0 12786 0 1 46
box -426 -400 426 400
use sky130_fd_pr__nfet_01v8_N5FCK4  XMB6 csdac_nom__devices
timestamp 1723353804
transform 1 0 14143 0 1 -193
box -246 -320 246 320
use sky130_fd_pr__nfet_01v8_8TEC39  XMB7 csdac_nom__devices
timestamp 1723353804
transform 1 0 15320 0 1 -252
box -246 -420 246 420
use sky130_fd_pr__nfet_01v8_SMGLWN  XMmirror csdac_nom__devices
timestamp 1723353804
transform 1 0 7486 0 1 5990
box -246 -260 246 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMN0 csdac_nom__devices
timestamp 1723353804
transform 1 0 6311 0 1 5480
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMN1
timestamp 1723353804
transform 1 0 5581 0 1 4780
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMN2
timestamp 1723353804
transform 1 0 9428 0 1 277
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMN3
timestamp 1723353804
transform 1 0 10925 0 1 118
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMN4
timestamp 1723353804
transform 1 0 12202 0 1 -41
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_648S5X  XMN5 csdac_nom__devices
timestamp 1723353804
transform 1 0 13739 0 1 -150
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_ATLS57  XMN6 csdac_nom__devices
timestamp 1723353804
transform 1 0 14916 0 1 -209
box -211 -410 211 410
use sky130_fd_pr__nfet_01v8_J2SMEF  XMN7 csdac_nom__devices
timestamp 1723353804
transform 1 0 16093 0 1 -268
box -211 -510 211 510
use sky130_fd_pr__nfet_01v8_L9ESAD  XMP0
timestamp 1723353804
transform 1 0 6721 0 1 5480
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMP1
timestamp 1723353804
transform 1 0 5991 0 1 4780
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMP2
timestamp 1723353804
transform 1 0 9059 0 1 330
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMP3
timestamp 1723353804
transform 1 0 10556 0 1 171
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMP4
timestamp 1723353804
transform 1 0 11833 0 1 12
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_648S5X  XMP5
timestamp 1723353804
transform 1 0 13370 0 1 -97
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_ATLS57  XMP6
timestamp 1723353804
transform 1 0 14547 0 1 -156
box -211 -410 211 410
use sky130_fd_pr__nfet_01v8_J2SMEF  XMP7
timestamp 1723353804
transform 1 0 15724 0 1 -215
box -211 -510 211 510
use sky130_fd_pr__pfet_01v8_XJ7GBL  XMprog csdac_nom__devices
timestamp 1723353804
transform 1 0 7971 0 1 5989
box -211 -269 211 269
use sky130_fd_pr__res_high_po_5p73_MRHKYZ  XR5 csdac_nom__devices
timestamp 1723353804
transform 1 0 14129 0 1 7402
box -739 -4582 739 4582
use sky130_fd_pr__res_high_po_5p73_MRHKYZ  XR6
timestamp 1723353804
transform 1 0 18415 0 1 3698
box -739 -4582 739 4582
<< labels >>
flabel metal1 7740 -7682 7940 -7482 0 FreeSans 256 90 0 0 Vpos
port 18 nsew
flabel metal1 7340 -7682 7540 -7482 0 FreeSans 256 90 0 0 Vneg
port 19 nsew
flabel metal1 6940 -7682 7140 -7482 0 FreeSans 256 90 0 0 Vbias
port 20 nsew
flabel metal1 6592 7110 6792 7310 0 FreeSans 256 90 0 0 p0
port 2 nsew
flabel metal1 6192 7110 6392 7310 0 FreeSans 256 90 0 0 n0
port 3 nsew
flabel metal1 5792 7110 5992 7310 0 FreeSans 256 90 0 0 p1
port 4 nsew
flabel metal1 5392 7110 5592 7310 0 FreeSans 256 90 0 0 n1
port 5 nsew
flabel metal1 4992 7110 5192 7310 0 FreeSans 256 90 0 0 p2
port 6 nsew
flabel metal1 4592 7110 4792 7310 0 FreeSans 256 90 0 0 n2
port 7 nsew
flabel metal1 4192 7110 4392 7310 0 FreeSans 256 90 0 0 p3
port 8 nsew
flabel metal1 3792 7110 3992 7310 0 FreeSans 256 90 0 0 n3
port 9 nsew
flabel metal1 3392 7110 3592 7310 0 FreeSans 256 90 0 0 p4
port 10 nsew
flabel metal1 2992 7110 3192 7310 0 FreeSans 256 90 0 0 n4
port 11 nsew
flabel metal1 2592 7110 2792 7310 0 FreeSans 256 90 0 0 p5
port 12 nsew
flabel metal1 2192 7110 2392 7310 0 FreeSans 256 90 0 0 n5
port 13 nsew
flabel metal1 1792 7110 1992 7310 0 FreeSans 256 90 0 0 p6
port 14 nsew
flabel metal1 1392 7110 1592 7310 0 FreeSans 256 90 0 0 n6
port 15 nsew
flabel metal1 992 7110 1192 7310 0 FreeSans 256 90 0 0 p7
port 16 nsew
flabel metal1 592 7110 792 7310 0 FreeSans 256 90 0 0 n7
port 17 nsew
flabel metal1 7392 7110 7592 7310 0 FreeSans 256 90 0 0 vss
port 1 nsew
flabel space 7872 7110 8072 7310 0 FreeSans 256 90 0 0 vcc
port 0 nsew
flabel metal1 6490 5190 6540 5250 0 FreeSans 320 0 0 0 IS0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1723783876
<< pwell >>
rect 6700 1410 6780 1450
rect 6900 1420 7000 1470
rect 1680 -1880 1740 -1820
rect 1540 -2260 1630 -2170
rect 1550 -2830 1620 -2670
rect 1920 -2960 2010 -2890
rect 1920 -3190 2010 -3120
rect 1550 -3280 1620 -3210
rect 1550 -3510 1620 -3440
rect 2290 -3720 2370 -3640
rect 1550 -4000 1620 -3850
rect 1550 -4440 1620 -4370
rect 1550 -4670 1620 -4600
rect 1550 -5100 1620 -5030
<< viali >>
rect 940 4860 1120 4910
rect 1380 4850 1630 4900
rect 850 4520 900 4810
rect 1280 4760 1330 4810
rect 1280 4530 1330 4580
rect 1680 4530 1720 4800
rect 940 4430 1120 4480
rect 1510 4440 1630 4480
rect 2040 3050 2350 3100
rect 1790 2760 1840 3010
rect 1890 2570 2090 2710
rect 6210 2380 6390 2430
rect 6820 2390 7080 2430
rect 6210 1970 6390 2020
rect 6220 1710 6380 1760
rect 1890 1560 2050 1690
rect 6720 1390 6760 1440
rect 7130 1390 7180 2340
rect 6220 1300 6380 1350
rect 6820 1300 7080 1340
rect 6260 850 6420 900
rect 7080 860 7200 910
rect 1890 630 2050 680
rect 1890 390 2060 450
rect 6260 440 6420 490
rect 6260 50 6420 100
rect 2540 -170 2780 -120
rect 1890 -320 2060 -280
rect 1890 -550 2060 -510
rect 2820 -610 2880 -210
rect 6260 -360 6420 -310
rect 2540 -700 2780 -650
rect 6830 -930 6880 -260
rect 7240 -930 7300 800
rect 6930 -1030 7190 -980
rect 1890 -1280 2060 -1220
rect 1800 -1450 1970 -1400
rect 6260 -1510 6420 -1460
rect 6950 -1500 7190 -1460
rect 2370 -1740 2980 -1690
rect 1800 -1970 1970 -1920
rect 1800 -2230 1970 -2180
rect 3010 -2350 3070 -1770
rect 6260 -1920 6420 -1870
rect 6260 -2310 6420 -2260
rect 2370 -2430 2980 -2380
rect 1800 -2740 1970 -2690
rect 6260 -2720 6420 -2670
rect 2070 -2850 2230 -2810
rect 2800 -3180 2980 -3130
rect 2070 -3270 2230 -3230
rect 2070 -3490 2230 -3450
rect 3020 -3500 3080 -3220
rect 2800 -3590 2980 -3540
rect 2070 -3910 2230 -3870
rect 1870 -4000 2030 -3960
rect 2460 -4340 3020 -4280
rect 1870 -4420 2030 -4380
rect 1870 -4660 2030 -4620
rect 3060 -4660 3120 -4380
rect 2460 -4760 3020 -4700
rect 6820 -4900 6880 -2620
rect 7240 -4900 7300 -1550
rect 8240 -4970 8310 3980
rect 9610 -4970 9770 3970
rect 11060 -4970 11150 3980
rect 1870 -5080 2030 -5040
<< metal1 >>
rect 1994 5256 2194 5456
rect 2394 5256 2594 5456
rect 2794 5256 2994 5456
rect 3194 5256 3394 5456
rect 3594 5256 3794 5456
rect 3994 5256 4194 5456
rect 4394 5256 4594 5456
rect 4794 5256 4994 5456
rect 5194 5256 5394 5456
rect 5594 5256 5794 5456
rect 5994 5256 6194 5456
rect 6394 5256 6594 5456
rect 6794 5256 6994 5456
rect 7194 5256 7394 5456
rect 7594 5256 7794 5456
rect 7994 5256 8194 5456
rect 840 4910 1140 4920
rect 840 4860 940 4910
rect 1120 4860 1140 4910
rect 840 4850 1140 4860
rect 1270 4900 1730 4910
rect 1270 4850 1380 4900
rect 1630 4850 1730 4900
rect 840 4810 910 4850
rect 1270 4840 1730 4850
rect 1270 4820 1350 4840
rect 840 4520 850 4810
rect 900 4720 910 4810
rect 990 4760 1280 4820
rect 1340 4760 1350 4820
rect 1670 4800 1730 4840
rect 990 4750 1350 4760
rect 1380 4750 1560 4800
rect 1380 4720 1460 4750
rect 1670 4720 1680 4800
rect 900 4620 1010 4720
rect 1050 4620 1460 4720
rect 1560 4620 1680 4720
rect 900 4520 910 4620
rect 990 4530 1280 4590
rect 1340 4530 1350 4590
rect 990 4520 1350 4530
rect 1380 4580 1460 4620
rect 1380 4530 1560 4580
rect 1670 4530 1680 4620
rect 1720 4530 1730 4800
rect 2060 4850 2120 5256
rect 2460 5000 2520 5256
rect 2865 5155 2915 5256
rect 2865 5105 3015 5155
rect 2460 4940 2860 5000
rect 2060 4790 2710 4850
rect 840 4490 910 4520
rect 840 4480 1140 4490
rect 840 4430 940 4480
rect 1120 4430 1140 4480
rect 840 4180 1140 4430
rect 840 4020 860 4180
rect 1120 4020 1140 4180
rect 840 4000 1140 4020
rect 1380 3370 1460 4530
rect 1670 4490 1730 4530
rect 1490 4480 1730 4490
rect 1490 4440 1510 4480
rect 1630 4440 1730 4480
rect 1490 4430 1730 4440
rect 1540 3800 1730 4430
rect 1540 3780 1850 3800
rect 1540 3620 1560 3780
rect 1820 3620 1850 3780
rect 1360 3350 1480 3370
rect 1360 3220 1380 3350
rect 1460 3220 1480 3350
rect 1360 3200 1480 3220
rect 1540 3010 1850 3620
rect 2030 3780 2360 3800
rect 2030 3620 2050 3780
rect 2340 3620 2360 3780
rect 1880 3340 1980 3350
rect 1880 3230 1890 3340
rect 1970 3230 1980 3340
rect 1880 3220 1980 3230
rect 1540 2760 1790 3010
rect 1840 2760 1850 3010
rect 1890 2830 1940 3220
rect 2030 3100 2360 3620
rect 2410 3340 2510 3350
rect 2410 3230 2420 3340
rect 2500 3230 2510 3340
rect 2410 3220 2510 3230
rect 2030 3050 2040 3100
rect 2350 3050 2360 3100
rect 2030 3000 2360 3050
rect 1970 2940 2390 3000
rect 2420 2830 2470 3220
rect 2650 3130 2710 4790
rect 2800 3130 2860 4940
rect 2965 3130 3015 5105
rect 3265 3130 3315 5256
rect 3675 5155 3725 5256
rect 3455 5105 3725 5155
rect 2644 3070 2650 3130
rect 2710 3070 2716 3130
rect 2794 3070 2800 3130
rect 2860 3070 2866 3130
rect 2950 3126 3030 3130
rect 2950 3074 2964 3126
rect 3016 3074 3030 3126
rect 2950 3070 3030 3074
rect 3250 3126 3330 3130
rect 3455 3126 3505 5105
rect 4075 4995 4125 5256
rect 3625 4945 4125 4995
rect 3625 3126 3675 4945
rect 4475 4835 4525 5256
rect 3785 4785 4525 4835
rect 3785 3126 3835 4785
rect 4875 4655 4925 5256
rect 3945 4605 4925 4655
rect 3945 3126 3995 4605
rect 5265 4495 5315 5256
rect 4085 4445 5315 4495
rect 4085 3126 4135 4445
rect 5665 4335 5715 5256
rect 4235 4285 5715 4335
rect 4235 3126 4285 4285
rect 6065 3595 6115 5256
rect 5005 3545 6115 3595
rect 3250 3074 3264 3126
rect 3316 3074 3330 3126
rect 3448 3074 3454 3126
rect 3506 3074 3512 3126
rect 3618 3074 3624 3126
rect 3676 3074 3682 3126
rect 3778 3074 3784 3126
rect 3836 3074 3842 3126
rect 3938 3074 3944 3126
rect 3996 3074 4002 3126
rect 4078 3074 4084 3126
rect 4136 3074 4142 3126
rect 4228 3074 4234 3126
rect 4286 3074 4292 3126
rect 3250 3070 3330 3074
rect 1970 2770 2390 2830
rect 1540 2730 1850 2760
rect 1540 2710 2110 2730
rect 1540 2690 1890 2710
rect 1540 2580 1560 2690
rect 1670 2580 1890 2690
rect 1540 2570 1890 2580
rect 2090 2570 2110 2710
rect 1540 2560 2110 2570
rect 1930 2460 2030 2520
rect 2090 2460 2100 2520
rect 2170 2420 2380 2770
rect 690 2400 1950 2420
rect 690 1860 710 2400
rect 870 1860 1950 2400
rect 690 1840 1950 1860
rect 1990 1840 2380 2420
rect 5005 2330 5055 3545
rect 6465 3435 6515 5256
rect 6860 4300 6920 5256
rect 7260 4460 7320 5256
rect 7668 5140 7728 5256
rect 8056 5140 8116 5256
rect 7668 5080 7808 5140
rect 7260 4400 7400 4460
rect 6860 4240 7260 4300
rect 5145 3385 6515 3435
rect 5145 2446 5195 3385
rect 7200 3130 7260 4240
rect 7340 3130 7400 4400
rect 7194 3070 7200 3130
rect 7260 3070 7266 3130
rect 7334 3070 7340 3130
rect 7400 3070 7406 3130
rect 7748 3128 7808 5080
rect 7886 5080 8116 5140
rect 7886 3128 7946 5080
rect 8650 4980 9270 5000
rect 8650 4820 8670 4980
rect 9250 4820 9270 4980
rect 8150 4580 8330 4600
rect 8150 4420 8170 4580
rect 8310 4420 8330 4580
rect 8150 3980 8330 4420
rect 7742 3068 7748 3128
rect 7808 3068 7814 3128
rect 7880 3068 7886 3128
rect 7946 3068 7952 3128
rect 5138 2394 5144 2446
rect 5196 2394 5202 2446
rect 5820 2440 6410 2450
rect 5820 2370 5830 2440
rect 5950 2430 6410 2440
rect 5950 2380 6210 2430
rect 6390 2380 6410 2430
rect 6800 2430 7670 2450
rect 5950 2370 6410 2380
rect 5820 2360 6410 2370
rect 6650 2390 6750 2400
rect 5005 2280 6600 2330
rect 6650 2310 6660 2390
rect 6740 2350 6750 2390
rect 6800 2390 6820 2430
rect 7080 2390 7490 2430
rect 6800 2380 7490 2390
rect 6740 2310 7000 2350
rect 6650 2300 7000 2310
rect 4730 2240 6280 2250
rect 4730 2160 4740 2240
rect 4920 2160 6280 2240
rect 4730 2150 6280 2160
rect 6320 2240 6510 2250
rect 6320 2160 6430 2240
rect 6500 2160 6510 2240
rect 6320 2150 6510 2160
rect 6550 2120 6600 2280
rect 6900 2270 7000 2300
rect 7120 2340 7490 2380
rect 5144 2096 5196 2102
rect 6260 2070 6600 2120
rect 5144 2038 5196 2044
rect 1930 1740 2030 1800
rect 2090 1740 2100 1800
rect 1540 1690 2110 1700
rect 1540 1680 1890 1690
rect 1540 1570 1560 1680
rect 1670 1570 1890 1680
rect 1540 1560 1890 1570
rect 2050 1560 2110 1690
rect 1540 1550 2110 1560
rect 1930 1450 2030 1510
rect 2090 1450 2100 1510
rect 2170 1410 2380 1840
rect 5145 1660 5195 2038
rect 5820 2030 6410 2040
rect 5820 1960 5830 2030
rect 5950 2020 6410 2030
rect 5950 1970 6210 2020
rect 6390 1970 6410 2020
rect 5950 1960 6410 1970
rect 5820 1950 6410 1960
rect 5460 1900 7085 1910
rect 5460 1830 5470 1900
rect 5650 1830 7085 1900
rect 5460 1820 7085 1830
rect 5820 1770 6410 1780
rect 5820 1700 5830 1770
rect 5950 1760 6410 1770
rect 5950 1710 6220 1760
rect 6380 1710 6410 1760
rect 5950 1700 6410 1710
rect 5820 1690 6410 1700
rect 5145 1610 6600 1660
rect 5090 1510 6280 1580
rect 5090 1430 5110 1510
rect 5270 1480 6280 1510
rect 6320 1570 6510 1580
rect 6320 1490 6430 1570
rect 6500 1490 6510 1570
rect 6320 1480 6510 1490
rect 5270 1430 5360 1480
rect 6550 1450 6600 1610
rect 5090 1410 5360 1430
rect 290 1390 1950 1410
rect 290 850 310 1390
rect 470 850 1950 1390
rect 290 830 1950 850
rect 1990 830 2380 1410
rect 6260 1400 6600 1450
rect 6700 1440 6780 1450
rect 6700 1390 6720 1440
rect 6760 1430 6780 1440
rect 6900 1430 7000 1470
rect 7120 1430 7130 2340
rect 6760 1390 7130 1430
rect 7180 1390 7490 2340
rect 5820 1360 6410 1370
rect 5820 1290 5830 1360
rect 5950 1350 6410 1360
rect 5950 1300 6220 1350
rect 6380 1300 6410 1350
rect 5950 1290 6410 1300
rect 5820 1280 6410 1290
rect 6700 1340 7490 1390
rect 6700 1300 6820 1340
rect 7080 1300 7490 1340
rect 7650 1300 7670 2430
rect 6700 1280 7670 1300
rect 5820 910 6440 920
rect 5820 850 5830 910
rect 5950 900 6440 910
rect 5950 850 6260 900
rect 6420 850 6440 900
rect 7060 910 7670 930
rect 5820 840 6440 850
rect 6910 860 7030 870
rect 6540 810 6620 820
rect 6540 800 6550 810
rect 1540 750 1690 770
rect 1540 640 1560 750
rect 1670 690 1690 750
rect 1930 730 2030 790
rect 2090 730 2100 790
rect 6310 750 6550 800
rect 6610 750 6620 810
rect 6910 780 6920 860
rect 7000 820 7030 860
rect 7060 860 7080 910
rect 7200 860 7490 910
rect 7060 850 7490 860
rect 7000 780 7110 820
rect 6910 770 7110 780
rect 6540 740 6620 750
rect 7010 740 7110 770
rect 7230 800 7490 850
rect 4730 710 4930 730
rect 1670 680 2110 690
rect 1670 640 1890 680
rect 1540 630 1890 640
rect 2050 630 2110 680
rect 1540 620 2110 630
rect 4730 630 4750 710
rect 4910 630 6320 710
rect 6360 700 6900 710
rect 6360 640 6810 700
rect 6890 640 6900 700
rect 6360 630 6900 640
rect 4730 610 4930 630
rect 6540 590 6620 600
rect 6310 540 6550 590
rect 6540 530 6550 540
rect 6610 530 6620 590
rect 6540 520 6620 530
rect 5820 490 6440 500
rect 1540 460 3150 470
rect 1540 390 1550 460
rect 1620 450 3150 460
rect 1620 400 1890 450
rect 1620 390 1630 400
rect 1540 380 1630 390
rect 1870 390 1890 400
rect 2060 440 3150 450
rect 2060 390 2970 440
rect 1870 380 2970 390
rect 2950 370 2970 380
rect 3130 370 3150 440
rect 5820 430 5830 490
rect 5950 440 6260 490
rect 6420 440 6440 490
rect 5950 430 6440 440
rect 5820 420 6440 430
rect 1670 360 1750 370
rect 1670 300 1680 360
rect 1740 340 1750 360
rect 2950 350 3150 370
rect 2593 340 2599 341
rect 1740 300 2599 340
rect 1670 290 2599 300
rect 2593 289 2599 290
rect 2651 289 2657 341
rect 5460 320 7200 330
rect 690 240 1940 260
rect 690 -110 710 240
rect 870 -110 1940 240
rect 690 -130 1940 -110
rect 1990 240 2190 250
rect 1990 -120 2100 240
rect 2180 -120 2190 240
rect 5460 230 5470 320
rect 5650 230 7200 320
rect 5460 220 7200 230
rect 5820 110 6440 120
rect 5820 50 5830 110
rect 5950 100 6440 110
rect 5950 50 6260 100
rect 6420 50 6440 100
rect 5820 40 6440 50
rect 6540 10 6620 20
rect 6540 0 6550 10
rect 6310 -50 6550 0
rect 6610 -50 6620 10
rect 6540 -60 6620 -50
rect 5090 -90 5290 -70
rect 1990 -130 2190 -120
rect 2520 -110 3150 -90
rect 2520 -120 2970 -110
rect 2520 -170 2540 -120
rect 2780 -170 2970 -120
rect 1670 -180 2000 -170
rect 2520 -180 2970 -170
rect 1670 -240 1680 -180
rect 1740 -220 2000 -180
rect 2800 -210 2970 -180
rect 1740 -240 1750 -220
rect 1670 -250 1750 -240
rect 1540 -260 1620 -250
rect 1540 -320 1550 -260
rect 1610 -290 1620 -260
rect 2230 -270 2700 -220
rect 1870 -280 2080 -270
rect 1870 -290 1890 -280
rect 1610 -320 1890 -290
rect 2060 -320 2080 -280
rect 1540 -330 2080 -320
rect 1090 -370 1290 -350
rect 2230 -370 2280 -270
rect 2800 -300 2820 -210
rect 1090 -460 1110 -370
rect 1270 -460 2280 -370
rect 1090 -480 1290 -460
rect 1540 -510 2080 -500
rect 1540 -570 1550 -510
rect 1610 -540 1890 -510
rect 1610 -570 1620 -540
rect 1870 -550 1890 -540
rect 2060 -550 2080 -510
rect 1870 -560 2080 -550
rect 2230 -550 2280 -460
rect 2320 -320 2600 -310
rect 2320 -500 2330 -320
rect 2460 -500 2600 -320
rect 2320 -510 2600 -500
rect 2710 -520 2820 -300
rect 1540 -580 1620 -570
rect 1670 -590 1750 -580
rect 1670 -650 1680 -590
rect 1740 -610 1750 -590
rect 2230 -600 2700 -550
rect 2800 -610 2820 -520
rect 2880 -610 2970 -210
rect 1740 -650 2000 -610
rect 2800 -640 2970 -610
rect 1670 -660 2000 -650
rect 2520 -650 2970 -640
rect 290 -710 1940 -690
rect 2520 -700 2540 -650
rect 2780 -700 2970 -650
rect 290 -1060 310 -710
rect 470 -1060 1940 -710
rect 290 -1080 1940 -1060
rect 1990 -710 2190 -700
rect 1990 -1070 2100 -710
rect 2180 -1070 2190 -710
rect 2520 -710 2970 -700
rect 3130 -710 3150 -110
rect 5090 -170 5110 -90
rect 5270 -170 6320 -90
rect 6360 -100 6900 -90
rect 6360 -160 6810 -100
rect 6890 -160 6900 -100
rect 6360 -170 6900 -160
rect 5090 -190 5290 -170
rect 6540 -210 6620 -200
rect 6310 -260 6550 -210
rect 6540 -270 6550 -260
rect 6610 -270 6620 -210
rect 6540 -280 6620 -270
rect 6810 -260 6900 -230
rect 5820 -310 6440 -300
rect 5820 -370 5830 -310
rect 5950 -360 6260 -310
rect 6420 -360 6440 -310
rect 5950 -370 6440 -360
rect 5820 -380 6440 -370
rect 2520 -730 3150 -710
rect 6810 -930 6830 -260
rect 6880 -900 6900 -260
rect 7010 -900 7110 -870
rect 7230 -900 7240 800
rect 6880 -930 7240 -900
rect 7300 -930 7490 800
rect 6810 -980 7490 -930
rect 6810 -1030 6930 -980
rect 7190 -1030 7490 -980
rect 7650 -1030 7670 910
rect 6810 -1050 7670 -1030
rect 1990 -1080 2190 -1070
rect 2593 -1120 2599 -1119
rect 1670 -1130 2599 -1120
rect 1670 -1190 1680 -1130
rect 1740 -1170 2599 -1130
rect 1740 -1190 1750 -1170
rect 2593 -1171 2599 -1170
rect 2651 -1171 2657 -1119
rect 1670 -1200 1750 -1190
rect 2950 -1200 3150 -1180
rect 2950 -1210 2970 -1200
rect 1540 -1220 1630 -1210
rect 1540 -1290 1550 -1220
rect 1620 -1230 1630 -1220
rect 1870 -1220 2970 -1210
rect 1870 -1230 1890 -1220
rect 1620 -1280 1890 -1230
rect 2060 -1280 2970 -1220
rect 1620 -1290 2970 -1280
rect 1540 -1300 2970 -1290
rect 1780 -1400 2970 -1300
rect 1780 -1450 1800 -1400
rect 1970 -1440 2970 -1400
rect 3130 -1440 3150 -1200
rect 1970 -1450 3150 -1440
rect 1780 -1460 3150 -1450
rect 5820 -1450 6440 -1440
rect 1670 -1480 1750 -1470
rect 1670 -1540 1680 -1480
rect 1740 -1500 1750 -1480
rect 2593 -1500 2599 -1499
rect 1740 -1540 2599 -1500
rect 1670 -1550 2599 -1540
rect 2593 -1551 2599 -1550
rect 2651 -1551 2657 -1499
rect 5820 -1510 5830 -1450
rect 5950 -1460 6440 -1450
rect 5950 -1510 6260 -1460
rect 6420 -1510 6440 -1460
rect 6930 -1460 7670 -1440
rect 5820 -1520 6440 -1510
rect 6800 -1500 6900 -1490
rect 6540 -1550 6620 -1540
rect 6540 -1560 6550 -1550
rect 690 -1600 1860 -1580
rect 690 -1760 710 -1600
rect 870 -1760 1860 -1600
rect 690 -1780 1860 -1760
rect 1900 -1590 2090 -1580
rect 1900 -1770 2010 -1590
rect 2080 -1770 2090 -1590
rect 6310 -1610 6550 -1560
rect 6610 -1610 6620 -1550
rect 6800 -1560 6810 -1500
rect 6890 -1540 6900 -1500
rect 6930 -1500 6950 -1460
rect 7190 -1500 7490 -1460
rect 6930 -1510 7490 -1500
rect 6890 -1560 7110 -1540
rect 6800 -1600 7110 -1560
rect 7230 -1550 7490 -1510
rect 6540 -1620 6620 -1610
rect 4730 -1650 4930 -1630
rect 2350 -1690 3350 -1680
rect 2350 -1740 2370 -1690
rect 2980 -1700 3350 -1690
rect 2980 -1740 3170 -1700
rect 2350 -1750 3170 -1740
rect 1900 -1780 2090 -1770
rect 3000 -1770 3170 -1750
rect 1670 -1820 1920 -1810
rect 1670 -1880 1680 -1820
rect 1740 -1860 1920 -1820
rect 2120 -1840 2890 -1790
rect 1740 -1880 1750 -1860
rect 1670 -1890 1750 -1880
rect 1540 -1900 1630 -1890
rect 1540 -1970 1550 -1900
rect 1620 -1920 1630 -1900
rect 1780 -1920 1990 -1910
rect 1620 -1970 1800 -1920
rect 1970 -1970 1990 -1920
rect 1540 -1980 1990 -1970
rect 1090 -1990 1290 -1980
rect 1090 -2140 1110 -1990
rect 1270 -2010 1290 -1990
rect 2120 -2010 2170 -1840
rect 3000 -1870 3010 -1770
rect 1270 -2130 2170 -2010
rect 1270 -2140 1290 -2130
rect 1090 -2160 1290 -2140
rect 1540 -2180 1990 -2160
rect 1540 -2250 1550 -2180
rect 1620 -2220 1800 -2180
rect 1620 -2250 1630 -2220
rect 1780 -2230 1800 -2220
rect 1970 -2230 1990 -2180
rect 1780 -2240 1990 -2230
rect 1540 -2260 1630 -2250
rect 1670 -2260 1750 -2250
rect 1670 -2320 1680 -2260
rect 1740 -2280 1750 -2260
rect 2120 -2280 2170 -2130
rect 2210 -1890 2430 -1880
rect 2210 -2230 2220 -1890
rect 2310 -2230 2430 -1890
rect 2210 -2240 2430 -2230
rect 2900 -2250 3010 -1870
rect 1740 -2320 1920 -2280
rect 1670 -2330 1920 -2320
rect 2120 -2330 2890 -2280
rect 3000 -2350 3010 -2250
rect 3070 -2350 3170 -1770
rect 290 -2380 1860 -2360
rect 290 -2540 310 -2380
rect 470 -2540 1860 -2380
rect 290 -2560 1860 -2540
rect 1900 -2370 2090 -2360
rect 3000 -2370 3170 -2350
rect 1900 -2550 2010 -2370
rect 2080 -2550 2090 -2370
rect 2350 -2380 3170 -2370
rect 2350 -2430 2370 -2380
rect 2980 -2420 3170 -2380
rect 3330 -2420 3350 -1700
rect 4730 -1730 4750 -1650
rect 4910 -1730 6320 -1650
rect 6360 -1660 6900 -1650
rect 6360 -1720 6810 -1660
rect 6890 -1720 6900 -1660
rect 6360 -1730 6900 -1720
rect 4730 -1750 4930 -1730
rect 6540 -1770 6620 -1760
rect 6310 -1820 6550 -1770
rect 6540 -1830 6550 -1820
rect 6610 -1830 6620 -1770
rect 6540 -1840 6620 -1830
rect 5820 -1870 6440 -1860
rect 5820 -1930 5830 -1870
rect 5950 -1920 6260 -1870
rect 6420 -1920 6440 -1870
rect 5950 -1930 6440 -1920
rect 5820 -1940 6440 -1930
rect 5460 -2040 7200 -2030
rect 5460 -2140 5470 -2040
rect 5650 -2140 7200 -2040
rect 5460 -2150 7200 -2140
rect 5820 -2250 6440 -2240
rect 5820 -2310 5830 -2250
rect 5950 -2260 6440 -2250
rect 5950 -2310 6260 -2260
rect 6420 -2310 6440 -2260
rect 5820 -2320 6440 -2310
rect 6540 -2350 6620 -2340
rect 6540 -2360 6550 -2350
rect 6310 -2410 6550 -2360
rect 6610 -2410 6620 -2350
rect 6540 -2420 6620 -2410
rect 2980 -2430 3350 -2420
rect 2350 -2440 3350 -2430
rect 5090 -2450 5290 -2430
rect 5090 -2530 5110 -2450
rect 5270 -2530 6320 -2450
rect 6360 -2460 6900 -2450
rect 6360 -2520 6810 -2460
rect 6890 -2520 6900 -2460
rect 6360 -2530 6900 -2520
rect 5090 -2550 5290 -2530
rect 1900 -2560 2090 -2550
rect 6540 -2570 6620 -2560
rect 2593 -2590 2599 -2589
rect 1670 -2600 2599 -2590
rect 1670 -2660 1680 -2600
rect 1740 -2640 2599 -2600
rect 1740 -2660 1750 -2640
rect 2593 -2641 2599 -2640
rect 2651 -2641 2657 -2589
rect 6310 -2620 6550 -2570
rect 6540 -2630 6550 -2620
rect 6610 -2630 6620 -2570
rect 6540 -2640 6620 -2630
rect 6810 -2620 6890 -2600
rect 1540 -2670 1630 -2660
rect 1670 -2670 1750 -2660
rect 5820 -2670 6440 -2660
rect 1540 -2830 1550 -2670
rect 1620 -2700 1630 -2670
rect 1780 -2690 3350 -2680
rect 1780 -2700 1800 -2690
rect 1620 -2740 1800 -2700
rect 1970 -2700 3350 -2690
rect 1970 -2740 3170 -2700
rect 1620 -2810 3170 -2740
rect 1620 -2830 2070 -2810
rect 1540 -2840 2070 -2830
rect 2050 -2850 2070 -2840
rect 2230 -2820 3170 -2810
rect 3330 -2820 3350 -2700
rect 5820 -2730 5830 -2670
rect 5950 -2720 6260 -2670
rect 6420 -2720 6440 -2670
rect 5950 -2730 6440 -2720
rect 5820 -2740 6440 -2730
rect 2230 -2840 3350 -2820
rect 2230 -2850 2250 -2840
rect 2050 -2870 2250 -2850
rect 1920 -2950 1930 -2890
rect 2000 -2910 2010 -2890
rect 2623 -2910 2629 -2909
rect 2000 -2950 2629 -2910
rect 690 -2970 890 -2950
rect 1920 -2960 2629 -2950
rect 2623 -2961 2629 -2960
rect 2681 -2961 2687 -2909
rect 690 -3110 710 -2970
rect 870 -2990 890 -2970
rect 870 -3090 2130 -2990
rect 2180 -3000 2380 -2990
rect 2180 -3080 2290 -3000
rect 2370 -3080 2380 -3000
rect 2180 -3090 2380 -3080
rect 870 -3110 890 -3090
rect 690 -3130 890 -3110
rect 1920 -3130 2200 -3120
rect 1920 -3190 1930 -3130
rect 2000 -3170 2200 -3130
rect 2780 -3130 3350 -3120
rect 2000 -3190 2010 -3170
rect 2780 -3180 2800 -3130
rect 2980 -3140 3350 -3130
rect 2980 -3180 3170 -3140
rect 2780 -3190 3170 -3180
rect 1540 -3210 1630 -3200
rect 1540 -3280 1550 -3210
rect 1620 -3220 1630 -3210
rect 2050 -3220 2260 -3210
rect 1620 -3230 2260 -3220
rect 1620 -3270 2070 -3230
rect 2230 -3270 2260 -3230
rect 1620 -3280 2260 -3270
rect 1540 -3290 2260 -3280
rect 2380 -3230 2750 -3200
rect 2940 -3220 3170 -3190
rect 2380 -3240 2900 -3230
rect 1090 -3310 1290 -3290
rect 1090 -3410 1110 -3310
rect 1270 -3320 1290 -3310
rect 2380 -3320 2420 -3240
rect 1270 -3400 2420 -3320
rect 1270 -3410 1290 -3400
rect 1090 -3430 1290 -3410
rect 1540 -3440 2260 -3430
rect 1540 -3510 1550 -3440
rect 1620 -3450 2260 -3440
rect 1620 -3490 2070 -3450
rect 2230 -3490 2260 -3450
rect 1620 -3500 2260 -3490
rect 1620 -3510 1630 -3500
rect 2050 -3510 2260 -3500
rect 2380 -3480 2420 -3400
rect 2450 -3280 2680 -3270
rect 2710 -3280 2900 -3240
rect 2450 -3440 2460 -3280
rect 2590 -3300 2680 -3280
rect 2940 -3300 3020 -3220
rect 2590 -3320 2690 -3300
rect 2920 -3320 3020 -3300
rect 2590 -3400 2700 -3320
rect 2910 -3400 3020 -3320
rect 2590 -3420 2690 -3400
rect 2920 -3420 3020 -3400
rect 2590 -3440 2680 -3420
rect 2450 -3450 2680 -3440
rect 2710 -3480 2900 -3440
rect 2380 -3490 2900 -3480
rect 1540 -3520 1630 -3510
rect 2380 -3520 2750 -3490
rect 2940 -3500 3020 -3420
rect 3080 -3500 3170 -3220
rect 2940 -3530 3170 -3500
rect 1920 -3590 1930 -3530
rect 2000 -3550 2010 -3530
rect 2780 -3540 3170 -3530
rect 2000 -3590 2200 -3550
rect 1920 -3600 2200 -3590
rect 2780 -3590 2800 -3540
rect 2980 -3580 3170 -3540
rect 3330 -3580 3350 -3140
rect 2980 -3590 3350 -3580
rect 2780 -3600 3350 -3590
rect 290 -3630 490 -3610
rect 290 -3730 310 -3630
rect 470 -3730 2130 -3630
rect 2180 -3640 2380 -3630
rect 2180 -3720 2290 -3640
rect 2370 -3720 2380 -3640
rect 2180 -3730 2380 -3720
rect 290 -3750 490 -3730
rect 2618 -3760 2624 -3759
rect 1920 -3770 2624 -3760
rect 1920 -3830 1930 -3770
rect 2000 -3810 2624 -3770
rect 2000 -3830 2010 -3810
rect 2618 -3811 2624 -3810
rect 2676 -3811 2682 -3759
rect 1540 -3850 1630 -3840
rect 1540 -4000 1550 -3850
rect 1620 -3860 1630 -3850
rect 2050 -3860 2260 -3850
rect 1620 -3870 3350 -3860
rect 1620 -3910 2070 -3870
rect 2230 -3880 3350 -3870
rect 2230 -3910 3170 -3880
rect 1620 -3960 3170 -3910
rect 1620 -3990 1870 -3960
rect 1540 -4010 1620 -4000
rect 1850 -4000 1870 -3990
rect 2030 -4000 3170 -3960
rect 3330 -4000 3350 -3880
rect 1850 -4020 3350 -4000
rect 1740 -4040 1820 -4030
rect 1740 -4100 1750 -4040
rect 1810 -4060 1820 -4040
rect 2623 -4060 2629 -4059
rect 1810 -4100 2629 -4060
rect 1740 -4110 2629 -4100
rect 2623 -4111 2629 -4110
rect 2681 -4111 2687 -4059
rect 690 -4140 890 -4120
rect 690 -4240 710 -4140
rect 870 -4240 1930 -4140
rect 1970 -4150 2190 -4140
rect 1970 -4230 2110 -4150
rect 1970 -4240 2190 -4230
rect 690 -4260 890 -4240
rect 1740 -4280 1990 -4270
rect 1740 -4340 1750 -4280
rect 1810 -4320 1990 -4280
rect 2440 -4280 3350 -4270
rect 1810 -4340 1820 -4320
rect 1740 -4350 1820 -4340
rect 2440 -4340 2460 -4280
rect 3020 -4290 3350 -4280
rect 3020 -4340 3170 -4290
rect 2440 -4350 3170 -4340
rect 1540 -4370 1620 -4360
rect 1540 -4440 1550 -4370
rect 1850 -4380 2060 -4360
rect 1850 -4390 1870 -4380
rect 1620 -4420 1870 -4390
rect 2030 -4420 2060 -4380
rect 3050 -4380 3170 -4350
rect 1620 -4440 2060 -4420
rect 2180 -4440 2940 -4390
rect 1090 -4470 1290 -4450
rect 2180 -4470 2220 -4440
rect 3050 -4470 3060 -4380
rect 1090 -4570 1110 -4470
rect 1270 -4570 2220 -4470
rect 2250 -4480 2530 -4470
rect 2250 -4560 2260 -4480
rect 2340 -4560 2530 -4480
rect 2250 -4570 2530 -4560
rect 2950 -4570 3060 -4470
rect 1090 -4590 1290 -4570
rect 2180 -4600 2220 -4570
rect 1540 -4670 1550 -4600
rect 1620 -4620 2060 -4600
rect 1620 -4660 1870 -4620
rect 2030 -4660 2060 -4620
rect 2180 -4650 2940 -4600
rect 1540 -4680 1620 -4670
rect 1850 -4680 2060 -4660
rect 3050 -4660 3060 -4570
rect 3120 -4660 3170 -4380
rect 3050 -4690 3170 -4660
rect 1740 -4700 1820 -4690
rect 1740 -4760 1750 -4700
rect 1810 -4720 1820 -4700
rect 2440 -4700 3170 -4690
rect 1810 -4760 1990 -4720
rect 1740 -4770 1990 -4760
rect 2440 -4760 2460 -4700
rect 3020 -4750 3170 -4700
rect 3330 -4750 3350 -4290
rect 3020 -4760 3350 -4750
rect 2440 -4770 3350 -4760
rect 290 -4800 490 -4780
rect 290 -4900 310 -4800
rect 470 -4900 1930 -4800
rect 1970 -4810 2190 -4800
rect 1970 -4890 2110 -4810
rect 1970 -4900 2190 -4890
rect 6810 -4900 6820 -2620
rect 6880 -4860 6890 -2620
rect 7010 -4860 7110 -4830
rect 7230 -4860 7240 -1550
rect 6880 -4900 7240 -4860
rect 7300 -4900 7490 -1550
rect 290 -4920 490 -4900
rect 2623 -4930 2629 -4929
rect 1740 -4940 2629 -4930
rect 1740 -5000 1750 -4940
rect 1810 -4980 2629 -4940
rect 1810 -5000 1820 -4980
rect 2623 -4981 2629 -4980
rect 2681 -4981 2687 -4929
rect 1740 -5010 1820 -5000
rect 6810 -4990 7490 -4900
rect 7650 -4990 7670 -1460
rect 6810 -5010 7670 -4990
rect 8150 -4970 8240 3980
rect 8310 -4970 8330 3980
rect 8650 3940 9270 4820
rect 10110 4980 10730 5000
rect 10110 4820 10130 4980
rect 10710 4820 10730 4980
rect 9600 4580 9780 4600
rect 9600 4420 9620 4580
rect 9760 4420 9780 4580
rect 9600 3970 9780 4420
rect 8370 3470 9550 3940
rect 8360 -4940 9560 -4460
rect 1540 -5030 1620 -5020
rect 1540 -5100 1550 -5030
rect 1850 -5040 3350 -5020
rect 1850 -5050 1870 -5040
rect 1620 -5080 1870 -5050
rect 2030 -5080 3170 -5040
rect 1620 -5100 3170 -5080
rect 3150 -5160 3170 -5100
rect 3330 -5160 3350 -5040
rect 8150 -5140 8330 -4970
rect 3150 -5180 3350 -5160
rect 8650 -6290 9270 -4940
rect 9600 -4970 9610 3970
rect 9770 -4970 9780 3970
rect 10110 3940 10730 4820
rect 11050 4580 11230 4600
rect 11050 4420 11070 4580
rect 11210 4420 11230 4580
rect 11050 3980 11230 4420
rect 9830 3470 11010 3940
rect 9820 -4940 11020 -4460
rect 9600 -5140 9780 -4970
rect 10110 -5890 10730 -4940
rect 11050 -4970 11060 3980
rect 11150 -4970 11230 3980
rect 11050 -5140 11230 -4970
rect 10110 -6050 10130 -5890
rect 10710 -6050 10730 -5890
rect 10110 -6070 10730 -6050
rect 8650 -6450 8670 -6290
rect 9250 -6450 9270 -6290
rect 8650 -6470 9270 -6450
<< via1 >>
rect 1280 4810 1340 4820
rect 1280 4760 1330 4810
rect 1330 4760 1340 4810
rect 1280 4580 1340 4590
rect 1280 4530 1330 4580
rect 1330 4530 1340 4580
rect 860 4020 1120 4180
rect 1560 3620 1820 3780
rect 1380 3220 1460 3350
rect 2050 3620 2340 3780
rect 1890 3230 1970 3340
rect 2420 3230 2500 3340
rect 2650 3070 2710 3130
rect 2800 3070 2860 3130
rect 2964 3074 3016 3126
rect 3264 3074 3316 3126
rect 3454 3074 3506 3126
rect 3624 3074 3676 3126
rect 3784 3074 3836 3126
rect 3944 3074 3996 3126
rect 4084 3074 4136 3126
rect 4234 3074 4286 3126
rect 1560 2580 1670 2690
rect 2030 2460 2090 2520
rect 710 1860 870 2400
rect 7200 3070 7260 3130
rect 7340 3070 7400 3130
rect 8670 4820 9250 4980
rect 8170 4420 8310 4580
rect 7748 3068 7808 3128
rect 7886 3068 7946 3128
rect 5144 2394 5196 2446
rect 5830 2370 5950 2440
rect 6660 2310 6740 2390
rect 4740 2160 4920 2240
rect 6430 2160 6500 2240
rect 5144 2044 5196 2096
rect 2030 1740 2090 1800
rect 1560 1570 1670 1680
rect 2030 1450 2090 1510
rect 5830 1960 5950 2030
rect 5470 1830 5650 1900
rect 5830 1700 5950 1770
rect 5110 1430 5270 1510
rect 6430 1490 6500 1570
rect 310 850 470 1390
rect 5830 1290 5950 1360
rect 7490 1300 7650 2430
rect 5830 850 5950 910
rect 1560 640 1670 750
rect 2030 730 2090 790
rect 6550 750 6610 810
rect 6920 780 7000 860
rect 4750 630 4910 710
rect 6810 640 6890 700
rect 6550 530 6610 590
rect 1550 390 1620 460
rect 2970 370 3130 440
rect 5830 430 5950 490
rect 1680 300 1740 360
rect 2599 289 2651 341
rect 710 -110 870 240
rect 2100 -120 2180 240
rect 5470 230 5650 320
rect 5830 50 5950 110
rect 6550 -50 6610 10
rect 1680 -240 1740 -180
rect 1550 -320 1610 -260
rect 1110 -460 1270 -370
rect 1550 -570 1610 -510
rect 2330 -500 2460 -320
rect 1680 -650 1740 -590
rect 310 -1060 470 -710
rect 2100 -1070 2180 -710
rect 2970 -710 3130 -110
rect 5110 -170 5270 -90
rect 6810 -160 6890 -100
rect 6550 -270 6610 -210
rect 5830 -370 5950 -310
rect 7490 -1030 7650 910
rect 1680 -1190 1740 -1130
rect 2599 -1171 2651 -1119
rect 1550 -1290 1620 -1220
rect 2970 -1440 3130 -1200
rect 1680 -1540 1740 -1480
rect 2599 -1551 2651 -1499
rect 5830 -1510 5950 -1450
rect 710 -1760 870 -1600
rect 2010 -1770 2080 -1590
rect 6550 -1610 6610 -1550
rect 6810 -1560 6890 -1500
rect 1680 -1880 1740 -1820
rect 1550 -1970 1620 -1900
rect 1110 -2140 1270 -1990
rect 1550 -2250 1620 -2180
rect 1680 -2320 1740 -2260
rect 2220 -2230 2310 -1890
rect 310 -2540 470 -2380
rect 2010 -2550 2080 -2370
rect 3170 -2420 3330 -1700
rect 4750 -1730 4910 -1650
rect 6810 -1720 6890 -1660
rect 6550 -1830 6610 -1770
rect 5830 -1930 5950 -1870
rect 5470 -2140 5650 -2040
rect 5830 -2310 5950 -2250
rect 6550 -2410 6610 -2350
rect 5110 -2530 5270 -2450
rect 6810 -2520 6890 -2460
rect 1680 -2660 1740 -2600
rect 2599 -2641 2651 -2589
rect 6550 -2630 6610 -2570
rect 1550 -2830 1620 -2670
rect 3170 -2820 3330 -2700
rect 5830 -2730 5950 -2670
rect 1930 -2950 2000 -2890
rect 2629 -2961 2681 -2909
rect 710 -3110 870 -2970
rect 2290 -3080 2370 -3000
rect 1930 -3190 2000 -3130
rect 1550 -3280 1620 -3210
rect 1110 -3410 1270 -3310
rect 1550 -3510 1620 -3440
rect 2460 -3440 2590 -3280
rect 1930 -3590 2000 -3530
rect 3170 -3580 3330 -3140
rect 310 -3730 470 -3630
rect 2290 -3720 2370 -3640
rect 1930 -3830 2000 -3770
rect 2624 -3811 2676 -3759
rect 1550 -4000 1620 -3850
rect 3170 -4000 3330 -3880
rect 1750 -4100 1810 -4040
rect 2629 -4111 2681 -4059
rect 710 -4240 870 -4140
rect 2110 -4230 2190 -4150
rect 1750 -4340 1810 -4280
rect 1550 -4440 1620 -4370
rect 1110 -4570 1270 -4470
rect 2260 -4560 2340 -4480
rect 1550 -4670 1620 -4600
rect 1750 -4760 1810 -4700
rect 3170 -4750 3330 -4290
rect 310 -4900 470 -4800
rect 2110 -4890 2190 -4810
rect 1750 -5000 1810 -4940
rect 2629 -4981 2681 -4929
rect 7490 -4990 7650 -1460
rect 10130 4820 10710 4980
rect 9620 4420 9760 4580
rect 1550 -5100 1620 -5030
rect 3170 -5160 3330 -5040
rect 11070 4420 11210 4580
rect 10130 -6050 10710 -5890
rect 8670 -6450 9250 -6290
<< metal2 >>
rect 8650 4980 9270 5000
rect 1270 4820 1350 4830
rect 1270 4760 1280 4820
rect 1340 4760 1350 4820
rect 8650 4820 8670 4980
rect 9250 4820 9270 4980
rect 8650 4800 9270 4820
rect 10110 4980 10730 5000
rect 10110 4820 10130 4980
rect 10710 4820 10730 4980
rect 10110 4800 10730 4820
rect 1270 4590 1350 4760
rect 1270 4530 1280 4590
rect 1340 4530 1350 4590
rect 1270 4510 1350 4530
rect 8150 4580 8330 4600
rect 8150 4420 8170 4580
rect 8310 4420 8330 4580
rect 8150 4400 8330 4420
rect 9600 4580 9780 4600
rect 9600 4420 9620 4580
rect 9760 4420 9780 4580
rect 9600 4400 9780 4420
rect 11050 4580 11230 4600
rect 11050 4420 11070 4580
rect 11210 4420 11230 4580
rect 11050 4400 11230 4420
rect 840 4180 1140 4200
rect 840 4020 860 4180
rect 1120 4020 1140 4180
rect 840 4000 1140 4020
rect 1540 3780 1840 3800
rect 1540 3620 1560 3780
rect 1820 3620 1840 3780
rect 1540 3600 1840 3620
rect 2030 3780 2360 3800
rect 2030 3620 2050 3780
rect 2340 3620 2360 3780
rect 2030 3600 2360 3620
rect 1090 3220 1380 3350
rect 1460 3340 5660 3350
rect 1460 3230 1890 3340
rect 1970 3230 2420 3340
rect 2500 3230 5660 3340
rect 1460 3220 5660 3230
rect 690 2400 890 2420
rect 690 1860 710 2400
rect 870 1860 890 2400
rect 690 1840 890 1860
rect 290 1390 490 1410
rect 290 850 310 1390
rect 470 850 490 1390
rect 290 830 490 850
rect 690 240 890 260
rect 690 -110 710 240
rect 870 -110 890 240
rect 690 -130 890 -110
rect 1090 -370 1290 3220
rect 2650 3130 2710 3136
rect 1540 2690 1690 2710
rect 1540 2580 1560 2690
rect 1670 2580 1690 2690
rect 1540 1680 1690 2580
rect 2650 2520 2710 3070
rect 2020 2460 2030 2520
rect 2090 2460 2710 2520
rect 2800 3130 2860 3136
rect 2440 1800 2500 2460
rect 2800 2370 2860 3070
rect 2964 3126 3016 3132
rect 2964 3068 3016 3074
rect 3264 3126 3316 3132
rect 3264 3068 3316 3074
rect 3454 3126 3506 3132
rect 3454 3068 3506 3074
rect 3624 3126 3676 3132
rect 3624 3068 3676 3074
rect 3784 3126 3836 3132
rect 3784 3068 3836 3074
rect 3944 3126 3996 3132
rect 3944 3068 3996 3074
rect 4084 3126 4136 3132
rect 4084 3068 4136 3074
rect 4234 3126 4286 3132
rect 4234 3068 4286 3074
rect 2020 1740 2030 1800
rect 2090 1740 2500 1800
rect 2580 2310 2860 2370
rect 1540 1570 1560 1680
rect 1670 1570 1690 1680
rect 1540 750 1690 1570
rect 2580 1510 2640 2310
rect 2965 2155 3015 3068
rect 2020 1450 2030 1510
rect 2090 1450 2640 1510
rect 2775 2105 3015 2155
rect 2440 790 2500 1450
rect 1540 640 1560 750
rect 1670 640 1690 750
rect 2020 730 2030 790
rect 2090 730 2500 790
rect 1540 620 1690 640
rect 1090 -460 1110 -370
rect 1270 -460 1290 -370
rect 290 -710 490 -690
rect 290 -1060 310 -710
rect 470 -1060 490 -710
rect 290 -1080 490 -1060
rect 690 -1600 890 -1580
rect 690 -1760 710 -1600
rect 870 -1760 890 -1600
rect 690 -1780 890 -1760
rect 1090 -1990 1290 -460
rect 1090 -2140 1110 -1990
rect 1270 -2140 1290 -1990
rect 290 -2380 490 -2360
rect 290 -2540 310 -2380
rect 470 -2540 490 -2380
rect 290 -2560 490 -2540
rect 690 -2970 890 -2950
rect 690 -3110 710 -2970
rect 870 -3110 890 -2970
rect 690 -3130 890 -3110
rect 1090 -3310 1290 -2140
rect 1090 -3410 1110 -3310
rect 1270 -3410 1290 -3310
rect 290 -3630 490 -3610
rect 290 -3730 310 -3630
rect 470 -3730 490 -3630
rect 290 -3750 490 -3730
rect 690 -4140 890 -4120
rect 690 -4240 710 -4140
rect 870 -4240 890 -4140
rect 690 -4260 890 -4240
rect 1090 -4470 1290 -3410
rect 1090 -4570 1110 -4470
rect 1270 -4570 1290 -4470
rect 290 -4800 490 -4780
rect 290 -4900 310 -4800
rect 470 -4900 490 -4800
rect 290 -4920 490 -4900
rect 1090 -5470 1290 -4570
rect 1540 460 1620 470
rect 1540 390 1550 460
rect 1540 -260 1620 390
rect 1670 360 1750 370
rect 1670 300 1680 360
rect 1740 300 1750 360
rect 1670 -180 1750 300
rect 2599 341 2651 347
rect 2775 340 2825 2105
rect 2950 440 3150 460
rect 2950 370 2970 440
rect 3130 370 3150 440
rect 2950 350 3150 370
rect 2651 290 2825 340
rect 2599 283 2651 289
rect 2090 240 2470 250
rect 2090 -120 2100 240
rect 2180 -120 2470 240
rect 2090 -130 2470 -120
rect 1670 -240 1680 -180
rect 1740 -240 1750 -180
rect 1670 -250 1750 -240
rect 1540 -320 1550 -260
rect 1610 -320 1620 -260
rect 1540 -510 1620 -320
rect 1540 -570 1550 -510
rect 1610 -570 1620 -510
rect 1540 -1220 1620 -570
rect 2320 -320 2470 -130
rect 2320 -500 2330 -320
rect 2460 -500 2470 -320
rect 1670 -590 1750 -580
rect 1670 -650 1680 -590
rect 1740 -650 1750 -590
rect 1670 -1130 1750 -650
rect 2320 -700 2470 -500
rect 2090 -710 2470 -700
rect 2090 -1070 2100 -710
rect 2180 -1070 2470 -710
rect 2950 -110 3150 -90
rect 2950 -710 2970 -110
rect 3130 -710 3150 -110
rect 2950 -730 3150 -710
rect 2090 -1080 2470 -1070
rect 3265 -1090 3315 3068
rect 1670 -1190 1680 -1130
rect 1740 -1190 1750 -1130
rect 2599 -1119 2651 -1113
rect 2840 -1120 3315 -1090
rect 2651 -1140 3315 -1120
rect 2651 -1170 2890 -1140
rect 2599 -1177 2651 -1171
rect 1670 -1200 1750 -1190
rect 2950 -1200 3150 -1180
rect 1540 -1290 1550 -1220
rect 1540 -1900 1620 -1290
rect 2950 -1440 2970 -1200
rect 3130 -1440 3150 -1200
rect 2950 -1460 3150 -1440
rect 1670 -1480 1750 -1470
rect 1670 -1540 1680 -1480
rect 1740 -1540 1750 -1480
rect 1670 -1820 1750 -1540
rect 2599 -1499 2651 -1493
rect 3455 -1500 3505 3068
rect 2651 -1550 3505 -1500
rect 2599 -1557 2651 -1551
rect 2000 -1590 2320 -1580
rect 2000 -1770 2010 -1590
rect 2080 -1770 2320 -1590
rect 2000 -1780 2320 -1770
rect 1670 -1880 1680 -1820
rect 1740 -1880 1750 -1820
rect 1670 -1890 1750 -1880
rect 2210 -1890 2320 -1780
rect 1540 -1970 1550 -1900
rect 1540 -2180 1620 -1970
rect 1540 -2250 1550 -2180
rect 2210 -2230 2220 -1890
rect 2310 -2230 2320 -1890
rect 1540 -2670 1620 -2250
rect 1670 -2260 1750 -2250
rect 1670 -2320 1680 -2260
rect 1740 -2320 1750 -2260
rect 1670 -2600 1750 -2320
rect 2210 -2360 2320 -2230
rect 2000 -2370 2320 -2360
rect 2000 -2550 2010 -2370
rect 2080 -2550 2320 -2370
rect 3150 -1700 3350 -1680
rect 3150 -2420 3170 -1700
rect 3330 -2420 3350 -1700
rect 3150 -2440 3350 -2420
rect 2000 -2560 2320 -2550
rect 1670 -2660 1680 -2600
rect 1740 -2660 1750 -2600
rect 2599 -2589 2651 -2583
rect 3625 -2590 3675 3068
rect 2651 -2640 3675 -2590
rect 2599 -2647 2651 -2641
rect 1670 -2670 1750 -2660
rect 1540 -2830 1550 -2670
rect 1540 -3210 1620 -2830
rect 3150 -2700 3350 -2680
rect 3150 -2820 3170 -2700
rect 3330 -2820 3350 -2700
rect 3150 -2840 3350 -2820
rect 1920 -2950 1930 -2890
rect 2000 -2950 2010 -2890
rect 1920 -3130 2010 -2950
rect 2629 -2909 2681 -2903
rect 3785 -2910 3835 3068
rect 2681 -2960 3835 -2910
rect 2629 -2967 2681 -2961
rect 2280 -3000 2600 -2990
rect 2280 -3080 2290 -3000
rect 2370 -3080 2600 -3000
rect 2280 -3090 2600 -3080
rect 1920 -3190 1930 -3130
rect 2000 -3190 2010 -3130
rect 1540 -3280 1550 -3210
rect 1540 -3440 1620 -3280
rect 1540 -3510 1550 -3440
rect 1540 -3850 1620 -3510
rect 2450 -3280 2600 -3090
rect 2450 -3440 2460 -3280
rect 2590 -3440 2600 -3280
rect 1920 -3590 1930 -3530
rect 2000 -3590 2010 -3530
rect 1920 -3770 2010 -3590
rect 2450 -3630 2600 -3440
rect 3150 -3140 3350 -3120
rect 3150 -3580 3170 -3140
rect 3330 -3580 3350 -3140
rect 3150 -3600 3350 -3580
rect 2280 -3640 2600 -3630
rect 2280 -3720 2290 -3640
rect 2370 -3720 2600 -3640
rect 2280 -3730 2600 -3720
rect 1920 -3830 1930 -3770
rect 2000 -3830 2010 -3770
rect 2624 -3759 2676 -3753
rect 3945 -3760 3995 3068
rect 2676 -3810 3995 -3760
rect 2624 -3817 2676 -3811
rect 1540 -4000 1550 -3850
rect 1540 -4370 1620 -4000
rect 3150 -3880 3350 -3860
rect 3150 -4000 3170 -3880
rect 3330 -4000 3350 -3880
rect 3150 -4020 3350 -4000
rect 1740 -4040 1820 -4030
rect 1740 -4100 1750 -4040
rect 1810 -4100 1820 -4040
rect 1740 -4280 1820 -4100
rect 2629 -4059 2681 -4053
rect 4085 -4060 4135 3068
rect 2681 -4110 4135 -4060
rect 2629 -4117 2681 -4111
rect 2100 -4150 2350 -4140
rect 2100 -4230 2110 -4150
rect 2190 -4230 2350 -4150
rect 2100 -4240 2350 -4230
rect 1740 -4340 1750 -4280
rect 1810 -4340 1820 -4280
rect 1740 -4350 1820 -4340
rect 1540 -4440 1550 -4370
rect 1540 -4600 1620 -4440
rect 1540 -4670 1550 -4600
rect 1540 -5030 1620 -4670
rect 2250 -4480 2350 -4240
rect 2250 -4560 2260 -4480
rect 2340 -4560 2350 -4480
rect 1740 -4700 1820 -4690
rect 1740 -4760 1750 -4700
rect 1810 -4760 1820 -4700
rect 1740 -4940 1820 -4760
rect 2250 -4800 2350 -4560
rect 3150 -4290 3350 -4270
rect 3150 -4750 3170 -4290
rect 3330 -4750 3350 -4290
rect 3150 -4770 3350 -4750
rect 2100 -4810 2350 -4800
rect 2100 -4890 2110 -4810
rect 2190 -4890 2350 -4810
rect 2100 -4900 2350 -4890
rect 1740 -5000 1750 -4940
rect 1810 -5000 1820 -4940
rect 2629 -4929 2681 -4923
rect 4235 -4930 4285 3068
rect 5144 2446 5196 2452
rect 5144 2388 5196 2394
rect 4730 2240 4930 2250
rect 4730 2160 4740 2240
rect 4920 2160 4930 2240
rect 4730 2150 4930 2160
rect 5145 2096 5195 2388
rect 5138 2044 5144 2096
rect 5196 2044 5202 2096
rect 5460 1900 5660 3220
rect 7200 3130 7260 3136
rect 5460 1830 5470 1900
rect 5650 1830 5660 1900
rect 5090 1510 5290 1530
rect 5090 1430 5110 1510
rect 5270 1430 5290 1510
rect 5090 1410 5290 1430
rect 4730 710 4930 730
rect 4730 630 4750 710
rect 4910 630 4930 710
rect 4730 610 4930 630
rect 5460 320 5660 1830
rect 5460 230 5470 320
rect 5650 230 5660 320
rect 5090 -90 5290 -70
rect 5090 -170 5110 -90
rect 5270 -170 5290 -90
rect 5090 -190 5290 -170
rect 4730 -1650 4930 -1630
rect 4730 -1730 4750 -1650
rect 4910 -1730 4930 -1650
rect 4730 -1750 4930 -1730
rect 5460 -2040 5660 230
rect 5460 -2140 5470 -2040
rect 5650 -2140 5660 -2040
rect 5090 -2450 5290 -2430
rect 5090 -2530 5110 -2450
rect 5270 -2530 5290 -2450
rect 5090 -2550 5290 -2530
rect 2681 -4980 4285 -4930
rect 2629 -4987 2681 -4981
rect 1740 -5010 1820 -5000
rect 1540 -5100 1550 -5030
rect 1540 -5110 1620 -5100
rect 3150 -5040 3350 -5020
rect 3150 -5160 3170 -5040
rect 3330 -5160 3350 -5040
rect 3150 -5180 3350 -5160
rect 5460 -5470 5660 -2140
rect 5820 3029 5960 3040
rect 5820 2911 5831 3029
rect 5949 2911 5960 3029
rect 5820 2440 5960 2911
rect 5820 2370 5830 2440
rect 5950 2370 5960 2440
rect 5820 2030 5960 2370
rect 6650 2390 6750 2400
rect 6650 2310 6660 2390
rect 6740 2310 6750 2390
rect 6650 2250 6750 2310
rect 6420 2240 6750 2250
rect 6420 2160 6430 2240
rect 6500 2160 6750 2240
rect 6420 2150 6750 2160
rect 5820 1960 5830 2030
rect 5950 1960 5960 2030
rect 5820 1770 5960 1960
rect 5820 1700 5830 1770
rect 5950 1700 5960 1770
rect 5820 1360 5960 1700
rect 6650 1580 6750 2150
rect 6420 1570 6750 1580
rect 6420 1490 6430 1570
rect 6500 1490 6750 1570
rect 6420 1480 6750 1490
rect 5820 1290 5830 1360
rect 5950 1290 5960 1360
rect 5820 910 5960 1290
rect 7200 1180 7260 3070
rect 5820 850 5830 910
rect 5950 850 5960 910
rect 5820 490 5960 850
rect 6550 1120 7260 1180
rect 7340 3130 7400 3136
rect 6550 820 6610 1120
rect 7340 1050 7400 3070
rect 7748 3128 7808 3134
rect 7470 2430 7670 2450
rect 7470 1300 7490 2430
rect 7650 1300 7670 2430
rect 7470 1280 7670 1300
rect 6680 990 7400 1050
rect 6540 810 6620 820
rect 6540 750 6550 810
rect 6610 750 6620 810
rect 6540 740 6620 750
rect 6550 600 6610 740
rect 6540 590 6620 600
rect 6540 530 6550 590
rect 6610 530 6620 590
rect 6540 520 6620 530
rect 5820 430 5830 490
rect 5950 430 5960 490
rect 5820 110 5960 430
rect 6680 150 6740 990
rect 7470 910 7670 930
rect 5820 50 5830 110
rect 5950 50 5960 110
rect 5820 -310 5960 50
rect 6550 90 6740 150
rect 6800 860 7010 870
rect 6800 780 6920 860
rect 7000 780 7010 860
rect 6800 770 7010 780
rect 6800 700 6900 770
rect 6800 640 6810 700
rect 6890 640 6900 700
rect 6550 20 6610 90
rect 6540 10 6620 20
rect 6540 -50 6550 10
rect 6610 -50 6620 10
rect 6540 -60 6620 -50
rect 6550 -200 6610 -60
rect 6800 -100 6900 640
rect 6800 -160 6810 -100
rect 6890 -160 6900 -100
rect 6800 -170 6900 -160
rect 6540 -210 6620 -200
rect 6540 -270 6550 -210
rect 6610 -270 6620 -210
rect 6540 -280 6620 -270
rect 5820 -370 5830 -310
rect 5950 -370 5960 -310
rect 5820 -1450 5960 -370
rect 7470 -1030 7490 910
rect 7650 -1030 7670 910
rect 7470 -1050 7670 -1030
rect 7748 -1180 7808 3068
rect 5820 -1510 5830 -1450
rect 5950 -1510 5960 -1450
rect 5820 -1870 5960 -1510
rect 6550 -1240 7808 -1180
rect 7886 3128 7946 3134
rect 6550 -1540 6610 -1240
rect 7886 -1310 7946 3068
rect 6680 -1370 7946 -1310
rect 6540 -1550 6620 -1540
rect 6540 -1610 6550 -1550
rect 6610 -1610 6620 -1550
rect 6540 -1620 6620 -1610
rect 6550 -1760 6610 -1620
rect 6540 -1770 6620 -1760
rect 6540 -1830 6550 -1770
rect 6610 -1830 6620 -1770
rect 6540 -1840 6620 -1830
rect 5820 -1930 5830 -1870
rect 5950 -1930 5960 -1870
rect 5820 -2250 5960 -1930
rect 6680 -2210 6740 -1370
rect 7470 -1460 7670 -1440
rect 5820 -2310 5830 -2250
rect 5950 -2310 5960 -2250
rect 5820 -2670 5960 -2310
rect 6550 -2270 6740 -2210
rect 6800 -1500 6900 -1490
rect 6800 -1560 6810 -1500
rect 6890 -1560 6900 -1500
rect 6800 -1660 6900 -1560
rect 6800 -1720 6810 -1660
rect 6890 -1720 6900 -1660
rect 6550 -2340 6610 -2270
rect 6540 -2350 6620 -2340
rect 6540 -2410 6550 -2350
rect 6610 -2410 6620 -2350
rect 6540 -2420 6620 -2410
rect 6550 -2560 6610 -2420
rect 6800 -2460 6900 -1720
rect 6800 -2520 6810 -2460
rect 6890 -2520 6900 -2460
rect 6800 -2530 6900 -2520
rect 6540 -2570 6620 -2560
rect 6540 -2630 6550 -2570
rect 6610 -2630 6620 -2570
rect 6540 -2640 6620 -2630
rect 5820 -2730 5830 -2670
rect 5950 -2730 5960 -2670
rect 5820 -2740 5960 -2730
rect 7470 -4990 7490 -1460
rect 7650 -4990 7670 -1460
rect 7470 -5010 7670 -4990
rect 10740 -5470 10980 -5450
rect 1090 -5670 10760 -5470
rect 10960 -5670 10980 -5470
rect 10740 -5690 10980 -5670
rect 10110 -5890 10730 -5870
rect 10110 -6050 10130 -5890
rect 10710 -6050 10730 -5890
rect 10110 -6070 10730 -6050
rect 8650 -6290 9270 -6270
rect 8650 -6450 8670 -6290
rect 9250 -6450 9270 -6290
rect 8650 -6470 9270 -6450
<< via2 >>
rect 8670 4820 9250 4980
rect 10130 4820 10710 4980
rect 8170 4420 8310 4580
rect 9620 4420 9760 4580
rect 11070 4420 11210 4580
rect 860 4020 1120 4180
rect 1560 3620 1820 3780
rect 2050 3620 2340 3780
rect 710 1860 870 2400
rect 310 850 470 1390
rect 710 -110 870 240
rect 310 -1060 470 -710
rect 710 -1760 870 -1600
rect 310 -2540 470 -2380
rect 710 -3110 870 -2970
rect 310 -3730 470 -3630
rect 710 -4240 870 -4140
rect 310 -4900 470 -4800
rect 2970 370 3130 440
rect 2970 -710 3130 -110
rect 2970 -1440 3130 -1200
rect 3170 -2420 3330 -1700
rect 3170 -2820 3330 -2700
rect 3170 -3580 3330 -3140
rect 3170 -4000 3330 -3880
rect 3170 -4750 3330 -4290
rect 4740 2160 4920 2240
rect 5110 1430 5270 1510
rect 4750 630 4910 710
rect 5110 -170 5270 -90
rect 4750 -1730 4910 -1650
rect 5110 -2530 5270 -2450
rect 3170 -5160 3330 -5040
rect 5831 2911 5949 3029
rect 7490 1300 7650 2430
rect 7490 -1030 7650 910
rect 7490 -4990 7650 -1460
rect 10760 -5670 10960 -5470
rect 10130 -6050 10710 -5890
rect 8670 -6450 9250 -6290
<< metal3 >>
rect 8650 4980 9270 5000
rect 8650 4820 8670 4980
rect 9250 4820 9270 4980
rect 8650 4800 9270 4820
rect 10110 4980 10730 5000
rect 10110 4820 10130 4980
rect 10710 4820 10730 4980
rect 10110 4800 10730 4820
rect 7470 4580 11230 4600
rect 7470 4420 8170 4580
rect 8310 4420 9620 4580
rect 9760 4420 11070 4580
rect 11210 4420 11230 4580
rect 7470 4400 11230 4420
rect 840 4180 1140 4200
rect 840 4020 860 4180
rect 1120 4020 1140 4180
rect 840 4000 1140 4020
rect 7470 3800 7670 4400
rect 634 3600 640 3800
rect 840 3780 7670 3800
rect 840 3620 1560 3780
rect 1820 3620 2050 3780
rect 2340 3620 7670 3780
rect 840 3600 7670 3620
rect 690 2400 890 2420
rect 690 1860 710 2400
rect 870 1860 890 2400
rect 290 1390 490 1410
rect 290 850 310 1390
rect 470 850 490 1390
rect 290 830 490 850
rect 690 240 890 1860
rect 690 -110 710 240
rect 870 -110 890 240
rect 290 -710 490 -690
rect 290 -1060 310 -710
rect 470 -1060 490 -710
rect 290 -1080 490 -1060
rect 690 -1600 890 -110
rect 2950 440 3150 3600
rect 5826 3029 5954 3600
rect 5826 2911 5831 3029
rect 5949 2911 5954 3029
rect 5826 2906 5954 2911
rect 7470 2430 7670 3600
rect 2950 370 2970 440
rect 3130 370 3150 440
rect 2950 -110 3150 370
rect 2950 -710 2970 -110
rect 3130 -710 3150 -110
rect 2950 -1200 3150 -710
rect 2950 -1440 2970 -1200
rect 3130 -1400 3150 -1200
rect 4730 2240 4930 2250
rect 4730 2160 4740 2240
rect 4920 2160 4930 2240
rect 4730 710 4930 2160
rect 5090 1510 5290 1530
rect 5090 1430 5110 1510
rect 5270 1430 5290 1510
rect 5090 1410 5290 1430
rect 4730 630 4750 710
rect 4910 630 4930 710
rect 3130 -1440 3350 -1400
rect 2950 -1600 3350 -1440
rect 690 -1760 710 -1600
rect 870 -1760 890 -1600
rect 290 -2380 490 -2360
rect 290 -2540 310 -2380
rect 470 -2540 490 -2380
rect 290 -2560 490 -2540
rect 690 -2970 890 -1760
rect 690 -3110 710 -2970
rect 870 -3110 890 -2970
rect 290 -3630 490 -3610
rect 290 -3730 310 -3630
rect 470 -3730 490 -3630
rect 290 -3750 490 -3730
rect 690 -4140 890 -3110
rect 690 -4240 710 -4140
rect 870 -4240 890 -4140
rect 290 -4800 490 -4780
rect 290 -4900 310 -4800
rect 470 -4900 490 -4800
rect 290 -4920 490 -4900
rect 690 -5870 890 -4240
rect 3150 -1700 3350 -1600
rect 3150 -2420 3170 -1700
rect 3330 -2420 3350 -1700
rect 3150 -2700 3350 -2420
rect 3150 -2820 3170 -2700
rect 3330 -2820 3350 -2700
rect 3150 -3140 3350 -2820
rect 3150 -3580 3170 -3140
rect 3330 -3580 3350 -3140
rect 3150 -3880 3350 -3580
rect 3150 -4000 3170 -3880
rect 3330 -4000 3350 -3880
rect 3150 -4290 3350 -4000
rect 3150 -4750 3170 -4290
rect 3330 -4750 3350 -4290
rect 3150 -5040 3350 -4750
rect 3150 -5160 3170 -5040
rect 3330 -5160 3350 -5040
rect 3150 -5180 3350 -5160
rect 4730 -1650 4930 630
rect 7470 1300 7490 2430
rect 7650 1300 7670 2430
rect 7470 910 7670 1300
rect 5090 -90 5290 -70
rect 5090 -170 5110 -90
rect 5270 -170 5290 -90
rect 5090 -190 5290 -170
rect 4730 -1730 4750 -1650
rect 4910 -1730 4930 -1650
rect 4730 -5870 4930 -1730
rect 7470 -1030 7490 910
rect 7650 -1030 7670 910
rect 7470 -1460 7670 -1030
rect 5090 -2450 5290 -2430
rect 5090 -2530 5110 -2450
rect 5270 -2530 5290 -2450
rect 5090 -2550 5290 -2530
rect 7470 -4990 7490 -1460
rect 7650 -4990 7670 -1460
rect 7470 -5010 7670 -4990
rect 10740 -5465 10980 -5450
rect 10740 -5675 10755 -5465
rect 10965 -5675 10980 -5465
rect 10740 -5690 10980 -5675
rect 690 -5890 10760 -5870
rect 690 -6050 10130 -5890
rect 10710 -6050 10760 -5890
rect 690 -6070 10760 -6050
rect 10960 -6070 10966 -5870
rect 8650 -6290 9270 -6270
rect 8650 -6450 8670 -6290
rect 9250 -6450 9270 -6290
rect 8650 -6470 9270 -6450
<< via3 >>
rect 8670 4820 9250 4980
rect 10130 4820 10710 4980
rect 860 4020 1120 4180
rect 640 3600 840 3800
rect 310 850 470 1390
rect 310 -1060 470 -710
rect 5110 1430 5270 1510
rect 310 -2540 470 -2380
rect 310 -3730 470 -3630
rect 310 -4900 470 -4800
rect 5110 -170 5270 -90
rect 5110 -2530 5270 -2450
rect 10755 -5470 10965 -5465
rect 10755 -5670 10760 -5470
rect 10760 -5670 10960 -5470
rect 10960 -5670 10965 -5470
rect 10755 -5675 10965 -5670
rect 10760 -6070 10960 -5870
rect 8670 -6450 9250 -6290
<< metal4 >>
rect 6580 4980 11230 5000
rect 6580 4820 8670 4980
rect 9250 4820 10130 4980
rect 10710 4820 11230 4980
rect 6580 4800 11230 4820
rect 6580 4200 6780 4800
rect 0 4180 6780 4200
rect 0 4020 860 4180
rect 1120 4020 6780 4180
rect 0 4000 6780 4020
rect 639 3800 841 3801
rect 0 3600 640 3800
rect 840 3600 841 3800
rect 639 3599 841 3600
rect 5090 1510 5290 1530
rect 5090 1430 5110 1510
rect 5270 1430 5290 1510
rect 290 1390 490 1410
rect 290 850 310 1390
rect 470 850 490 1390
rect 290 -710 490 850
rect 290 -1060 310 -710
rect 470 -1060 490 -710
rect 290 -2380 490 -1060
rect 290 -2540 310 -2380
rect 470 -2540 490 -2380
rect 290 -3630 490 -2540
rect 290 -3730 310 -3630
rect 470 -3730 490 -3630
rect 290 -4800 490 -3730
rect 290 -4900 310 -4800
rect 470 -4900 490 -4800
rect 290 -6270 490 -4900
rect 5090 -90 5290 1430
rect 5090 -170 5110 -90
rect 5270 -170 5290 -90
rect 5090 -2450 5290 -170
rect 5090 -2530 5110 -2450
rect 5270 -2530 5290 -2450
rect 5090 -6270 5290 -2530
rect 10740 -5465 10980 -5450
rect 10740 -5675 10755 -5465
rect 10965 -5470 10980 -5465
rect 10965 -5670 11390 -5470
rect 10965 -5675 10980 -5670
rect 10740 -5690 10980 -5675
rect 10759 -5870 10961 -5869
rect 10759 -6070 10760 -5870
rect 10960 -6070 11390 -5870
rect 10759 -6071 10961 -6070
rect 290 -6290 11390 -6270
rect 290 -6450 8670 -6290
rect 9250 -6450 11390 -6290
rect 290 -6470 11390 -6450
use sky130_fd_pr__nfet_01v8_ATLS57  sky130_fd_pr__nfet_01v8_ATLS57_0 csdac_nom__devices
timestamp 1723780759
transform -1 0 1971 0 -1 -890
box -211 -410 211 410
use sky130_fd_pr__nfet_01v8_HZS9GD  XMB0 csdac_nom__devices
timestamp 1723780759
transform 0 1 7060 -1 0 -3224
box -1796 -260 1796 260
use sky130_fd_pr__nfet_01v8_FMHZDY  XMB1 csdac_nom__devices
timestamp 1723780759
transform 0 1 7060 -1 0 -64
box -996 -260 996 260
use sky130_fd_pr__nfet_01v8_AHZR5K  XMB2 csdac_nom__devices
timestamp 1723780759
transform 0 1 6950 -1 0 1866
box -596 -260 596 260
use sky130_fd_pr__nfet_01v8_BHEWB6  XMB3 csdac_nom__devices
timestamp 1723780759
transform 1 0 2736 0 1 -4520
box -406 -260 406 260
use sky130_fd_pr__nfet_01v8_FMMQLY  XMB4 csdac_nom__devices
timestamp 1723780759
transform 1 0 2806 0 1 -3360
box -296 -260 296 260
use sky130_fd_pr__nfet_01v8_C4RU6Y  XMB5 csdac_nom__devices
timestamp 1723780759
transform 1 0 2666 0 1 -2060
box -426 -400 426 400
use sky130_fd_pr__nfet_01v8_N5FCK4  XMB6 csdac_nom__devices
timestamp 1723780759
transform 1 0 2656 0 1 -410
box -246 -320 246 320
use sky130_fd_pr__nfet_01v8_8TEC39  XMB7 csdac_nom__devices
timestamp 1723780759
transform 0 -1 2180 1 0 2886
box -246 -420 246 420
use sky130_fd_pr__nfet_01v8_SMGLWN  XMmirror csdac_nom__devices
timestamp 1723780759
transform 1 0 1505 0 1 4667
box -246 -260 246 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMN0 csdac_nom__devices
timestamp 1723780759
transform 1 0 6341 0 1 -1690
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMN1
timestamp 1723780759
transform 1 0 6341 0 1 670
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMN2
timestamp 1723780759
transform 1 0 6301 0 1 2200
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMN3
timestamp 1723780759
transform 1 0 1951 0 1 -4190
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMN4
timestamp 1723780759
transform 1 0 2151 0 1 -3040
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_648S5X  XMN5 csdac_nom__devices
timestamp 1723780759
transform 1 0 1881 0 1 -1680
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_ATLS57  XMN6
timestamp 1723780759
transform -1 0 1971 0 -1 60
box -211 -410 211 410
use sky130_fd_pr__nfet_01v8_J2SMEF  XMN7 csdac_nom__devices
timestamp 1723780759
transform 1 0 1971 0 1 2130
box -211 -510 211 510
use sky130_fd_pr__nfet_01v8_L9ESAD  XMP0
timestamp 1723780759
transform 1 0 6341 0 1 -2490
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMP1
timestamp 1723780759
transform 1 0 6341 0 1 -130
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMP2
timestamp 1723780759
transform 1 0 6301 0 1 1530
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMP3
timestamp 1723780759
transform 1 0 1951 0 1 -4850
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XMP4
timestamp 1723780759
transform 1 0 2151 0 1 -3680
box -211 -260 211 260
use sky130_fd_pr__nfet_01v8_648S5X  XMP5
timestamp 1723780759
transform 1 0 1881 0 1 -2460
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_J2SMEF  XMP7
timestamp 1723780759
transform 1 0 1971 0 1 1120
box -211 -510 211 510
use sky130_fd_pr__pfet_01v8_XJ7GBL  XMprog csdac_nom__devices
timestamp 1723780759
transform 1 0 1031 0 1 4669
box -211 -269 211 269
use sky130_fd_pr__res_high_po_5p73_MRHKYZ  XR5 csdac_nom__devices
timestamp 1723782672
transform 1 0 8959 0 1 -498
box -739 -4582 739 4582
use sky130_fd_pr__res_high_po_5p73_MRHKYZ  XR6
timestamp 1723782672
transform 1 0 10419 0 1 -498
box -739 -4582 739 4582
<< labels >>
flabel metal1 2170 830 2380 2830 0 FreeSans 800 0 0 0 IS7
flabel metal2 2320 -320 2470 250 0 FreeSans 800 0 0 0 IS6
flabel metal2 2080 -1780 2320 -1580 0 FreeSans 800 0 0 0 IS5
flabel metal2 2450 -3280 2600 -2990 0 FreeSans 800 0 0 0 IS4
flabel metal2 2250 -4480 2350 -4140 0 FreeSans 800 0 0 0 IS3
flabel metal2 6500 2150 6750 2250 0 FreeSans 800 0 0 0 IS2
flabel metal2 6800 -100 6900 640 0 FreeSans 800 0 0 0 IS1
flabel metal2 6800 -2460 6900 -1720 0 FreeSans 800 0 0 0 IS0
flabel metal4 0 4000 300 4200 0 FreeSans 1120 0 0 0 vcc
port 21 nsew
flabel metal4 0 3600 300 3800 0 FreeSans 1120 0 0 0 vss
port 22 nsew
flabel metal4 11090 -6470 11390 -6270 0 FreeSans 640 0 0 0 Vpos
port 23 nsew
flabel metal4 11090 -6070 11390 -5870 0 FreeSans 640 0 0 0 Vneg
port 24 nsew
flabel metal4 11090 -5670 11390 -5470 0 FreeSans 640 0 0 0 Vbias
port 25 nsew
flabel metal1 3194 5256 3394 5456 0 FreeSans 640 0 0 0 p6
port 14 nsew
flabel metal1 3594 5256 3794 5456 0 FreeSans 640 0 0 0 n5
port 13 nsew
flabel metal1 3994 5256 4194 5456 0 FreeSans 640 0 0 0 p5
port 12 nsew
flabel metal1 4394 5256 4594 5456 0 FreeSans 640 0 0 0 n4
port 11 nsew
flabel metal1 4794 5256 4994 5456 0 FreeSans 640 0 0 0 p4
port 10 nsew
flabel metal1 5194 5256 5394 5456 0 FreeSans 640 0 0 0 n3
port 9 nsew
flabel metal1 5594 5256 5794 5456 0 FreeSans 640 0 0 0 p3
port 8 nsew
flabel metal1 5994 5256 6194 5456 0 FreeSans 640 0 0 0 n2
port 7 nsew
flabel metal1 6394 5256 6594 5456 0 FreeSans 640 0 0 0 p2
port 6 nsew
flabel metal1 6794 5256 6994 5456 0 FreeSans 640 0 0 0 n1
port 5 nsew
flabel metal1 7194 5256 7394 5456 0 FreeSans 640 0 0 0 p1
port 4 nsew
flabel metal1 7594 5256 7794 5456 0 FreeSans 640 0 0 0 n0
port 3 nsew
flabel metal1 7994 5256 8194 5456 0 FreeSans 640 0 0 0 p0
port 2 nsew
flabel metal1 2794 5256 2994 5456 0 FreeSans 640 0 0 0 n6
port 15 nsew
flabel metal1 2394 5256 2594 5456 0 FreeSans 640 0 0 0 p7
port 16 nsew
flabel metal1 1994 5256 2194 5456 0 FreeSans 640 0 0 0 n7
port 17 nsew
<< end >>

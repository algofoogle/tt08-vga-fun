magic
tech sky130A
timestamp 1723780759
<< pwell >>
rect -123 -210 123 210
<< nmos >>
rect -25 -105 25 105
<< ndiff >>
rect -54 99 -25 105
rect -54 -99 -48 99
rect -31 -99 -25 99
rect -54 -105 -25 -99
rect 25 99 54 105
rect 25 -99 31 99
rect 48 -99 54 99
rect 25 -105 54 -99
<< ndiffc >>
rect -48 -99 -31 99
rect 31 -99 48 99
<< psubdiff >>
rect -105 175 -57 192
rect 57 175 105 192
rect -105 144 -88 175
rect 88 144 105 175
rect -105 -175 -88 -144
rect 88 -175 105 -144
rect -105 -192 -57 -175
rect 57 -192 105 -175
<< psubdiffcont >>
rect -57 175 57 192
rect -105 -144 -88 144
rect 88 -144 105 144
rect -57 -192 57 -175
<< poly >>
rect -25 141 25 149
rect -25 124 -17 141
rect 17 124 25 141
rect -25 105 25 124
rect -25 -124 25 -105
rect -25 -141 -17 -124
rect 17 -141 25 -124
rect -25 -149 25 -141
<< polycont >>
rect -17 124 17 141
rect -17 -141 17 -124
<< locali >>
rect -105 175 -57 192
rect 57 175 105 192
rect -105 144 -88 175
rect 88 144 105 175
rect -25 124 -17 141
rect 17 124 25 141
rect -48 99 -31 107
rect -48 -107 -31 -99
rect 31 99 48 107
rect 31 -107 48 -99
rect -25 -141 -17 -124
rect 17 -141 25 -124
rect -105 -175 -88 -144
rect 88 -175 105 -144
rect -105 -192 -57 -175
rect 57 -192 105 -175
<< viali >>
rect -17 124 17 141
rect -48 -99 -31 99
rect 31 -99 48 99
rect -17 -141 17 -124
<< metal1 >>
rect -23 141 23 144
rect -23 124 -17 141
rect 17 124 23 141
rect -23 121 23 124
rect -51 99 -28 105
rect -51 -99 -48 99
rect -31 -99 -28 99
rect -51 -105 -28 -99
rect 28 99 51 105
rect 28 -99 31 99
rect 48 -99 51 99
rect 28 -105 51 -99
rect -23 -124 23 -121
rect -23 -141 -17 -124
rect 17 -141 23 -124
rect -23 -144 23 -141
<< properties >>
string FIXED_BBOX -96 -183 96 183
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2.1 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
